
/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : pfb_8Mmax_16iw_16ow_10tps_dp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data                                                     
//
//
/*****************************************************************************/


module pfb_8Mmax_16iw_16ow_10tps_dp_rom
(
  input clk, 
  input wea,
  input [6:0] addra,
  input [6:0] addrb,
  input [24:0] dia,
  output [24:0] dob
);

(* rom_style = "block" *) reg [24:0] rom [127:0];
reg [6:0] addra_d;
reg [6:0] addrb_d;
reg [24:0] dob_d;
reg [24:0] rom_pipea;
reg [24:0] dia_d;
reg wea_d;

assign dob = dob_d;

initial
begin
    rom[0] = 25'b1111011111111110101111101;
    rom[1] = 25'b1111100001010001111110100;
    rom[2] = 25'b1111100101000101111100000;
    rom[3] = 25'b1111101011001001101110101;
    rom[4] = 25'b1111110011000010010100100;
    rom[5] = 25'b1111111100001100001001000;
    rom[6] = 25'b0000000101111101001110010;
    rom[7] = 25'b0000001111100111110001100;
    rom[8] = 25'b0000011000011101000000100;
    rom[9] = 25'b0000011111110000001001010;
    rom[10] = 25'b0000100100111001010110010;
    rom[11] = 25'b0000100111011000100000011;
    rom[12] = 25'b0000100110110111101000011;
    rom[13] = 25'b0000100011001100110001001;
    rom[14] = 25'b0000011100011011010001100;
    rom[15] = 25'b0000010010110100010111011;
    rom[16] = 25'b0000000110110110111000101;
    rom[17] = 25'b1111111001001110010000000;
    rom[18] = 25'b1111101010110000100111100;
    rom[19] = 25'b1111011100011100010101101;
    rom[20] = 25'b1111001111010100110011011;
    rom[21] = 25'b1111000100011110110101110;
    rom[22] = 25'b1110111100111100110110100;
    rom[23] = 25'b1110111001101010111001000;
    rom[24] = 25'b1110111011011010111010101;
    rom[25] = 25'b1111000010110001011011101;
    rom[26] = 25'b1111010000000010101110011;
    rom[27] = 25'b1111100011010000111000101;
    rom[28] = 25'b1111111100001010110000011;
    rom[29] = 25'b0000011010001011111001011;
    rom[30] = 25'b0000111100011101100110000;
    rom[31] = 25'b0001100001111000111011000;
    rom[32] = 25'b0010001001001001101110110;
    rom[33] = 25'b0010110000110010011101111;
    rom[34] = 25'b0011010111010000100100000;
    rom[35] = 25'b0011111011000001010000100;
    rom[36] = 25'b0100011010100110011111000;
    rom[37] = 25'b0100110100101011101000011;
    rom[38] = 25'b0101001000001001110111000;
    rom[39] = 25'b0101010100001011110001001;
    rom[40] = 25'b0101011000010000001010001;
    rom[41] = 25'b0101010100001011110001001;
    rom[42] = 25'b0101001000001001110111000;
    rom[43] = 25'b0100110100101011101000011;
    rom[44] = 25'b0100011010100110011111000;
    rom[45] = 25'b0011111011000001010000100;
    rom[46] = 25'b0011010111010000100100000;
    rom[47] = 25'b0010110000110010011101111;
    rom[48] = 25'b0010001001001001101110110;
    rom[49] = 25'b0001100001111000111011000;
    rom[50] = 25'b0000111100011101100110000;
    rom[51] = 25'b0000011010001011111001011;
    rom[52] = 25'b1111111100001010110000011;
    rom[53] = 25'b1111100011010000111000101;
    rom[54] = 25'b1111010000000010101110011;
    rom[55] = 25'b1111000010110001011011101;
    rom[56] = 25'b1110111011011010111010101;
    rom[57] = 25'b1110111001101010111001000;
    rom[58] = 25'b1110111100111100110110100;
    rom[59] = 25'b1111000100011110110101110;
    rom[60] = 25'b1111001111010100110011011;
    rom[61] = 25'b1111011100011100010101101;
    rom[62] = 25'b1111101010110000100111100;
    rom[63] = 25'b1111111001001110010000000;
    rom[64] = 25'b0000000110110110111000101;
    rom[65] = 25'b0000010010110100010111011;
    rom[66] = 25'b0000011100011011010001100;
    rom[67] = 25'b0000100011001100110001001;
    rom[68] = 25'b0000100110110111101000011;
    rom[69] = 25'b0000100111011000100000011;
    rom[70] = 25'b0000100100111001010110010;
    rom[71] = 25'b0000011111110000001001010;
    rom[72] = 25'b0000011000011101000000100;
    rom[73] = 25'b0000001111100111110001100;
    rom[74] = 25'b0000000101111101001110010;
    rom[75] = 25'b1111111100001100001001000;
    rom[76] = 25'b1111110011000010010100100;
    rom[77] = 25'b1111101011001001101110101;
    rom[78] = 25'b1111100101000101111100000;
    rom[79] = 25'b1111100001010001111110100;
    rom[80] = 25'b0000000000000000000000000;
    rom[81] = 25'b0000000000000000000000000;
    rom[82] = 25'b0000000000000000000000000;
    rom[83] = 25'b0000000000000000000000000;
    rom[84] = 25'b0000000000000000000000000;
    rom[85] = 25'b0000000000000000000000000;
    rom[86] = 25'b0000000000000000000000000;
    rom[87] = 25'b0000000000000000000000000;
    rom[88] = 25'b0000000000000000000000000;
    rom[89] = 25'b0000000000000000000000000;
    rom[90] = 25'b0000000000000000000000000;
    rom[91] = 25'b0000000000000000000000000;
    rom[92] = 25'b0000000000000000000000000;
    rom[93] = 25'b0000000000000000000000000;
    rom[94] = 25'b0000000000000000000000000;
    rom[95] = 25'b0000000000000000000000000;
    rom[96] = 25'b0000000000000000000000000;
    rom[97] = 25'b0000000000000000000000000;
    rom[98] = 25'b0000000000000000000000000;
    rom[99] = 25'b0000000000000000000000000;
    rom[100] = 25'b0000000000000000000000000;
    rom[101] = 25'b0000000000000000000000000;
    rom[102] = 25'b0000000000000000000000000;
    rom[103] = 25'b0000000000000000000000000;
    rom[104] = 25'b0000000000000000000000000;
    rom[105] = 25'b0000000000000000000000000;
    rom[106] = 25'b0000000000000000000000000;
    rom[107] = 25'b0000000000000000000000000;
    rom[108] = 25'b0000000000000000000000000;
    rom[109] = 25'b0000000000000000000000000;
    rom[110] = 25'b0000000000000000000000000;
    rom[111] = 25'b0000000000000000000000000;
    rom[112] = 25'b0000000000000000000000000;
    rom[113] = 25'b0000000000000000000000000;
    rom[114] = 25'b0000000000000000000000000;
    rom[115] = 25'b0000000000000000000000000;
    rom[116] = 25'b0000000000000000000000000;
    rom[117] = 25'b0000000000000000000000000;
    rom[118] = 25'b0000000000000000000000000;
    rom[119] = 25'b0000000000000000000000000;
    rom[120] = 25'b0000000000000000000000000;
    rom[121] = 25'b0000000000000000000000000;
    rom[122] = 25'b0000000000000000000000000;
    rom[123] = 25'b0000000000000000000000000;
    rom[124] = 25'b0000000000000000000000000;
    rom[125] = 25'b0000000000000000000000000;
    rom[126] = 25'b0000000000000000000000000;
    rom[127] = 25'b0000000000000000000000000;
end

// port a
always @(posedge clk)
begin
    if (wea_d == 1'b1) begin
      rom[addra_d] <= dia_d;
    end
    wea_d <= wea;
    dia_d <= dia;
    addra_d <= addra;
end

// port b
always @(posedge clk)
begin
    addrb_d <= addrb;
    rom_pipea <= rom[addrb_d];
    dob_d <= rom_pipea;
end

endmodule
