
//     Licensed to the Apache Software Foundation (ASF) under one
// or more contributor license agreements.  See the NOTICE file
// distributed with this work for additional information
// regarding copyright ownership.  The ASF licenses this file
// to you under the Apache License, Version 2.0 (the
// "License"); you may not use this file except in compliance
// with the License.  You may obtain a copy of the License at
// 
//   http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing,
// software distributed under the License is distributed on an
// "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY
// KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations
// under the License.  


/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : pfb_2048Mmax_16iw_16ow_32tps_dp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data                                                     
//
//
/*****************************************************************************/


module pfb_2048Mmax_16iw_16ow_32tps_dp_rom
(
  input clk, 
  input wea,
  input [24:0] dia,
  input [15:0] addra,
  input [15:0] addrb,
  output [24:0] dob
);

(* rom_style = "block" *) reg [24:0] rom [65535:0];
reg [15:0] addrb_d;
reg [24:0] dob_d;
reg [24:0] rom_pipea;
reg [15:0] addra_d;
reg [24:0] dia_d;
reg wea_d;

assign dob = dob_d;

initial
begin
    rom[0] = 25'b1111111111111111110011100;
    rom[1] = 25'b1111111111111111110011100;
    rom[2] = 25'b1111111111111111110011100;
    rom[3] = 25'b1111111111111111110011100;
    rom[4] = 25'b1111111111111111110011100;
    rom[5] = 25'b1111111111111111110011100;
    rom[6] = 25'b1111111111111111110011100;
    rom[7] = 25'b1111111111111111110011100;
    rom[8] = 25'b1111111111111111110011100;
    rom[9] = 25'b1111111111111111110011100;
    rom[10] = 25'b1111111111111111110011100;
    rom[11] = 25'b1111111111111111110011100;
    rom[12] = 25'b1111111111111111110011100;
    rom[13] = 25'b1111111111111111110011100;
    rom[14] = 25'b1111111111111111110011100;
    rom[15] = 25'b1111111111111111110011100;
    rom[16] = 25'b1111111111111111110011100;
    rom[17] = 25'b1111111111111111110011100;
    rom[18] = 25'b1111111111111111110011100;
    rom[19] = 25'b1111111111111111110011100;
    rom[20] = 25'b1111111111111111110011100;
    rom[21] = 25'b1111111111111111110011100;
    rom[22] = 25'b1111111111111111110011100;
    rom[23] = 25'b1111111111111111110011100;
    rom[24] = 25'b1111111111111111110011100;
    rom[25] = 25'b1111111111111111110011100;
    rom[26] = 25'b1111111111111111110011100;
    rom[27] = 25'b1111111111111111110011100;
    rom[28] = 25'b1111111111111111110011100;
    rom[29] = 25'b1111111111111111110011100;
    rom[30] = 25'b1111111111111111110011100;
    rom[31] = 25'b1111111111111111110011100;
    rom[32] = 25'b1111111111111111110011100;
    rom[33] = 25'b1111111111111111110011100;
    rom[34] = 25'b1111111111111111110011100;
    rom[35] = 25'b1111111111111111110011100;
    rom[36] = 25'b1111111111111111110011100;
    rom[37] = 25'b1111111111111111110011100;
    rom[38] = 25'b1111111111111111110011100;
    rom[39] = 25'b1111111111111111110011100;
    rom[40] = 25'b1111111111111111110011100;
    rom[41] = 25'b1111111111111111110011100;
    rom[42] = 25'b1111111111111111110011100;
    rom[43] = 25'b1111111111111111110011100;
    rom[44] = 25'b1111111111111111110011011;
    rom[45] = 25'b1111111111111111110011011;
    rom[46] = 25'b1111111111111111110011011;
    rom[47] = 25'b1111111111111111110011011;
    rom[48] = 25'b1111111111111111110011011;
    rom[49] = 25'b1111111111111111110011011;
    rom[50] = 25'b1111111111111111110011011;
    rom[51] = 25'b1111111111111111110011011;
    rom[52] = 25'b1111111111111111110011011;
    rom[53] = 25'b1111111111111111110011011;
    rom[54] = 25'b1111111111111111110011011;
    rom[55] = 25'b1111111111111111110011011;
    rom[56] = 25'b1111111111111111110011011;
    rom[57] = 25'b1111111111111111110011011;
    rom[58] = 25'b1111111111111111110011011;
    rom[59] = 25'b1111111111111111110011011;
    rom[60] = 25'b1111111111111111110011011;
    rom[61] = 25'b1111111111111111110011011;
    rom[62] = 25'b1111111111111111110011011;
    rom[63] = 25'b1111111111111111110011011;
    rom[64] = 25'b1111111111111111110011011;
    rom[65] = 25'b1111111111111111110011011;
    rom[66] = 25'b1111111111111111110011011;
    rom[67] = 25'b1111111111111111110011011;
    rom[68] = 25'b1111111111111111110011011;
    rom[69] = 25'b1111111111111111110011011;
    rom[70] = 25'b1111111111111111110011011;
    rom[71] = 25'b1111111111111111110011011;
    rom[72] = 25'b1111111111111111110011011;
    rom[73] = 25'b1111111111111111110011011;
    rom[74] = 25'b1111111111111111110011011;
    rom[75] = 25'b1111111111111111110011011;
    rom[76] = 25'b1111111111111111110011011;
    rom[77] = 25'b1111111111111111110011011;
    rom[78] = 25'b1111111111111111110011011;
    rom[79] = 25'b1111111111111111110011011;
    rom[80] = 25'b1111111111111111110011011;
    rom[81] = 25'b1111111111111111110011011;
    rom[82] = 25'b1111111111111111110011011;
    rom[83] = 25'b1111111111111111110011011;
    rom[84] = 25'b1111111111111111110011010;
    rom[85] = 25'b1111111111111111110011010;
    rom[86] = 25'b1111111111111111110011010;
    rom[87] = 25'b1111111111111111110011010;
    rom[88] = 25'b1111111111111111110011010;
    rom[89] = 25'b1111111111111111110011010;
    rom[90] = 25'b1111111111111111110011010;
    rom[91] = 25'b1111111111111111110011010;
    rom[92] = 25'b1111111111111111110011010;
    rom[93] = 25'b1111111111111111110011010;
    rom[94] = 25'b1111111111111111110011010;
    rom[95] = 25'b1111111111111111110011010;
    rom[96] = 25'b1111111111111111110011010;
    rom[97] = 25'b1111111111111111110011010;
    rom[98] = 25'b1111111111111111110011001;
    rom[99] = 25'b1111111111111111110011001;
    rom[100] = 25'b1111111111111111110011001;
    rom[101] = 25'b1111111111111111110011001;
    rom[102] = 25'b1111111111111111110011001;
    rom[103] = 25'b1111111111111111110011001;
    rom[104] = 25'b1111111111111111110011001;
    rom[105] = 25'b1111111111111111110011001;
    rom[106] = 25'b1111111111111111110011001;
    rom[107] = 25'b1111111111111111110011001;
    rom[108] = 25'b1111111111111111110011001;
    rom[109] = 25'b1111111111111111110011001;
    rom[110] = 25'b1111111111111111110011000;
    rom[111] = 25'b1111111111111111110011000;
    rom[112] = 25'b1111111111111111110011000;
    rom[113] = 25'b1111111111111111110011000;
    rom[114] = 25'b1111111111111111110011000;
    rom[115] = 25'b1111111111111111110011000;
    rom[116] = 25'b1111111111111111110011000;
    rom[117] = 25'b1111111111111111110011000;
    rom[118] = 25'b1111111111111111110011000;
    rom[119] = 25'b1111111111111111110011000;
    rom[120] = 25'b1111111111111111110011000;
    rom[121] = 25'b1111111111111111110011000;
    rom[122] = 25'b1111111111111111110011000;
    rom[123] = 25'b1111111111111111110011000;
    rom[124] = 25'b1111111111111111110011000;
    rom[125] = 25'b1111111111111111110011000;
    rom[126] = 25'b1111111111111111110011000;
    rom[127] = 25'b1111111111111111110011000;
    rom[128] = 25'b1111111111111111110011000;
    rom[129] = 25'b1111111111111111110011000;
    rom[130] = 25'b1111111111111111110011000;
    rom[131] = 25'b1111111111111111110011000;
    rom[132] = 25'b1111111111111111110010111;
    rom[133] = 25'b1111111111111111110010111;
    rom[134] = 25'b1111111111111111110010111;
    rom[135] = 25'b1111111111111111110010111;
    rom[136] = 25'b1111111111111111110010111;
    rom[137] = 25'b1111111111111111110010111;
    rom[138] = 25'b1111111111111111110010111;
    rom[139] = 25'b1111111111111111110010111;
    rom[140] = 25'b1111111111111111110010111;
    rom[141] = 25'b1111111111111111110010110;
    rom[142] = 25'b1111111111111111110010110;
    rom[143] = 25'b1111111111111111110010110;
    rom[144] = 25'b1111111111111111110010110;
    rom[145] = 25'b1111111111111111110010110;
    rom[146] = 25'b1111111111111111110010110;
    rom[147] = 25'b1111111111111111110010110;
    rom[148] = 25'b1111111111111111110010110;
    rom[149] = 25'b1111111111111111110010110;
    rom[150] = 25'b1111111111111111110010101;
    rom[151] = 25'b1111111111111111110010101;
    rom[152] = 25'b1111111111111111110010101;
    rom[153] = 25'b1111111111111111110010101;
    rom[154] = 25'b1111111111111111110010101;
    rom[155] = 25'b1111111111111111110010101;
    rom[156] = 25'b1111111111111111110010101;
    rom[157] = 25'b1111111111111111110010101;
    rom[158] = 25'b1111111111111111110010101;
    rom[159] = 25'b1111111111111111110010101;
    rom[160] = 25'b1111111111111111110010101;
    rom[161] = 25'b1111111111111111110010101;
    rom[162] = 25'b1111111111111111110010101;
    rom[163] = 25'b1111111111111111110010101;
    rom[164] = 25'b1111111111111111110010101;
    rom[165] = 25'b1111111111111111110010101;
    rom[166] = 25'b1111111111111111110010100;
    rom[167] = 25'b1111111111111111110010100;
    rom[168] = 25'b1111111111111111110010100;
    rom[169] = 25'b1111111111111111110010100;
    rom[170] = 25'b1111111111111111110010100;
    rom[171] = 25'b1111111111111111110010100;
    rom[172] = 25'b1111111111111111110010100;
    rom[173] = 25'b1111111111111111110010100;
    rom[174] = 25'b1111111111111111110010011;
    rom[175] = 25'b1111111111111111110010011;
    rom[176] = 25'b1111111111111111110010011;
    rom[177] = 25'b1111111111111111110010011;
    rom[178] = 25'b1111111111111111110010011;
    rom[179] = 25'b1111111111111111110010011;
    rom[180] = 25'b1111111111111111110010011;
    rom[181] = 25'b1111111111111111110010010;
    rom[182] = 25'b1111111111111111110010010;
    rom[183] = 25'b1111111111111111110010010;
    rom[184] = 25'b1111111111111111110010010;
    rom[185] = 25'b1111111111111111110010010;
    rom[186] = 25'b1111111111111111110010010;
    rom[187] = 25'b1111111111111111110010010;
    rom[188] = 25'b1111111111111111110010010;
    rom[189] = 25'b1111111111111111110010010;
    rom[190] = 25'b1111111111111111110010010;
    rom[191] = 25'b1111111111111111110010010;
    rom[192] = 25'b1111111111111111110010010;
    rom[193] = 25'b1111111111111111110010010;
    rom[194] = 25'b1111111111111111110010010;
    rom[195] = 25'b1111111111111111110010001;
    rom[196] = 25'b1111111111111111110010001;
    rom[197] = 25'b1111111111111111110010001;
    rom[198] = 25'b1111111111111111110010001;
    rom[199] = 25'b1111111111111111110010001;
    rom[200] = 25'b1111111111111111110010001;
    rom[201] = 25'b1111111111111111110010001;
    rom[202] = 25'b1111111111111111110010000;
    rom[203] = 25'b1111111111111111110010000;
    rom[204] = 25'b1111111111111111110010000;
    rom[205] = 25'b1111111111111111110010000;
    rom[206] = 25'b1111111111111111110010000;
    rom[207] = 25'b1111111111111111110010000;
    rom[208] = 25'b1111111111111111110001111;
    rom[209] = 25'b1111111111111111110001111;
    rom[210] = 25'b1111111111111111110001111;
    rom[211] = 25'b1111111111111111110001111;
    rom[212] = 25'b1111111111111111110001111;
    rom[213] = 25'b1111111111111111110001111;
    rom[214] = 25'b1111111111111111110001111;
    rom[215] = 25'b1111111111111111110001111;
    rom[216] = 25'b1111111111111111110001111;
    rom[217] = 25'b1111111111111111110001111;
    rom[218] = 25'b1111111111111111110001111;
    rom[219] = 25'b1111111111111111110001111;
    rom[220] = 25'b1111111111111111110001110;
    rom[221] = 25'b1111111111111111110001110;
    rom[222] = 25'b1111111111111111110001110;
    rom[223] = 25'b1111111111111111110001110;
    rom[224] = 25'b1111111111111111110001110;
    rom[225] = 25'b1111111111111111110001110;
    rom[226] = 25'b1111111111111111110001101;
    rom[227] = 25'b1111111111111111110001101;
    rom[228] = 25'b1111111111111111110001101;
    rom[229] = 25'b1111111111111111110001101;
    rom[230] = 25'b1111111111111111110001101;
    rom[231] = 25'b1111111111111111110001101;
    rom[232] = 25'b1111111111111111110001100;
    rom[233] = 25'b1111111111111111110001100;
    rom[234] = 25'b1111111111111111110001100;
    rom[235] = 25'b1111111111111111110001100;
    rom[236] = 25'b1111111111111111110001100;
    rom[237] = 25'b1111111111111111110001100;
    rom[238] = 25'b1111111111111111110001100;
    rom[239] = 25'b1111111111111111110001100;
    rom[240] = 25'b1111111111111111110001100;
    rom[241] = 25'b1111111111111111110001100;
    rom[242] = 25'b1111111111111111110001100;
    rom[243] = 25'b1111111111111111110001011;
    rom[244] = 25'b1111111111111111110001011;
    rom[245] = 25'b1111111111111111110001011;
    rom[246] = 25'b1111111111111111110001011;
    rom[247] = 25'b1111111111111111110001011;
    rom[248] = 25'b1111111111111111110001010;
    rom[249] = 25'b1111111111111111110001010;
    rom[250] = 25'b1111111111111111110001010;
    rom[251] = 25'b1111111111111111110001010;
    rom[252] = 25'b1111111111111111110001010;
    rom[253] = 25'b1111111111111111110001001;
    rom[254] = 25'b1111111111111111110001001;
    rom[255] = 25'b1111111111111111110001001;
    rom[256] = 25'b1111111111111111110001001;
    rom[257] = 25'b1111111111111111110001001;
    rom[258] = 25'b1111111111111111110001001;
    rom[259] = 25'b1111111111111111110001001;
    rom[260] = 25'b1111111111111111110001001;
    rom[261] = 25'b1111111111111111110001001;
    rom[262] = 25'b1111111111111111110001001;
    rom[263] = 25'b1111111111111111110001000;
    rom[264] = 25'b1111111111111111110001000;
    rom[265] = 25'b1111111111111111110001000;
    rom[266] = 25'b1111111111111111110001000;
    rom[267] = 25'b1111111111111111110001000;
    rom[268] = 25'b1111111111111111110000111;
    rom[269] = 25'b1111111111111111110000111;
    rom[270] = 25'b1111111111111111110000111;
    rom[271] = 25'b1111111111111111110000111;
    rom[272] = 25'b1111111111111111110000111;
    rom[273] = 25'b1111111111111111110000110;
    rom[274] = 25'b1111111111111111110000110;
    rom[275] = 25'b1111111111111111110000110;
    rom[276] = 25'b1111111111111111110000110;
    rom[277] = 25'b1111111111111111110000110;
    rom[278] = 25'b1111111111111111110000110;
    rom[279] = 25'b1111111111111111110000110;
    rom[280] = 25'b1111111111111111110000110;
    rom[281] = 25'b1111111111111111110000110;
    rom[282] = 25'b1111111111111111110000110;
    rom[283] = 25'b1111111111111111110000101;
    rom[284] = 25'b1111111111111111110000101;
    rom[285] = 25'b1111111111111111110000101;
    rom[286] = 25'b1111111111111111110000101;
    rom[287] = 25'b1111111111111111110000100;
    rom[288] = 25'b1111111111111111110000100;
    rom[289] = 25'b1111111111111111110000100;
    rom[290] = 25'b1111111111111111110000100;
    rom[291] = 25'b1111111111111111110000100;
    rom[292] = 25'b1111111111111111110000011;
    rom[293] = 25'b1111111111111111110000011;
    rom[294] = 25'b1111111111111111110000011;
    rom[295] = 25'b1111111111111111110000011;
    rom[296] = 25'b1111111111111111110000011;
    rom[297] = 25'b1111111111111111110000011;
    rom[298] = 25'b1111111111111111110000011;
    rom[299] = 25'b1111111111111111110000011;
    rom[300] = 25'b1111111111111111110000011;
    rom[301] = 25'b1111111111111111110000010;
    rom[302] = 25'b1111111111111111110000010;
    rom[303] = 25'b1111111111111111110000010;
    rom[304] = 25'b1111111111111111110000010;
    rom[305] = 25'b1111111111111111110000001;
    rom[306] = 25'b1111111111111111110000001;
    rom[307] = 25'b1111111111111111110000001;
    rom[308] = 25'b1111111111111111110000001;
    rom[309] = 25'b1111111111111111110000001;
    rom[310] = 25'b1111111111111111110000000;
    rom[311] = 25'b1111111111111111110000000;
    rom[312] = 25'b1111111111111111110000000;
    rom[313] = 25'b1111111111111111110000000;
    rom[314] = 25'b1111111111111111110000000;
    rom[315] = 25'b1111111111111111110000000;
    rom[316] = 25'b1111111111111111110000000;
    rom[317] = 25'b1111111111111111110000000;
    rom[318] = 25'b1111111111111111101111111;
    rom[319] = 25'b1111111111111111101111111;
    rom[320] = 25'b1111111111111111101111111;
    rom[321] = 25'b1111111111111111101111111;
    rom[322] = 25'b1111111111111111101111110;
    rom[323] = 25'b1111111111111111101111110;
    rom[324] = 25'b1111111111111111101111110;
    rom[325] = 25'b1111111111111111101111110;
    rom[326] = 25'b1111111111111111101111110;
    rom[327] = 25'b1111111111111111101111110;
    rom[328] = 25'b1111111111111111101111110;
    rom[329] = 25'b1111111111111111101111110;
    rom[330] = 25'b1111111111111111101111101;
    rom[331] = 25'b1111111111111111101111101;
    rom[332] = 25'b1111111111111111101111101;
    rom[333] = 25'b1111111111111111101111101;
    rom[334] = 25'b1111111111111111101111101;
    rom[335] = 25'b1111111111111111101111100;
    rom[336] = 25'b1111111111111111101111100;
    rom[337] = 25'b1111111111111111101111100;
    rom[338] = 25'b1111111111111111101111011;
    rom[339] = 25'b1111111111111111101111011;
    rom[340] = 25'b1111111111111111101111011;
    rom[341] = 25'b1111111111111111101111011;
    rom[342] = 25'b1111111111111111101111011;
    rom[343] = 25'b1111111111111111101111011;
    rom[344] = 25'b1111111111111111101111011;
    rom[345] = 25'b1111111111111111101111011;
    rom[346] = 25'b1111111111111111101111010;
    rom[347] = 25'b1111111111111111101111010;
    rom[348] = 25'b1111111111111111101111010;
    rom[349] = 25'b1111111111111111101111010;
    rom[350] = 25'b1111111111111111101111001;
    rom[351] = 25'b1111111111111111101111001;
    rom[352] = 25'b1111111111111111101111001;
    rom[353] = 25'b1111111111111111101111001;
    rom[354] = 25'b1111111111111111101111000;
    rom[355] = 25'b1111111111111111101111000;
    rom[356] = 25'b1111111111111111101111000;
    rom[357] = 25'b1111111111111111101111000;
    rom[358] = 25'b1111111111111111101111000;
    rom[359] = 25'b1111111111111111101111000;
    rom[360] = 25'b1111111111111111101111000;
    rom[361] = 25'b1111111111111111101111000;
    rom[362] = 25'b1111111111111111101110111;
    rom[363] = 25'b1111111111111111101110111;
    rom[364] = 25'b1111111111111111101110111;
    rom[365] = 25'b1111111111111111101110110;
    rom[366] = 25'b1111111111111111101110110;
    rom[367] = 25'b1111111111111111101110110;
    rom[368] = 25'b1111111111111111101110110;
    rom[369] = 25'b1111111111111111101110101;
    rom[370] = 25'b1111111111111111101110101;
    rom[371] = 25'b1111111111111111101110101;
    rom[372] = 25'b1111111111111111101110101;
    rom[373] = 25'b1111111111111111101110101;
    rom[374] = 25'b1111111111111111101110101;
    rom[375] = 25'b1111111111111111101110101;
    rom[376] = 25'b1111111111111111101110100;
    rom[377] = 25'b1111111111111111101110100;
    rom[378] = 25'b1111111111111111101110100;
    rom[379] = 25'b1111111111111111101110100;
    rom[380] = 25'b1111111111111111101110011;
    rom[381] = 25'b1111111111111111101110011;
    rom[382] = 25'b1111111111111111101110011;
    rom[383] = 25'b1111111111111111101110010;
    rom[384] = 25'b1111111111111111101110010;
    rom[385] = 25'b1111111111111111101110010;
    rom[386] = 25'b1111111111111111101110010;
    rom[387] = 25'b1111111111111111101110010;
    rom[388] = 25'b1111111111111111101110010;
    rom[389] = 25'b1111111111111111101110010;
    rom[390] = 25'b1111111111111111101110010;
    rom[391] = 25'b1111111111111111101110001;
    rom[392] = 25'b1111111111111111101110001;
    rom[393] = 25'b1111111111111111101110001;
    rom[394] = 25'b1111111111111111101110000;
    rom[395] = 25'b1111111111111111101110000;
    rom[396] = 25'b1111111111111111101110000;
    rom[397] = 25'b1111111111111111101101111;
    rom[398] = 25'b1111111111111111101101111;
    rom[399] = 25'b1111111111111111101101111;
    rom[400] = 25'b1111111111111111101101111;
    rom[401] = 25'b1111111111111111101101111;
    rom[402] = 25'b1111111111111111101101111;
    rom[403] = 25'b1111111111111111101101111;
    rom[404] = 25'b1111111111111111101101110;
    rom[405] = 25'b1111111111111111101101110;
    rom[406] = 25'b1111111111111111101101110;
    rom[407] = 25'b1111111111111111101101110;
    rom[408] = 25'b1111111111111111101101101;
    rom[409] = 25'b1111111111111111101101101;
    rom[410] = 25'b1111111111111111101101101;
    rom[411] = 25'b1111111111111111101101100;
    rom[412] = 25'b1111111111111111101101100;
    rom[413] = 25'b1111111111111111101101100;
    rom[414] = 25'b1111111111111111101101100;
    rom[415] = 25'b1111111111111111101101100;
    rom[416] = 25'b1111111111111111101101100;
    rom[417] = 25'b1111111111111111101101100;
    rom[418] = 25'b1111111111111111101101011;
    rom[419] = 25'b1111111111111111101101011;
    rom[420] = 25'b1111111111111111101101011;
    rom[421] = 25'b1111111111111111101101010;
    rom[422] = 25'b1111111111111111101101010;
    rom[423] = 25'b1111111111111111101101010;
    rom[424] = 25'b1111111111111111101101001;
    rom[425] = 25'b1111111111111111101101001;
    rom[426] = 25'b1111111111111111101101001;
    rom[427] = 25'b1111111111111111101101001;
    rom[428] = 25'b1111111111111111101101001;
    rom[429] = 25'b1111111111111111101101001;
    rom[430] = 25'b1111111111111111101101001;
    rom[431] = 25'b1111111111111111101101000;
    rom[432] = 25'b1111111111111111101101000;
    rom[433] = 25'b1111111111111111101101000;
    rom[434] = 25'b1111111111111111101100111;
    rom[435] = 25'b1111111111111111101100111;
    rom[436] = 25'b1111111111111111101100111;
    rom[437] = 25'b1111111111111111101100110;
    rom[438] = 25'b1111111111111111101100110;
    rom[439] = 25'b1111111111111111101100110;
    rom[440] = 25'b1111111111111111101100110;
    rom[441] = 25'b1111111111111111101100110;
    rom[442] = 25'b1111111111111111101100110;
    rom[443] = 25'b1111111111111111101100101;
    rom[444] = 25'b1111111111111111101100101;
    rom[445] = 25'b1111111111111111101100101;
    rom[446] = 25'b1111111111111111101100101;
    rom[447] = 25'b1111111111111111101100100;
    rom[448] = 25'b1111111111111111101100100;
    rom[449] = 25'b1111111111111111101100100;
    rom[450] = 25'b1111111111111111101100011;
    rom[451] = 25'b1111111111111111101100011;
    rom[452] = 25'b1111111111111111101100011;
    rom[453] = 25'b1111111111111111101100011;
    rom[454] = 25'b1111111111111111101100011;
    rom[455] = 25'b1111111111111111101100011;
    rom[456] = 25'b1111111111111111101100010;
    rom[457] = 25'b1111111111111111101100010;
    rom[458] = 25'b1111111111111111101100010;
    rom[459] = 25'b1111111111111111101100001;
    rom[460] = 25'b1111111111111111101100001;
    rom[461] = 25'b1111111111111111101100001;
    rom[462] = 25'b1111111111111111101100000;
    rom[463] = 25'b1111111111111111101100000;
    rom[464] = 25'b1111111111111111101100000;
    rom[465] = 25'b1111111111111111101100000;
    rom[466] = 25'b1111111111111111101100000;
    rom[467] = 25'b1111111111111111101100000;
    rom[468] = 25'b1111111111111111101011111;
    rom[469] = 25'b1111111111111111101011111;
    rom[470] = 25'b1111111111111111101011111;
    rom[471] = 25'b1111111111111111101011110;
    rom[472] = 25'b1111111111111111101011110;
    rom[473] = 25'b1111111111111111101011110;
    rom[474] = 25'b1111111111111111101011101;
    rom[475] = 25'b1111111111111111101011101;
    rom[476] = 25'b1111111111111111101011101;
    rom[477] = 25'b1111111111111111101011101;
    rom[478] = 25'b1111111111111111101011101;
    rom[479] = 25'b1111111111111111101011101;
    rom[480] = 25'b1111111111111111101011100;
    rom[481] = 25'b1111111111111111101011100;
    rom[482] = 25'b1111111111111111101011100;
    rom[483] = 25'b1111111111111111101011011;
    rom[484] = 25'b1111111111111111101011011;
    rom[485] = 25'b1111111111111111101011011;
    rom[486] = 25'b1111111111111111101011010;
    rom[487] = 25'b1111111111111111101011010;
    rom[488] = 25'b1111111111111111101011010;
    rom[489] = 25'b1111111111111111101011010;
    rom[490] = 25'b1111111111111111101011010;
    rom[491] = 25'b1111111111111111101011010;
    rom[492] = 25'b1111111111111111101011001;
    rom[493] = 25'b1111111111111111101011001;
    rom[494] = 25'b1111111111111111101011001;
    rom[495] = 25'b1111111111111111101011000;
    rom[496] = 25'b1111111111111111101011000;
    rom[497] = 25'b1111111111111111101011000;
    rom[498] = 25'b1111111111111111101010111;
    rom[499] = 25'b1111111111111111101010111;
    rom[500] = 25'b1111111111111111101010111;
    rom[501] = 25'b1111111111111111101010111;
    rom[502] = 25'b1111111111111111101010111;
    rom[503] = 25'b1111111111111111101010110;
    rom[504] = 25'b1111111111111111101010110;
    rom[505] = 25'b1111111111111111101010110;
    rom[506] = 25'b1111111111111111101010101;
    rom[507] = 25'b1111111111111111101010101;
    rom[508] = 25'b1111111111111111101010101;
    rom[509] = 25'b1111111111111111101010100;
    rom[510] = 25'b1111111111111111101010100;
    rom[511] = 25'b1111111111111111101010100;
    rom[512] = 25'b1111111111111111101010100;
    rom[513] = 25'b1111111111111111101010100;
    rom[514] = 25'b1111111111111111101010100;
    rom[515] = 25'b1111111111111111101010011;
    rom[516] = 25'b1111111111111111101010011;
    rom[517] = 25'b1111111111111111101010010;
    rom[518] = 25'b1111111111111111101010010;
    rom[519] = 25'b1111111111111111101010010;
    rom[520] = 25'b1111111111111111101010001;
    rom[521] = 25'b1111111111111111101010001;
    rom[522] = 25'b1111111111111111101010001;
    rom[523] = 25'b1111111111111111101010001;
    rom[524] = 25'b1111111111111111101010001;
    rom[525] = 25'b1111111111111111101010001;
    rom[526] = 25'b1111111111111111101010000;
    rom[527] = 25'b1111111111111111101010000;
    rom[528] = 25'b1111111111111111101001111;
    rom[529] = 25'b1111111111111111101001111;
    rom[530] = 25'b1111111111111111101001111;
    rom[531] = 25'b1111111111111111101001110;
    rom[532] = 25'b1111111111111111101001110;
    rom[533] = 25'b1111111111111111101001110;
    rom[534] = 25'b1111111111111111101001110;
    rom[535] = 25'b1111111111111111101001110;
    rom[536] = 25'b1111111111111111101001110;
    rom[537] = 25'b1111111111111111101001101;
    rom[538] = 25'b1111111111111111101001101;
    rom[539] = 25'b1111111111111111101001100;
    rom[540] = 25'b1111111111111111101001100;
    rom[541] = 25'b1111111111111111101001100;
    rom[542] = 25'b1111111111111111101001011;
    rom[543] = 25'b1111111111111111101001011;
    rom[544] = 25'b1111111111111111101001011;
    rom[545] = 25'b1111111111111111101001011;
    rom[546] = 25'b1111111111111111101001011;
    rom[547] = 25'b1111111111111111101001010;
    rom[548] = 25'b1111111111111111101001010;
    rom[549] = 25'b1111111111111111101001010;
    rom[550] = 25'b1111111111111111101001001;
    rom[551] = 25'b1111111111111111101001001;
    rom[552] = 25'b1111111111111111101001001;
    rom[553] = 25'b1111111111111111101001000;
    rom[554] = 25'b1111111111111111101001000;
    rom[555] = 25'b1111111111111111101001000;
    rom[556] = 25'b1111111111111111101001000;
    rom[557] = 25'b1111111111111111101001000;
    rom[558] = 25'b1111111111111111101000111;
    rom[559] = 25'b1111111111111111101000111;
    rom[560] = 25'b1111111111111111101000111;
    rom[561] = 25'b1111111111111111101000110;
    rom[562] = 25'b1111111111111111101000110;
    rom[563] = 25'b1111111111111111101000101;
    rom[564] = 25'b1111111111111111101000101;
    rom[565] = 25'b1111111111111111101000101;
    rom[566] = 25'b1111111111111111101000101;
    rom[567] = 25'b1111111111111111101000101;
    rom[568] = 25'b1111111111111111101000101;
    rom[569] = 25'b1111111111111111101000100;
    rom[570] = 25'b1111111111111111101000100;
    rom[571] = 25'b1111111111111111101000011;
    rom[572] = 25'b1111111111111111101000011;
    rom[573] = 25'b1111111111111111101000011;
    rom[574] = 25'b1111111111111111101000010;
    rom[575] = 25'b1111111111111111101000010;
    rom[576] = 25'b1111111111111111101000010;
    rom[577] = 25'b1111111111111111101000010;
    rom[578] = 25'b1111111111111111101000010;
    rom[579] = 25'b1111111111111111101000001;
    rom[580] = 25'b1111111111111111101000001;
    rom[581] = 25'b1111111111111111101000000;
    rom[582] = 25'b1111111111111111101000000;
    rom[583] = 25'b1111111111111111101000000;
    rom[584] = 25'b1111111111111111100111111;
    rom[585] = 25'b1111111111111111100111111;
    rom[586] = 25'b1111111111111111100111111;
    rom[587] = 25'b1111111111111111100111111;
    rom[588] = 25'b1111111111111111100111111;
    rom[589] = 25'b1111111111111111100111110;
    rom[590] = 25'b1111111111111111100111110;
    rom[591] = 25'b1111111111111111100111110;
    rom[592] = 25'b1111111111111111100111101;
    rom[593] = 25'b1111111111111111100111101;
    rom[594] = 25'b1111111111111111100111101;
    rom[595] = 25'b1111111111111111100111101;
    rom[596] = 25'b1111111111111111100111101;
    rom[597] = 25'b1111111111111111100111100;
    rom[598] = 25'b1111111111111111100111100;
    rom[599] = 25'b1111111111111111100111011;
    rom[600] = 25'b1111111111111111100111011;
    rom[601] = 25'b1111111111111111100111011;
    rom[602] = 25'b1111111111111111100111010;
    rom[603] = 25'b1111111111111111100111010;
    rom[604] = 25'b1111111111111111100111010;
    rom[605] = 25'b1111111111111111100111010;
    rom[606] = 25'b1111111111111111100111010;
    rom[607] = 25'b1111111111111111100111001;
    rom[608] = 25'b1111111111111111100111001;
    rom[609] = 25'b1111111111111111100111000;
    rom[610] = 25'b1111111111111111100111000;
    rom[611] = 25'b1111111111111111100111000;
    rom[612] = 25'b1111111111111111100110111;
    rom[613] = 25'b1111111111111111100110111;
    rom[614] = 25'b1111111111111111100110111;
    rom[615] = 25'b1111111111111111100110111;
    rom[616] = 25'b1111111111111111100110111;
    rom[617] = 25'b1111111111111111100110110;
    rom[618] = 25'b1111111111111111100110110;
    rom[619] = 25'b1111111111111111100110101;
    rom[620] = 25'b1111111111111111100110101;
    rom[621] = 25'b1111111111111111100110101;
    rom[622] = 25'b1111111111111111100110100;
    rom[623] = 25'b1111111111111111100110100;
    rom[624] = 25'b1111111111111111100110100;
    rom[625] = 25'b1111111111111111100110100;
    rom[626] = 25'b1111111111111111100110100;
    rom[627] = 25'b1111111111111111100110011;
    rom[628] = 25'b1111111111111111100110011;
    rom[629] = 25'b1111111111111111100110010;
    rom[630] = 25'b1111111111111111100110010;
    rom[631] = 25'b1111111111111111100110001;
    rom[632] = 25'b1111111111111111100110001;
    rom[633] = 25'b1111111111111111100110001;
    rom[634] = 25'b1111111111111111100110001;
    rom[635] = 25'b1111111111111111100110001;
    rom[636] = 25'b1111111111111111100110000;
    rom[637] = 25'b1111111111111111100110000;
    rom[638] = 25'b1111111111111111100110000;
    rom[639] = 25'b1111111111111111100101111;
    rom[640] = 25'b1111111111111111100101111;
    rom[641] = 25'b1111111111111111100101110;
    rom[642] = 25'b1111111111111111100101110;
    rom[643] = 25'b1111111111111111100101110;
    rom[644] = 25'b1111111111111111100101110;
    rom[645] = 25'b1111111111111111100101110;
    rom[646] = 25'b1111111111111111100101101;
    rom[647] = 25'b1111111111111111100101101;
    rom[648] = 25'b1111111111111111100101100;
    rom[649] = 25'b1111111111111111100101100;
    rom[650] = 25'b1111111111111111100101100;
    rom[651] = 25'b1111111111111111100101011;
    rom[652] = 25'b1111111111111111100101011;
    rom[653] = 25'b1111111111111111100101011;
    rom[654] = 25'b1111111111111111100101011;
    rom[655] = 25'b1111111111111111100101011;
    rom[656] = 25'b1111111111111111100101010;
    rom[657] = 25'b1111111111111111100101010;
    rom[658] = 25'b1111111111111111100101001;
    rom[659] = 25'b1111111111111111100101001;
    rom[660] = 25'b1111111111111111100101000;
    rom[661] = 25'b1111111111111111100101000;
    rom[662] = 25'b1111111111111111100101000;
    rom[663] = 25'b1111111111111111100101000;
    rom[664] = 25'b1111111111111111100101000;
    rom[665] = 25'b1111111111111111100100111;
    rom[666] = 25'b1111111111111111100100111;
    rom[667] = 25'b1111111111111111100100110;
    rom[668] = 25'b1111111111111111100100110;
    rom[669] = 25'b1111111111111111100100110;
    rom[670] = 25'b1111111111111111100100101;
    rom[671] = 25'b1111111111111111100100101;
    rom[672] = 25'b1111111111111111100100101;
    rom[673] = 25'b1111111111111111100100101;
    rom[674] = 25'b1111111111111111100100101;
    rom[675] = 25'b1111111111111111100100100;
    rom[676] = 25'b1111111111111111100100100;
    rom[677] = 25'b1111111111111111100100011;
    rom[678] = 25'b1111111111111111100100011;
    rom[679] = 25'b1111111111111111100100010;
    rom[680] = 25'b1111111111111111100100010;
    rom[681] = 25'b1111111111111111100100010;
    rom[682] = 25'b1111111111111111100100010;
    rom[683] = 25'b1111111111111111100100010;
    rom[684] = 25'b1111111111111111100100001;
    rom[685] = 25'b1111111111111111100100001;
    rom[686] = 25'b1111111111111111100100000;
    rom[687] = 25'b1111111111111111100100000;
    rom[688] = 25'b1111111111111111100100000;
    rom[689] = 25'b1111111111111111100011111;
    rom[690] = 25'b1111111111111111100011111;
    rom[691] = 25'b1111111111111111100011111;
    rom[692] = 25'b1111111111111111100011111;
    rom[693] = 25'b1111111111111111100011110;
    rom[694] = 25'b1111111111111111100011110;
    rom[695] = 25'b1111111111111111100011110;
    rom[696] = 25'b1111111111111111100011101;
    rom[697] = 25'b1111111111111111100011101;
    rom[698] = 25'b1111111111111111100011100;
    rom[699] = 25'b1111111111111111100011100;
    rom[700] = 25'b1111111111111111100011100;
    rom[701] = 25'b1111111111111111100011100;
    rom[702] = 25'b1111111111111111100011011;
    rom[703] = 25'b1111111111111111100011011;
    rom[704] = 25'b1111111111111111100011011;
    rom[705] = 25'b1111111111111111100011010;
    rom[706] = 25'b1111111111111111100011010;
    rom[707] = 25'b1111111111111111100011001;
    rom[708] = 25'b1111111111111111100011001;
    rom[709] = 25'b1111111111111111100011001;
    rom[710] = 25'b1111111111111111100011001;
    rom[711] = 25'b1111111111111111100011001;
    rom[712] = 25'b1111111111111111100011000;
    rom[713] = 25'b1111111111111111100011000;
    rom[714] = 25'b1111111111111111100010111;
    rom[715] = 25'b1111111111111111100010111;
    rom[716] = 25'b1111111111111111100010110;
    rom[717] = 25'b1111111111111111100010110;
    rom[718] = 25'b1111111111111111100010110;
    rom[719] = 25'b1111111111111111100010110;
    rom[720] = 25'b1111111111111111100010110;
    rom[721] = 25'b1111111111111111100010101;
    rom[722] = 25'b1111111111111111100010101;
    rom[723] = 25'b1111111111111111100010100;
    rom[724] = 25'b1111111111111111100010100;
    rom[725] = 25'b1111111111111111100010011;
    rom[726] = 25'b1111111111111111100010011;
    rom[727] = 25'b1111111111111111100010011;
    rom[728] = 25'b1111111111111111100010011;
    rom[729] = 25'b1111111111111111100010011;
    rom[730] = 25'b1111111111111111100010010;
    rom[731] = 25'b1111111111111111100010010;
    rom[732] = 25'b1111111111111111100010001;
    rom[733] = 25'b1111111111111111100010001;
    rom[734] = 25'b1111111111111111100010000;
    rom[735] = 25'b1111111111111111100010000;
    rom[736] = 25'b1111111111111111100010000;
    rom[737] = 25'b1111111111111111100010000;
    rom[738] = 25'b1111111111111111100010000;
    rom[739] = 25'b1111111111111111100001111;
    rom[740] = 25'b1111111111111111100001111;
    rom[741] = 25'b1111111111111111100001110;
    rom[742] = 25'b1111111111111111100001110;
    rom[743] = 25'b1111111111111111100001101;
    rom[744] = 25'b1111111111111111100001101;
    rom[745] = 25'b1111111111111111100001101;
    rom[746] = 25'b1111111111111111100001101;
    rom[747] = 25'b1111111111111111100001101;
    rom[748] = 25'b1111111111111111100001100;
    rom[749] = 25'b1111111111111111100001100;
    rom[750] = 25'b1111111111111111100001011;
    rom[751] = 25'b1111111111111111100001011;
    rom[752] = 25'b1111111111111111100001010;
    rom[753] = 25'b1111111111111111100001010;
    rom[754] = 25'b1111111111111111100001010;
    rom[755] = 25'b1111111111111111100001010;
    rom[756] = 25'b1111111111111111100001010;
    rom[757] = 25'b1111111111111111100001001;
    rom[758] = 25'b1111111111111111100001001;
    rom[759] = 25'b1111111111111111100001000;
    rom[760] = 25'b1111111111111111100001000;
    rom[761] = 25'b1111111111111111100000111;
    rom[762] = 25'b1111111111111111100000111;
    rom[763] = 25'b1111111111111111100000111;
    rom[764] = 25'b1111111111111111100000111;
    rom[765] = 25'b1111111111111111100000111;
    rom[766] = 25'b1111111111111111100000110;
    rom[767] = 25'b1111111111111111100000110;
    rom[768] = 25'b1111111111111111100000101;
    rom[769] = 25'b1111111111111111100000101;
    rom[770] = 25'b1111111111111111100000100;
    rom[771] = 25'b1111111111111111100000100;
    rom[772] = 25'b1111111111111111100000100;
    rom[773] = 25'b1111111111111111100000100;
    rom[774] = 25'b1111111111111111100000100;
    rom[775] = 25'b1111111111111111100000011;
    rom[776] = 25'b1111111111111111100000011;
    rom[777] = 25'b1111111111111111100000010;
    rom[778] = 25'b1111111111111111100000010;
    rom[779] = 25'b1111111111111111100000001;
    rom[780] = 25'b1111111111111111100000001;
    rom[781] = 25'b1111111111111111100000001;
    rom[782] = 25'b1111111111111111100000001;
    rom[783] = 25'b1111111111111111100000000;
    rom[784] = 25'b1111111111111111100000000;
    rom[785] = 25'b1111111111111111100000000;
    rom[786] = 25'b1111111111111111011111111;
    rom[787] = 25'b1111111111111111011111111;
    rom[788] = 25'b1111111111111111011111110;
    rom[789] = 25'b1111111111111111011111110;
    rom[790] = 25'b1111111111111111011111110;
    rom[791] = 25'b1111111111111111011111110;
    rom[792] = 25'b1111111111111111011111101;
    rom[793] = 25'b1111111111111111011111101;
    rom[794] = 25'b1111111111111111011111100;
    rom[795] = 25'b1111111111111111011111100;
    rom[796] = 25'b1111111111111111011111100;
    rom[797] = 25'b1111111111111111011111100;
    rom[798] = 25'b1111111111111111011111100;
    rom[799] = 25'b1111111111111111011111011;
    rom[800] = 25'b1111111111111111011111011;
    rom[801] = 25'b1111111111111111011111010;
    rom[802] = 25'b1111111111111111011111010;
    rom[803] = 25'b1111111111111111011111001;
    rom[804] = 25'b1111111111111111011111001;
    rom[805] = 25'b1111111111111111011111001;
    rom[806] = 25'b1111111111111111011111001;
    rom[807] = 25'b1111111111111111011111001;
    rom[808] = 25'b1111111111111111011111000;
    rom[809] = 25'b1111111111111111011111000;
    rom[810] = 25'b1111111111111111011110111;
    rom[811] = 25'b1111111111111111011110111;
    rom[812] = 25'b1111111111111111011110110;
    rom[813] = 25'b1111111111111111011110110;
    rom[814] = 25'b1111111111111111011110110;
    rom[815] = 25'b1111111111111111011110110;
    rom[816] = 25'b1111111111111111011110101;
    rom[817] = 25'b1111111111111111011110101;
    rom[818] = 25'b1111111111111111011110100;
    rom[819] = 25'b1111111111111111011110100;
    rom[820] = 25'b1111111111111111011110100;
    rom[821] = 25'b1111111111111111011110011;
    rom[822] = 25'b1111111111111111011110011;
    rom[823] = 25'b1111111111111111011110011;
    rom[824] = 25'b1111111111111111011110011;
    rom[825] = 25'b1111111111111111011110010;
    rom[826] = 25'b1111111111111111011110010;
    rom[827] = 25'b1111111111111111011110001;
    rom[828] = 25'b1111111111111111011110001;
    rom[829] = 25'b1111111111111111011110000;
    rom[830] = 25'b1111111111111111011110000;
    rom[831] = 25'b1111111111111111011110000;
    rom[832] = 25'b1111111111111111011110000;
    rom[833] = 25'b1111111111111111011110000;
    rom[834] = 25'b1111111111111111011101111;
    rom[835] = 25'b1111111111111111011101111;
    rom[836] = 25'b1111111111111111011101110;
    rom[837] = 25'b1111111111111111011101110;
    rom[838] = 25'b1111111111111111011101101;
    rom[839] = 25'b1111111111111111011101101;
    rom[840] = 25'b1111111111111111011101101;
    rom[841] = 25'b1111111111111111011101101;
    rom[842] = 25'b1111111111111111011101100;
    rom[843] = 25'b1111111111111111011101100;
    rom[844] = 25'b1111111111111111011101011;
    rom[845] = 25'b1111111111111111011101011;
    rom[846] = 25'b1111111111111111011101011;
    rom[847] = 25'b1111111111111111011101010;
    rom[848] = 25'b1111111111111111011101010;
    rom[849] = 25'b1111111111111111011101010;
    rom[850] = 25'b1111111111111111011101010;
    rom[851] = 25'b1111111111111111011101001;
    rom[852] = 25'b1111111111111111011101001;
    rom[853] = 25'b1111111111111111011101000;
    rom[854] = 25'b1111111111111111011101000;
    rom[855] = 25'b1111111111111111011100111;
    rom[856] = 25'b1111111111111111011100111;
    rom[857] = 25'b1111111111111111011100111;
    rom[858] = 25'b1111111111111111011100111;
    rom[859] = 25'b1111111111111111011100111;
    rom[860] = 25'b1111111111111111011100110;
    rom[861] = 25'b1111111111111111011100110;
    rom[862] = 25'b1111111111111111011100101;
    rom[863] = 25'b1111111111111111011100101;
    rom[864] = 25'b1111111111111111011100100;
    rom[865] = 25'b1111111111111111011100100;
    rom[866] = 25'b1111111111111111011100100;
    rom[867] = 25'b1111111111111111011100100;
    rom[868] = 25'b1111111111111111011100011;
    rom[869] = 25'b1111111111111111011100011;
    rom[870] = 25'b1111111111111111011100010;
    rom[871] = 25'b1111111111111111011100010;
    rom[872] = 25'b1111111111111111011100001;
    rom[873] = 25'b1111111111111111011100001;
    rom[874] = 25'b1111111111111111011100001;
    rom[875] = 25'b1111111111111111011100001;
    rom[876] = 25'b1111111111111111011100001;
    rom[877] = 25'b1111111111111111011100000;
    rom[878] = 25'b1111111111111111011100000;
    rom[879] = 25'b1111111111111111011011111;
    rom[880] = 25'b1111111111111111011011111;
    rom[881] = 25'b1111111111111111011011110;
    rom[882] = 25'b1111111111111111011011110;
    rom[883] = 25'b1111111111111111011011110;
    rom[884] = 25'b1111111111111111011011110;
    rom[885] = 25'b1111111111111111011011101;
    rom[886] = 25'b1111111111111111011011101;
    rom[887] = 25'b1111111111111111011011101;
    rom[888] = 25'b1111111111111111011011100;
    rom[889] = 25'b1111111111111111011011100;
    rom[890] = 25'b1111111111111111011011011;
    rom[891] = 25'b1111111111111111011011011;
    rom[892] = 25'b1111111111111111011011011;
    rom[893] = 25'b1111111111111111011011011;
    rom[894] = 25'b1111111111111111011011010;
    rom[895] = 25'b1111111111111111011011010;
    rom[896] = 25'b1111111111111111011011001;
    rom[897] = 25'b1111111111111111011011001;
    rom[898] = 25'b1111111111111111011011000;
    rom[899] = 25'b1111111111111111011011000;
    rom[900] = 25'b1111111111111111011011000;
    rom[901] = 25'b1111111111111111011011000;
    rom[902] = 25'b1111111111111111011011000;
    rom[903] = 25'b1111111111111111011010111;
    rom[904] = 25'b1111111111111111011010111;
    rom[905] = 25'b1111111111111111011010110;
    rom[906] = 25'b1111111111111111011010110;
    rom[907] = 25'b1111111111111111011010101;
    rom[908] = 25'b1111111111111111011010101;
    rom[909] = 25'b1111111111111111011010101;
    rom[910] = 25'b1111111111111111011010101;
    rom[911] = 25'b1111111111111111011010100;
    rom[912] = 25'b1111111111111111011010100;
    rom[913] = 25'b1111111111111111011010011;
    rom[914] = 25'b1111111111111111011010011;
    rom[915] = 25'b1111111111111111011010010;
    rom[916] = 25'b1111111111111111011010010;
    rom[917] = 25'b1111111111111111011010010;
    rom[918] = 25'b1111111111111111011010010;
    rom[919] = 25'b1111111111111111011010010;
    rom[920] = 25'b1111111111111111011010001;
    rom[921] = 25'b1111111111111111011010001;
    rom[922] = 25'b1111111111111111011010000;
    rom[923] = 25'b1111111111111111011010000;
    rom[924] = 25'b1111111111111111011001111;
    rom[925] = 25'b1111111111111111011001111;
    rom[926] = 25'b1111111111111111011001111;
    rom[927] = 25'b1111111111111111011001111;
    rom[928] = 25'b1111111111111111011001110;
    rom[929] = 25'b1111111111111111011001110;
    rom[930] = 25'b1111111111111111011001101;
    rom[931] = 25'b1111111111111111011001101;
    rom[932] = 25'b1111111111111111011001101;
    rom[933] = 25'b1111111111111111011001100;
    rom[934] = 25'b1111111111111111011001100;
    rom[935] = 25'b1111111111111111011001100;
    rom[936] = 25'b1111111111111111011001100;
    rom[937] = 25'b1111111111111111011001011;
    rom[938] = 25'b1111111111111111011001011;
    rom[939] = 25'b1111111111111111011001010;
    rom[940] = 25'b1111111111111111011001010;
    rom[941] = 25'b1111111111111111011001001;
    rom[942] = 25'b1111111111111111011001001;
    rom[943] = 25'b1111111111111111011001001;
    rom[944] = 25'b1111111111111111011001001;
    rom[945] = 25'b1111111111111111011001000;
    rom[946] = 25'b1111111111111111011001000;
    rom[947] = 25'b1111111111111111011001000;
    rom[948] = 25'b1111111111111111011000111;
    rom[949] = 25'b1111111111111111011000111;
    rom[950] = 25'b1111111111111111011000110;
    rom[951] = 25'b1111111111111111011000110;
    rom[952] = 25'b1111111111111111011000110;
    rom[953] = 25'b1111111111111111011000110;
    rom[954] = 25'b1111111111111111011000101;
    rom[955] = 25'b1111111111111111011000101;
    rom[956] = 25'b1111111111111111011000100;
    rom[957] = 25'b1111111111111111011000100;
    rom[958] = 25'b1111111111111111011000011;
    rom[959] = 25'b1111111111111111011000011;
    rom[960] = 25'b1111111111111111011000011;
    rom[961] = 25'b1111111111111111011000011;
    rom[962] = 25'b1111111111111111011000011;
    rom[963] = 25'b1111111111111111011000010;
    rom[964] = 25'b1111111111111111011000010;
    rom[965] = 25'b1111111111111111011000001;
    rom[966] = 25'b1111111111111111011000001;
    rom[967] = 25'b1111111111111111011000000;
    rom[968] = 25'b1111111111111111011000000;
    rom[969] = 25'b1111111111111111011000000;
    rom[970] = 25'b1111111111111111011000000;
    rom[971] = 25'b1111111111111111010111111;
    rom[972] = 25'b1111111111111111010111111;
    rom[973] = 25'b1111111111111111010111111;
    rom[974] = 25'b1111111111111111010111110;
    rom[975] = 25'b1111111111111111010111110;
    rom[976] = 25'b1111111111111111010111110;
    rom[977] = 25'b1111111111111111010111110;
    rom[978] = 25'b1111111111111111010111101;
    rom[979] = 25'b1111111111111111010111101;
    rom[980] = 25'b1111111111111111010111100;
    rom[981] = 25'b1111111111111111010111100;
    rom[982] = 25'b1111111111111111010111011;
    rom[983] = 25'b1111111111111111010111011;
    rom[984] = 25'b1111111111111111010111011;
    rom[985] = 25'b1111111111111111010111011;
    rom[986] = 25'b1111111111111111010111010;
    rom[987] = 25'b1111111111111111010111010;
    rom[988] = 25'b1111111111111111010111010;
    rom[989] = 25'b1111111111111111010111001;
    rom[990] = 25'b1111111111111111010111001;
    rom[991] = 25'b1111111111111111010111000;
    rom[992] = 25'b1111111111111111010111000;
    rom[993] = 25'b1111111111111111010111000;
    rom[994] = 25'b1111111111111111010111000;
    rom[995] = 25'b1111111111111111010110111;
    rom[996] = 25'b1111111111111111010110111;
    rom[997] = 25'b1111111111111111010110110;
    rom[998] = 25'b1111111111111111010110110;
    rom[999] = 25'b1111111111111111010110110;
    rom[1000] = 25'b1111111111111111010110101;
    rom[1001] = 25'b1111111111111111010110101;
    rom[1002] = 25'b1111111111111111010110101;
    rom[1003] = 25'b1111111111111111010110101;
    rom[1004] = 25'b1111111111111111010110100;
    rom[1005] = 25'b1111111111111111010110100;
    rom[1006] = 25'b1111111111111111010110011;
    rom[1007] = 25'b1111111111111111010110011;
    rom[1008] = 25'b1111111111111111010110010;
    rom[1009] = 25'b1111111111111111010110010;
    rom[1010] = 25'b1111111111111111010110010;
    rom[1011] = 25'b1111111111111111010110010;
    rom[1012] = 25'b1111111111111111010110010;
    rom[1013] = 25'b1111111111111111010110001;
    rom[1014] = 25'b1111111111111111010110001;
    rom[1015] = 25'b1111111111111111010110000;
    rom[1016] = 25'b1111111111111111010110000;
    rom[1017] = 25'b1111111111111111010101111;
    rom[1018] = 25'b1111111111111111010101111;
    rom[1019] = 25'b1111111111111111010101111;
    rom[1020] = 25'b1111111111111111010101111;
    rom[1021] = 25'b1111111111111111010101110;
    rom[1022] = 25'b1111111111111111010101110;
    rom[1023] = 25'b1111111111111111010101110;
    rom[1024] = 25'b1111111111111111010101101;
    rom[1025] = 25'b1111111111111111010101101;
    rom[1026] = 25'b1111111111111111010101100;
    rom[1027] = 25'b1111111111111111010101100;
    rom[1028] = 25'b1111111111111111010101100;
    rom[1029] = 25'b1111111111111111010101100;
    rom[1030] = 25'b1111111111111111010101011;
    rom[1031] = 25'b1111111111111111010101011;
    rom[1032] = 25'b1111111111111111010101010;
    rom[1033] = 25'b1111111111111111010101010;
    rom[1034] = 25'b1111111111111111010101010;
    rom[1035] = 25'b1111111111111111010101001;
    rom[1036] = 25'b1111111111111111010101001;
    rom[1037] = 25'b1111111111111111010101001;
    rom[1038] = 25'b1111111111111111010101001;
    rom[1039] = 25'b1111111111111111010101000;
    rom[1040] = 25'b1111111111111111010101000;
    rom[1041] = 25'b1111111111111111010100111;
    rom[1042] = 25'b1111111111111111010100111;
    rom[1043] = 25'b1111111111111111010100110;
    rom[1044] = 25'b1111111111111111010100110;
    rom[1045] = 25'b1111111111111111010100110;
    rom[1046] = 25'b1111111111111111010100110;
    rom[1047] = 25'b1111111111111111010100110;
    rom[1048] = 25'b1111111111111111010100101;
    rom[1049] = 25'b1111111111111111010100101;
    rom[1050] = 25'b1111111111111111010100100;
    rom[1051] = 25'b1111111111111111010100100;
    rom[1052] = 25'b1111111111111111010100011;
    rom[1053] = 25'b1111111111111111010100011;
    rom[1054] = 25'b1111111111111111010100011;
    rom[1055] = 25'b1111111111111111010100011;
    rom[1056] = 25'b1111111111111111010100011;
    rom[1057] = 25'b1111111111111111010100010;
    rom[1058] = 25'b1111111111111111010100010;
    rom[1059] = 25'b1111111111111111010100001;
    rom[1060] = 25'b1111111111111111010100001;
    rom[1061] = 25'b1111111111111111010100000;
    rom[1062] = 25'b1111111111111111010100000;
    rom[1063] = 25'b1111111111111111010100000;
    rom[1064] = 25'b1111111111111111010100000;
    rom[1065] = 25'b1111111111111111010100000;
    rom[1066] = 25'b1111111111111111010011111;
    rom[1067] = 25'b1111111111111111010011111;
    rom[1068] = 25'b1111111111111111010011110;
    rom[1069] = 25'b1111111111111111010011110;
    rom[1070] = 25'b1111111111111111010011101;
    rom[1071] = 25'b1111111111111111010011101;
    rom[1072] = 25'b1111111111111111010011101;
    rom[1073] = 25'b1111111111111111010011101;
    rom[1074] = 25'b1111111111111111010011101;
    rom[1075] = 25'b1111111111111111010011100;
    rom[1076] = 25'b1111111111111111010011100;
    rom[1077] = 25'b1111111111111111010011011;
    rom[1078] = 25'b1111111111111111010011011;
    rom[1079] = 25'b1111111111111111010011010;
    rom[1080] = 25'b1111111111111111010011010;
    rom[1081] = 25'b1111111111111111010011010;
    rom[1082] = 25'b1111111111111111010011010;
    rom[1083] = 25'b1111111111111111010011010;
    rom[1084] = 25'b1111111111111111010011001;
    rom[1085] = 25'b1111111111111111010011001;
    rom[1086] = 25'b1111111111111111010011000;
    rom[1087] = 25'b1111111111111111010011000;
    rom[1088] = 25'b1111111111111111010010111;
    rom[1089] = 25'b1111111111111111010010111;
    rom[1090] = 25'b1111111111111111010010111;
    rom[1091] = 25'b1111111111111111010010111;
    rom[1092] = 25'b1111111111111111010010111;
    rom[1093] = 25'b1111111111111111010010110;
    rom[1094] = 25'b1111111111111111010010110;
    rom[1095] = 25'b1111111111111111010010101;
    rom[1096] = 25'b1111111111111111010010101;
    rom[1097] = 25'b1111111111111111010010100;
    rom[1098] = 25'b1111111111111111010010100;
    rom[1099] = 25'b1111111111111111010010100;
    rom[1100] = 25'b1111111111111111010010100;
    rom[1101] = 25'b1111111111111111010010100;
    rom[1102] = 25'b1111111111111111010010011;
    rom[1103] = 25'b1111111111111111010010011;
    rom[1104] = 25'b1111111111111111010010010;
    rom[1105] = 25'b1111111111111111010010010;
    rom[1106] = 25'b1111111111111111010010001;
    rom[1107] = 25'b1111111111111111010010001;
    rom[1108] = 25'b1111111111111111010010001;
    rom[1109] = 25'b1111111111111111010010001;
    rom[1110] = 25'b1111111111111111010010001;
    rom[1111] = 25'b1111111111111111010010000;
    rom[1112] = 25'b1111111111111111010010000;
    rom[1113] = 25'b1111111111111111010001111;
    rom[1114] = 25'b1111111111111111010001111;
    rom[1115] = 25'b1111111111111111010001111;
    rom[1116] = 25'b1111111111111111010001110;
    rom[1117] = 25'b1111111111111111010001110;
    rom[1118] = 25'b1111111111111111010001110;
    rom[1119] = 25'b1111111111111111010001110;
    rom[1120] = 25'b1111111111111111010001101;
    rom[1121] = 25'b1111111111111111010001101;
    rom[1122] = 25'b1111111111111111010001101;
    rom[1123] = 25'b1111111111111111010001100;
    rom[1124] = 25'b1111111111111111010001100;
    rom[1125] = 25'b1111111111111111010001011;
    rom[1126] = 25'b1111111111111111010001011;
    rom[1127] = 25'b1111111111111111010001011;
    rom[1128] = 25'b1111111111111111010001011;
    rom[1129] = 25'b1111111111111111010001011;
    rom[1130] = 25'b1111111111111111010001010;
    rom[1131] = 25'b1111111111111111010001010;
    rom[1132] = 25'b1111111111111111010001001;
    rom[1133] = 25'b1111111111111111010001001;
    rom[1134] = 25'b1111111111111111010001000;
    rom[1135] = 25'b1111111111111111010001000;
    rom[1136] = 25'b1111111111111111010001000;
    rom[1137] = 25'b1111111111111111010001000;
    rom[1138] = 25'b1111111111111111010001000;
    rom[1139] = 25'b1111111111111111010000111;
    rom[1140] = 25'b1111111111111111010000111;
    rom[1141] = 25'b1111111111111111010000110;
    rom[1142] = 25'b1111111111111111010000110;
    rom[1143] = 25'b1111111111111111010000110;
    rom[1144] = 25'b1111111111111111010000101;
    rom[1145] = 25'b1111111111111111010000101;
    rom[1146] = 25'b1111111111111111010000101;
    rom[1147] = 25'b1111111111111111010000101;
    rom[1148] = 25'b1111111111111111010000100;
    rom[1149] = 25'b1111111111111111010000100;
    rom[1150] = 25'b1111111111111111010000100;
    rom[1151] = 25'b1111111111111111010000011;
    rom[1152] = 25'b1111111111111111010000011;
    rom[1153] = 25'b1111111111111111010000010;
    rom[1154] = 25'b1111111111111111010000010;
    rom[1155] = 25'b1111111111111111010000010;
    rom[1156] = 25'b1111111111111111010000010;
    rom[1157] = 25'b1111111111111111010000010;
    rom[1158] = 25'b1111111111111111010000001;
    rom[1159] = 25'b1111111111111111010000001;
    rom[1160] = 25'b1111111111111111010000000;
    rom[1161] = 25'b1111111111111111010000000;
    rom[1162] = 25'b1111111111111111010000000;
    rom[1163] = 25'b1111111111111111001111111;
    rom[1164] = 25'b1111111111111111001111111;
    rom[1165] = 25'b1111111111111111001111111;
    rom[1166] = 25'b1111111111111111001111111;
    rom[1167] = 25'b1111111111111111001111111;
    rom[1168] = 25'b1111111111111111001111110;
    rom[1169] = 25'b1111111111111111001111110;
    rom[1170] = 25'b1111111111111111001111101;
    rom[1171] = 25'b1111111111111111001111101;
    rom[1172] = 25'b1111111111111111001111101;
    rom[1173] = 25'b1111111111111111001111101;
    rom[1174] = 25'b1111111111111111001111101;
    rom[1175] = 25'b1111111111111111001111100;
    rom[1176] = 25'b1111111111111111001111100;
    rom[1177] = 25'b1111111111111111001111011;
    rom[1178] = 25'b1111111111111111001111011;
    rom[1179] = 25'b1111111111111111001111011;
    rom[1180] = 25'b1111111111111111001111010;
    rom[1181] = 25'b1111111111111111001111010;
    rom[1182] = 25'b1111111111111111001111010;
    rom[1183] = 25'b1111111111111111001111010;
    rom[1184] = 25'b1111111111111111001111010;
    rom[1185] = 25'b1111111111111111001111001;
    rom[1186] = 25'b1111111111111111001111001;
    rom[1187] = 25'b1111111111111111001111000;
    rom[1188] = 25'b1111111111111111001111000;
    rom[1189] = 25'b1111111111111111001111000;
    rom[1190] = 25'b1111111111111111001110111;
    rom[1191] = 25'b1111111111111111001110111;
    rom[1192] = 25'b1111111111111111001110111;
    rom[1193] = 25'b1111111111111111001110111;
    rom[1194] = 25'b1111111111111111001110111;
    rom[1195] = 25'b1111111111111111001110110;
    rom[1196] = 25'b1111111111111111001110110;
    rom[1197] = 25'b1111111111111111001110101;
    rom[1198] = 25'b1111111111111111001110101;
    rom[1199] = 25'b1111111111111111001110101;
    rom[1200] = 25'b1111111111111111001110100;
    rom[1201] = 25'b1111111111111111001110100;
    rom[1202] = 25'b1111111111111111001110100;
    rom[1203] = 25'b1111111111111111001110100;
    rom[1204] = 25'b1111111111111111001110100;
    rom[1205] = 25'b1111111111111111001110011;
    rom[1206] = 25'b1111111111111111001110011;
    rom[1207] = 25'b1111111111111111001110010;
    rom[1208] = 25'b1111111111111111001110010;
    rom[1209] = 25'b1111111111111111001110010;
    rom[1210] = 25'b1111111111111111001110001;
    rom[1211] = 25'b1111111111111111001110001;
    rom[1212] = 25'b1111111111111111001110001;
    rom[1213] = 25'b1111111111111111001110001;
    rom[1214] = 25'b1111111111111111001110001;
    rom[1215] = 25'b1111111111111111001110000;
    rom[1216] = 25'b1111111111111111001110000;
    rom[1217] = 25'b1111111111111111001101111;
    rom[1218] = 25'b1111111111111111001101111;
    rom[1219] = 25'b1111111111111111001101111;
    rom[1220] = 25'b1111111111111111001101110;
    rom[1221] = 25'b1111111111111111001101110;
    rom[1222] = 25'b1111111111111111001101110;
    rom[1223] = 25'b1111111111111111001101110;
    rom[1224] = 25'b1111111111111111001101110;
    rom[1225] = 25'b1111111111111111001101101;
    rom[1226] = 25'b1111111111111111001101101;
    rom[1227] = 25'b1111111111111111001101101;
    rom[1228] = 25'b1111111111111111001101100;
    rom[1229] = 25'b1111111111111111001101100;
    rom[1230] = 25'b1111111111111111001101011;
    rom[1231] = 25'b1111111111111111001101011;
    rom[1232] = 25'b1111111111111111001101011;
    rom[1233] = 25'b1111111111111111001101011;
    rom[1234] = 25'b1111111111111111001101011;
    rom[1235] = 25'b1111111111111111001101011;
    rom[1236] = 25'b1111111111111111001101010;
    rom[1237] = 25'b1111111111111111001101010;
    rom[1238] = 25'b1111111111111111001101001;
    rom[1239] = 25'b1111111111111111001101001;
    rom[1240] = 25'b1111111111111111001101001;
    rom[1241] = 25'b1111111111111111001101000;
    rom[1242] = 25'b1111111111111111001101000;
    rom[1243] = 25'b1111111111111111001101000;
    rom[1244] = 25'b1111111111111111001101000;
    rom[1245] = 25'b1111111111111111001101000;
    rom[1246] = 25'b1111111111111111001100111;
    rom[1247] = 25'b1111111111111111001100111;
    rom[1248] = 25'b1111111111111111001100111;
    rom[1249] = 25'b1111111111111111001100110;
    rom[1250] = 25'b1111111111111111001100110;
    rom[1251] = 25'b1111111111111111001100110;
    rom[1252] = 25'b1111111111111111001100101;
    rom[1253] = 25'b1111111111111111001100101;
    rom[1254] = 25'b1111111111111111001100101;
    rom[1255] = 25'b1111111111111111001100101;
    rom[1256] = 25'b1111111111111111001100101;
    rom[1257] = 25'b1111111111111111001100100;
    rom[1258] = 25'b1111111111111111001100100;
    rom[1259] = 25'b1111111111111111001100100;
    rom[1260] = 25'b1111111111111111001100011;
    rom[1261] = 25'b1111111111111111001100011;
    rom[1262] = 25'b1111111111111111001100010;
    rom[1263] = 25'b1111111111111111001100010;
    rom[1264] = 25'b1111111111111111001100010;
    rom[1265] = 25'b1111111111111111001100010;
    rom[1266] = 25'b1111111111111111001100010;
    rom[1267] = 25'b1111111111111111001100010;
    rom[1268] = 25'b1111111111111111001100001;
    rom[1269] = 25'b1111111111111111001100001;
    rom[1270] = 25'b1111111111111111001100001;
    rom[1271] = 25'b1111111111111111001100000;
    rom[1272] = 25'b1111111111111111001100000;
    rom[1273] = 25'b1111111111111111001100000;
    rom[1274] = 25'b1111111111111111001011111;
    rom[1275] = 25'b1111111111111111001011111;
    rom[1276] = 25'b1111111111111111001011111;
    rom[1277] = 25'b1111111111111111001011111;
    rom[1278] = 25'b1111111111111111001011111;
    rom[1279] = 25'b1111111111111111001011110;
    rom[1280] = 25'b1111111111111111001011110;
    rom[1281] = 25'b1111111111111111001011110;
    rom[1282] = 25'b1111111111111111001011101;
    rom[1283] = 25'b1111111111111111001011101;
    rom[1284] = 25'b1111111111111111001011101;
    rom[1285] = 25'b1111111111111111001011100;
    rom[1286] = 25'b1111111111111111001011100;
    rom[1287] = 25'b1111111111111111001011100;
    rom[1288] = 25'b1111111111111111001011100;
    rom[1289] = 25'b1111111111111111001011100;
    rom[1290] = 25'b1111111111111111001011011;
    rom[1291] = 25'b1111111111111111001011011;
    rom[1292] = 25'b1111111111111111001011011;
    rom[1293] = 25'b1111111111111111001011010;
    rom[1294] = 25'b1111111111111111001011010;
    rom[1295] = 25'b1111111111111111001011010;
    rom[1296] = 25'b1111111111111111001011001;
    rom[1297] = 25'b1111111111111111001011001;
    rom[1298] = 25'b1111111111111111001011001;
    rom[1299] = 25'b1111111111111111001011001;
    rom[1300] = 25'b1111111111111111001011001;
    rom[1301] = 25'b1111111111111111001011001;
    rom[1302] = 25'b1111111111111111001011000;
    rom[1303] = 25'b1111111111111111001011000;
    rom[1304] = 25'b1111111111111111001011000;
    rom[1305] = 25'b1111111111111111001010111;
    rom[1306] = 25'b1111111111111111001010111;
    rom[1307] = 25'b1111111111111111001010111;
    rom[1308] = 25'b1111111111111111001010110;
    rom[1309] = 25'b1111111111111111001010110;
    rom[1310] = 25'b1111111111111111001010110;
    rom[1311] = 25'b1111111111111111001010110;
    rom[1312] = 25'b1111111111111111001010110;
    rom[1313] = 25'b1111111111111111001010110;
    rom[1314] = 25'b1111111111111111001010101;
    rom[1315] = 25'b1111111111111111001010101;
    rom[1316] = 25'b1111111111111111001010101;
    rom[1317] = 25'b1111111111111111001010100;
    rom[1318] = 25'b1111111111111111001010100;
    rom[1319] = 25'b1111111111111111001010100;
    rom[1320] = 25'b1111111111111111001010011;
    rom[1321] = 25'b1111111111111111001010011;
    rom[1322] = 25'b1111111111111111001010011;
    rom[1323] = 25'b1111111111111111001010011;
    rom[1324] = 25'b1111111111111111001010011;
    rom[1325] = 25'b1111111111111111001010011;
    rom[1326] = 25'b1111111111111111001010010;
    rom[1327] = 25'b1111111111111111001010010;
    rom[1328] = 25'b1111111111111111001010010;
    rom[1329] = 25'b1111111111111111001010001;
    rom[1330] = 25'b1111111111111111001010001;
    rom[1331] = 25'b1111111111111111001010001;
    rom[1332] = 25'b1111111111111111001010000;
    rom[1333] = 25'b1111111111111111001010000;
    rom[1334] = 25'b1111111111111111001010000;
    rom[1335] = 25'b1111111111111111001010000;
    rom[1336] = 25'b1111111111111111001010000;
    rom[1337] = 25'b1111111111111111001010000;
    rom[1338] = 25'b1111111111111111001010000;
    rom[1339] = 25'b1111111111111111001001111;
    rom[1340] = 25'b1111111111111111001001111;
    rom[1341] = 25'b1111111111111111001001111;
    rom[1342] = 25'b1111111111111111001001110;
    rom[1343] = 25'b1111111111111111001001110;
    rom[1344] = 25'b1111111111111111001001110;
    rom[1345] = 25'b1111111111111111001001101;
    rom[1346] = 25'b1111111111111111001001101;
    rom[1347] = 25'b1111111111111111001001101;
    rom[1348] = 25'b1111111111111111001001101;
    rom[1349] = 25'b1111111111111111001001101;
    rom[1350] = 25'b1111111111111111001001101;
    rom[1351] = 25'b1111111111111111001001100;
    rom[1352] = 25'b1111111111111111001001100;
    rom[1353] = 25'b1111111111111111001001100;
    rom[1354] = 25'b1111111111111111001001100;
    rom[1355] = 25'b1111111111111111001001011;
    rom[1356] = 25'b1111111111111111001001011;
    rom[1357] = 25'b1111111111111111001001011;
    rom[1358] = 25'b1111111111111111001001010;
    rom[1359] = 25'b1111111111111111001001010;
    rom[1360] = 25'b1111111111111111001001010;
    rom[1361] = 25'b1111111111111111001001010;
    rom[1362] = 25'b1111111111111111001001010;
    rom[1363] = 25'b1111111111111111001001010;
    rom[1364] = 25'b1111111111111111001001010;
    rom[1365] = 25'b1111111111111111001001001;
    rom[1366] = 25'b1111111111111111001001001;
    rom[1367] = 25'b1111111111111111001001001;
    rom[1368] = 25'b1111111111111111001001000;
    rom[1369] = 25'b1111111111111111001001000;
    rom[1370] = 25'b1111111111111111001001000;
    rom[1371] = 25'b1111111111111111001000111;
    rom[1372] = 25'b1111111111111111001000111;
    rom[1373] = 25'b1111111111111111001000111;
    rom[1374] = 25'b1111111111111111001000111;
    rom[1375] = 25'b1111111111111111001000111;
    rom[1376] = 25'b1111111111111111001000111;
    rom[1377] = 25'b1111111111111111001000111;
    rom[1378] = 25'b1111111111111111001000110;
    rom[1379] = 25'b1111111111111111001000110;
    rom[1380] = 25'b1111111111111111001000110;
    rom[1381] = 25'b1111111111111111001000110;
    rom[1382] = 25'b1111111111111111001000101;
    rom[1383] = 25'b1111111111111111001000101;
    rom[1384] = 25'b1111111111111111001000101;
    rom[1385] = 25'b1111111111111111001000100;
    rom[1386] = 25'b1111111111111111001000100;
    rom[1387] = 25'b1111111111111111001000100;
    rom[1388] = 25'b1111111111111111001000100;
    rom[1389] = 25'b1111111111111111001000100;
    rom[1390] = 25'b1111111111111111001000100;
    rom[1391] = 25'b1111111111111111001000100;
    rom[1392] = 25'b1111111111111111001000011;
    rom[1393] = 25'b1111111111111111001000011;
    rom[1394] = 25'b1111111111111111001000011;
    rom[1395] = 25'b1111111111111111001000011;
    rom[1396] = 25'b1111111111111111001000010;
    rom[1397] = 25'b1111111111111111001000010;
    rom[1398] = 25'b1111111111111111001000010;
    rom[1399] = 25'b1111111111111111001000010;
    rom[1400] = 25'b1111111111111111001000001;
    rom[1401] = 25'b1111111111111111001000001;
    rom[1402] = 25'b1111111111111111001000001;
    rom[1403] = 25'b1111111111111111001000001;
    rom[1404] = 25'b1111111111111111001000001;
    rom[1405] = 25'b1111111111111111001000001;
    rom[1406] = 25'b1111111111111111001000001;
    rom[1407] = 25'b1111111111111111001000000;
    rom[1408] = 25'b1111111111111111001000000;
    rom[1409] = 25'b1111111111111111001000000;
    rom[1410] = 25'b1111111111111111001000000;
    rom[1411] = 25'b1111111111111111000111111;
    rom[1412] = 25'b1111111111111111000111111;
    rom[1413] = 25'b1111111111111111000111111;
    rom[1414] = 25'b1111111111111111000111111;
    rom[1415] = 25'b1111111111111111000111110;
    rom[1416] = 25'b1111111111111111000111110;
    rom[1417] = 25'b1111111111111111000111110;
    rom[1418] = 25'b1111111111111111000111110;
    rom[1419] = 25'b1111111111111111000111110;
    rom[1420] = 25'b1111111111111111000111110;
    rom[1421] = 25'b1111111111111111000111110;
    rom[1422] = 25'b1111111111111111000111110;
    rom[1423] = 25'b1111111111111111000111101;
    rom[1424] = 25'b1111111111111111000111101;
    rom[1425] = 25'b1111111111111111000111101;
    rom[1426] = 25'b1111111111111111000111101;
    rom[1427] = 25'b1111111111111111000111100;
    rom[1428] = 25'b1111111111111111000111100;
    rom[1429] = 25'b1111111111111111000111100;
    rom[1430] = 25'b1111111111111111000111100;
    rom[1431] = 25'b1111111111111111000111100;
    rom[1432] = 25'b1111111111111111000111100;
    rom[1433] = 25'b1111111111111111000111100;
    rom[1434] = 25'b1111111111111111000111100;
    rom[1435] = 25'b1111111111111111000111011;
    rom[1436] = 25'b1111111111111111000111011;
    rom[1437] = 25'b1111111111111111000111011;
    rom[1438] = 25'b1111111111111111000111011;
    rom[1439] = 25'b1111111111111111000111010;
    rom[1440] = 25'b1111111111111111000111010;
    rom[1441] = 25'b1111111111111111000111010;
    rom[1442] = 25'b1111111111111111000111010;
    rom[1443] = 25'b1111111111111111000111001;
    rom[1444] = 25'b1111111111111111000111001;
    rom[1445] = 25'b1111111111111111000111001;
    rom[1446] = 25'b1111111111111111000111001;
    rom[1447] = 25'b1111111111111111000111001;
    rom[1448] = 25'b1111111111111111000111001;
    rom[1449] = 25'b1111111111111111000111001;
    rom[1450] = 25'b1111111111111111000111001;
    rom[1451] = 25'b1111111111111111000111001;
    rom[1452] = 25'b1111111111111111000111000;
    rom[1453] = 25'b1111111111111111000111000;
    rom[1454] = 25'b1111111111111111000111000;
    rom[1455] = 25'b1111111111111111000111000;
    rom[1456] = 25'b1111111111111111000111000;
    rom[1457] = 25'b1111111111111111000110111;
    rom[1458] = 25'b1111111111111111000110111;
    rom[1459] = 25'b1111111111111111000110111;
    rom[1460] = 25'b1111111111111111000110111;
    rom[1461] = 25'b1111111111111111000110110;
    rom[1462] = 25'b1111111111111111000110110;
    rom[1463] = 25'b1111111111111111000110110;
    rom[1464] = 25'b1111111111111111000110110;
    rom[1465] = 25'b1111111111111111000110110;
    rom[1466] = 25'b1111111111111111000110110;
    rom[1467] = 25'b1111111111111111000110110;
    rom[1468] = 25'b1111111111111111000110110;
    rom[1469] = 25'b1111111111111111000110110;
    rom[1470] = 25'b1111111111111111000110101;
    rom[1471] = 25'b1111111111111111000110101;
    rom[1472] = 25'b1111111111111111000110101;
    rom[1473] = 25'b1111111111111111000110101;
    rom[1474] = 25'b1111111111111111000110101;
    rom[1475] = 25'b1111111111111111000110100;
    rom[1476] = 25'b1111111111111111000110100;
    rom[1477] = 25'b1111111111111111000110100;
    rom[1478] = 25'b1111111111111111000110100;
    rom[1479] = 25'b1111111111111111000110100;
    rom[1480] = 25'b1111111111111111000110011;
    rom[1481] = 25'b1111111111111111000110011;
    rom[1482] = 25'b1111111111111111000110011;
    rom[1483] = 25'b1111111111111111000110011;
    rom[1484] = 25'b1111111111111111000110011;
    rom[1485] = 25'b1111111111111111000110011;
    rom[1486] = 25'b1111111111111111000110011;
    rom[1487] = 25'b1111111111111111000110011;
    rom[1488] = 25'b1111111111111111000110011;
    rom[1489] = 25'b1111111111111111000110011;
    rom[1490] = 25'b1111111111111111000110010;
    rom[1491] = 25'b1111111111111111000110010;
    rom[1492] = 25'b1111111111111111000110010;
    rom[1493] = 25'b1111111111111111000110010;
    rom[1494] = 25'b1111111111111111000110010;
    rom[1495] = 25'b1111111111111111000110010;
    rom[1496] = 25'b1111111111111111000110001;
    rom[1497] = 25'b1111111111111111000110001;
    rom[1498] = 25'b1111111111111111000110001;
    rom[1499] = 25'b1111111111111111000110001;
    rom[1500] = 25'b1111111111111111000110001;
    rom[1501] = 25'b1111111111111111000110000;
    rom[1502] = 25'b1111111111111111000110000;
    rom[1503] = 25'b1111111111111111000110000;
    rom[1504] = 25'b1111111111111111000110000;
    rom[1505] = 25'b1111111111111111000110000;
    rom[1506] = 25'b1111111111111111000110000;
    rom[1507] = 25'b1111111111111111000110000;
    rom[1508] = 25'b1111111111111111000110000;
    rom[1509] = 25'b1111111111111111000110000;
    rom[1510] = 25'b1111111111111111000110000;
    rom[1511] = 25'b1111111111111111000110000;
    rom[1512] = 25'b1111111111111111000110000;
    rom[1513] = 25'b1111111111111111000101111;
    rom[1514] = 25'b1111111111111111000101111;
    rom[1515] = 25'b1111111111111111000101111;
    rom[1516] = 25'b1111111111111111000101111;
    rom[1517] = 25'b1111111111111111000101111;
    rom[1518] = 25'b1111111111111111000101111;
    rom[1519] = 25'b1111111111111111000101110;
    rom[1520] = 25'b1111111111111111000101110;
    rom[1521] = 25'b1111111111111111000101110;
    rom[1522] = 25'b1111111111111111000101110;
    rom[1523] = 25'b1111111111111111000101110;
    rom[1524] = 25'b1111111111111111000101110;
    rom[1525] = 25'b1111111111111111000101101;
    rom[1526] = 25'b1111111111111111000101101;
    rom[1527] = 25'b1111111111111111000101101;
    rom[1528] = 25'b1111111111111111000101101;
    rom[1529] = 25'b1111111111111111000101101;
    rom[1530] = 25'b1111111111111111000101101;
    rom[1531] = 25'b1111111111111111000101101;
    rom[1532] = 25'b1111111111111111000101101;
    rom[1533] = 25'b1111111111111111000101101;
    rom[1534] = 25'b1111111111111111000101101;
    rom[1535] = 25'b1111111111111111000101101;
    rom[1536] = 25'b1111111111111111000101101;
    rom[1537] = 25'b1111111111111111000101101;
    rom[1538] = 25'b1111111111111111000101100;
    rom[1539] = 25'b1111111111111111000101100;
    rom[1540] = 25'b1111111111111111000101100;
    rom[1541] = 25'b1111111111111111000101100;
    rom[1542] = 25'b1111111111111111000101100;
    rom[1543] = 25'b1111111111111111000101100;
    rom[1544] = 25'b1111111111111111000101100;
    rom[1545] = 25'b1111111111111111000101100;
    rom[1546] = 25'b1111111111111111000101011;
    rom[1547] = 25'b1111111111111111000101011;
    rom[1548] = 25'b1111111111111111000101011;
    rom[1549] = 25'b1111111111111111000101011;
    rom[1550] = 25'b1111111111111111000101011;
    rom[1551] = 25'b1111111111111111000101011;
    rom[1552] = 25'b1111111111111111000101011;
    rom[1553] = 25'b1111111111111111000101010;
    rom[1554] = 25'b1111111111111111000101010;
    rom[1555] = 25'b1111111111111111000101010;
    rom[1556] = 25'b1111111111111111000101010;
    rom[1557] = 25'b1111111111111111000101010;
    rom[1558] = 25'b1111111111111111000101010;
    rom[1559] = 25'b1111111111111111000101010;
    rom[1560] = 25'b1111111111111111000101010;
    rom[1561] = 25'b1111111111111111000101010;
    rom[1562] = 25'b1111111111111111000101010;
    rom[1563] = 25'b1111111111111111000101010;
    rom[1564] = 25'b1111111111111111000101010;
    rom[1565] = 25'b1111111111111111000101010;
    rom[1566] = 25'b1111111111111111000101010;
    rom[1567] = 25'b1111111111111111000101010;
    rom[1568] = 25'b1111111111111111000101010;
    rom[1569] = 25'b1111111111111111000101010;
    rom[1570] = 25'b1111111111111111000101001;
    rom[1571] = 25'b1111111111111111000101001;
    rom[1572] = 25'b1111111111111111000101001;
    rom[1573] = 25'b1111111111111111000101001;
    rom[1574] = 25'b1111111111111111000101001;
    rom[1575] = 25'b1111111111111111000101001;
    rom[1576] = 25'b1111111111111111000101001;
    rom[1577] = 25'b1111111111111111000101001;
    rom[1578] = 25'b1111111111111111000101001;
    rom[1579] = 25'b1111111111111111000101001;
    rom[1580] = 25'b1111111111111111000101000;
    rom[1581] = 25'b1111111111111111000101000;
    rom[1582] = 25'b1111111111111111000101000;
    rom[1583] = 25'b1111111111111111000101000;
    rom[1584] = 25'b1111111111111111000101000;
    rom[1585] = 25'b1111111111111111000101000;
    rom[1586] = 25'b1111111111111111000101000;
    rom[1587] = 25'b1111111111111111000101000;
    rom[1588] = 25'b1111111111111111000101000;
    rom[1589] = 25'b1111111111111111000101000;
    rom[1590] = 25'b1111111111111111000100111;
    rom[1591] = 25'b1111111111111111000100111;
    rom[1592] = 25'b1111111111111111000100111;
    rom[1593] = 25'b1111111111111111000100111;
    rom[1594] = 25'b1111111111111111000100111;
    rom[1595] = 25'b1111111111111111000100111;
    rom[1596] = 25'b1111111111111111000100111;
    rom[1597] = 25'b1111111111111111000100111;
    rom[1598] = 25'b1111111111111111000100111;
    rom[1599] = 25'b1111111111111111000100111;
    rom[1600] = 25'b1111111111111111000100111;
    rom[1601] = 25'b1111111111111111000100111;
    rom[1602] = 25'b1111111111111111000100111;
    rom[1603] = 25'b1111111111111111000100111;
    rom[1604] = 25'b1111111111111111000100111;
    rom[1605] = 25'b1111111111111111000100111;
    rom[1606] = 25'b1111111111111111000100111;
    rom[1607] = 25'b1111111111111111000100111;
    rom[1608] = 25'b1111111111111111000100111;
    rom[1609] = 25'b1111111111111111000100111;
    rom[1610] = 25'b1111111111111111000100111;
    rom[1611] = 25'b1111111111111111000100111;
    rom[1612] = 25'b1111111111111111000100111;
    rom[1613] = 25'b1111111111111111000100111;
    rom[1614] = 25'b1111111111111111000100111;
    rom[1615] = 25'b1111111111111111000100111;
    rom[1616] = 25'b1111111111111111000100111;
    rom[1617] = 25'b1111111111111111000100111;
    rom[1618] = 25'b1111111111111111000100110;
    rom[1619] = 25'b1111111111111111000100110;
    rom[1620] = 25'b1111111111111111000100110;
    rom[1621] = 25'b1111111111111111000100110;
    rom[1622] = 25'b1111111111111111000100110;
    rom[1623] = 25'b1111111111111111000100110;
    rom[1624] = 25'b1111111111111111000100110;
    rom[1625] = 25'b1111111111111111000100110;
    rom[1626] = 25'b1111111111111111000100110;
    rom[1627] = 25'b1111111111111111000100110;
    rom[1628] = 25'b1111111111111111000100110;
    rom[1629] = 25'b1111111111111111000100110;
    rom[1630] = 25'b1111111111111111000100110;
    rom[1631] = 25'b1111111111111111000100110;
    rom[1632] = 25'b1111111111111111000100110;
    rom[1633] = 25'b1111111111111111000100110;
    rom[1634] = 25'b1111111111111111000100110;
    rom[1635] = 25'b1111111111111111000100110;
    rom[1636] = 25'b1111111111111111000100110;
    rom[1637] = 25'b1111111111111111000100110;
    rom[1638] = 25'b1111111111111111000100110;
    rom[1639] = 25'b1111111111111111000100110;
    rom[1640] = 25'b1111111111111111000100110;
    rom[1641] = 25'b1111111111111111000100101;
    rom[1642] = 25'b1111111111111111000100101;
    rom[1643] = 25'b1111111111111111000100101;
    rom[1644] = 25'b1111111111111111000100101;
    rom[1645] = 25'b1111111111111111000100101;
    rom[1646] = 25'b1111111111111111000100101;
    rom[1647] = 25'b1111111111111111000100101;
    rom[1648] = 25'b1111111111111111000100101;
    rom[1649] = 25'b1111111111111111000100101;
    rom[1650] = 25'b1111111111111111000100101;
    rom[1651] = 25'b1111111111111111000100101;
    rom[1652] = 25'b1111111111111111000100101;
    rom[1653] = 25'b1111111111111111000100101;
    rom[1654] = 25'b1111111111111111000100101;
    rom[1655] = 25'b1111111111111111000100101;
    rom[1656] = 25'b1111111111111111000100101;
    rom[1657] = 25'b1111111111111111000100101;
    rom[1658] = 25'b1111111111111111000100101;
    rom[1659] = 25'b1111111111111111000100101;
    rom[1660] = 25'b1111111111111111000100101;
    rom[1661] = 25'b1111111111111111000100101;
    rom[1662] = 25'b1111111111111111000100101;
    rom[1663] = 25'b1111111111111111000100101;
    rom[1664] = 25'b1111111111111111000100101;
    rom[1665] = 25'b1111111111111111000100101;
    rom[1666] = 25'b1111111111111111000100101;
    rom[1667] = 25'b1111111111111111000100101;
    rom[1668] = 25'b1111111111111111000100101;
    rom[1669] = 25'b1111111111111111000100101;
    rom[1670] = 25'b1111111111111111000100101;
    rom[1671] = 25'b1111111111111111000100101;
    rom[1672] = 25'b1111111111111111000100101;
    rom[1673] = 25'b1111111111111111000100101;
    rom[1674] = 25'b1111111111111111000100101;
    rom[1675] = 25'b1111111111111111000100101;
    rom[1676] = 25'b1111111111111111000100101;
    rom[1677] = 25'b1111111111111111000100101;
    rom[1678] = 25'b1111111111111111000100101;
    rom[1679] = 25'b1111111111111111000100101;
    rom[1680] = 25'b1111111111111111000100101;
    rom[1681] = 25'b1111111111111111000100101;
    rom[1682] = 25'b1111111111111111000100101;
    rom[1683] = 25'b1111111111111111000100101;
    rom[1684] = 25'b1111111111111111000100101;
    rom[1685] = 25'b1111111111111111000100101;
    rom[1686] = 25'b1111111111111111000100101;
    rom[1687] = 25'b1111111111111111000100101;
    rom[1688] = 25'b1111111111111111000100101;
    rom[1689] = 25'b1111111111111111000100101;
    rom[1690] = 25'b1111111111111111000100110;
    rom[1691] = 25'b1111111111111111000100110;
    rom[1692] = 25'b1111111111111111000100110;
    rom[1693] = 25'b1111111111111111000100110;
    rom[1694] = 25'b1111111111111111000100110;
    rom[1695] = 25'b1111111111111111000100110;
    rom[1696] = 25'b1111111111111111000100110;
    rom[1697] = 25'b1111111111111111000100110;
    rom[1698] = 25'b1111111111111111000100110;
    rom[1699] = 25'b1111111111111111000100110;
    rom[1700] = 25'b1111111111111111000100110;
    rom[1701] = 25'b1111111111111111000100110;
    rom[1702] = 25'b1111111111111111000100110;
    rom[1703] = 25'b1111111111111111000100110;
    rom[1704] = 25'b1111111111111111000100110;
    rom[1705] = 25'b1111111111111111000100110;
    rom[1706] = 25'b1111111111111111000100110;
    rom[1707] = 25'b1111111111111111000100110;
    rom[1708] = 25'b1111111111111111000100110;
    rom[1709] = 25'b1111111111111111000100110;
    rom[1710] = 25'b1111111111111111000100110;
    rom[1711] = 25'b1111111111111111000100110;
    rom[1712] = 25'b1111111111111111000100110;
    rom[1713] = 25'b1111111111111111000100111;
    rom[1714] = 25'b1111111111111111000100111;
    rom[1715] = 25'b1111111111111111000100111;
    rom[1716] = 25'b1111111111111111000100111;
    rom[1717] = 25'b1111111111111111000100111;
    rom[1718] = 25'b1111111111111111000100111;
    rom[1719] = 25'b1111111111111111000100111;
    rom[1720] = 25'b1111111111111111000100111;
    rom[1721] = 25'b1111111111111111000100111;
    rom[1722] = 25'b1111111111111111000100111;
    rom[1723] = 25'b1111111111111111000100111;
    rom[1724] = 25'b1111111111111111000100111;
    rom[1725] = 25'b1111111111111111000100111;
    rom[1726] = 25'b1111111111111111000100111;
    rom[1727] = 25'b1111111111111111000100111;
    rom[1728] = 25'b1111111111111111000100111;
    rom[1729] = 25'b1111111111111111000100111;
    rom[1730] = 25'b1111111111111111000100111;
    rom[1731] = 25'b1111111111111111000100111;
    rom[1732] = 25'b1111111111111111000100111;
    rom[1733] = 25'b1111111111111111000100111;
    rom[1734] = 25'b1111111111111111000100111;
    rom[1735] = 25'b1111111111111111000100111;
    rom[1736] = 25'b1111111111111111000100111;
    rom[1737] = 25'b1111111111111111000100111;
    rom[1738] = 25'b1111111111111111000100111;
    rom[1739] = 25'b1111111111111111000101000;
    rom[1740] = 25'b1111111111111111000101000;
    rom[1741] = 25'b1111111111111111000101000;
    rom[1742] = 25'b1111111111111111000101000;
    rom[1743] = 25'b1111111111111111000101000;
    rom[1744] = 25'b1111111111111111000101000;
    rom[1745] = 25'b1111111111111111000101000;
    rom[1746] = 25'b1111111111111111000101000;
    rom[1747] = 25'b1111111111111111000101000;
    rom[1748] = 25'b1111111111111111000101000;
    rom[1749] = 25'b1111111111111111000101001;
    rom[1750] = 25'b1111111111111111000101001;
    rom[1751] = 25'b1111111111111111000101001;
    rom[1752] = 25'b1111111111111111000101001;
    rom[1753] = 25'b1111111111111111000101001;
    rom[1754] = 25'b1111111111111111000101001;
    rom[1755] = 25'b1111111111111111000101001;
    rom[1756] = 25'b1111111111111111000101001;
    rom[1757] = 25'b1111111111111111000101001;
    rom[1758] = 25'b1111111111111111000101010;
    rom[1759] = 25'b1111111111111111000101010;
    rom[1760] = 25'b1111111111111111000101010;
    rom[1761] = 25'b1111111111111111000101010;
    rom[1762] = 25'b1111111111111111000101010;
    rom[1763] = 25'b1111111111111111000101010;
    rom[1764] = 25'b1111111111111111000101010;
    rom[1765] = 25'b1111111111111111000101010;
    rom[1766] = 25'b1111111111111111000101010;
    rom[1767] = 25'b1111111111111111000101010;
    rom[1768] = 25'b1111111111111111000101010;
    rom[1769] = 25'b1111111111111111000101010;
    rom[1770] = 25'b1111111111111111000101010;
    rom[1771] = 25'b1111111111111111000101010;
    rom[1772] = 25'b1111111111111111000101010;
    rom[1773] = 25'b1111111111111111000101010;
    rom[1774] = 25'b1111111111111111000101011;
    rom[1775] = 25'b1111111111111111000101011;
    rom[1776] = 25'b1111111111111111000101011;
    rom[1777] = 25'b1111111111111111000101011;
    rom[1778] = 25'b1111111111111111000101011;
    rom[1779] = 25'b1111111111111111000101011;
    rom[1780] = 25'b1111111111111111000101011;
    rom[1781] = 25'b1111111111111111000101100;
    rom[1782] = 25'b1111111111111111000101100;
    rom[1783] = 25'b1111111111111111000101100;
    rom[1784] = 25'b1111111111111111000101100;
    rom[1785] = 25'b1111111111111111000101100;
    rom[1786] = 25'b1111111111111111000101100;
    rom[1787] = 25'b1111111111111111000101101;
    rom[1788] = 25'b1111111111111111000101101;
    rom[1789] = 25'b1111111111111111000101101;
    rom[1790] = 25'b1111111111111111000101101;
    rom[1791] = 25'b1111111111111111000101101;
    rom[1792] = 25'b1111111111111111000101101;
    rom[1793] = 25'b1111111111111111000101101;
    rom[1794] = 25'b1111111111111111000101101;
    rom[1795] = 25'b1111111111111111000101101;
    rom[1796] = 25'b1111111111111111000101101;
    rom[1797] = 25'b1111111111111111000101101;
    rom[1798] = 25'b1111111111111111000101101;
    rom[1799] = 25'b1111111111111111000101110;
    rom[1800] = 25'b1111111111111111000101110;
    rom[1801] = 25'b1111111111111111000101110;
    rom[1802] = 25'b1111111111111111000101110;
    rom[1803] = 25'b1111111111111111000101110;
    rom[1804] = 25'b1111111111111111000101110;
    rom[1805] = 25'b1111111111111111000101111;
    rom[1806] = 25'b1111111111111111000101111;
    rom[1807] = 25'b1111111111111111000101111;
    rom[1808] = 25'b1111111111111111000101111;
    rom[1809] = 25'b1111111111111111000101111;
    rom[1810] = 25'b1111111111111111000101111;
    rom[1811] = 25'b1111111111111111000110000;
    rom[1812] = 25'b1111111111111111000110000;
    rom[1813] = 25'b1111111111111111000110000;
    rom[1814] = 25'b1111111111111111000110000;
    rom[1815] = 25'b1111111111111111000110000;
    rom[1816] = 25'b1111111111111111000110000;
    rom[1817] = 25'b1111111111111111000110000;
    rom[1818] = 25'b1111111111111111000110000;
    rom[1819] = 25'b1111111111111111000110000;
    rom[1820] = 25'b1111111111111111000110000;
    rom[1821] = 25'b1111111111111111000110001;
    rom[1822] = 25'b1111111111111111000110001;
    rom[1823] = 25'b1111111111111111000110001;
    rom[1824] = 25'b1111111111111111000110001;
    rom[1825] = 25'b1111111111111111000110001;
    rom[1826] = 25'b1111111111111111000110010;
    rom[1827] = 25'b1111111111111111000110010;
    rom[1828] = 25'b1111111111111111000110010;
    rom[1829] = 25'b1111111111111111000110010;
    rom[1830] = 25'b1111111111111111000110011;
    rom[1831] = 25'b1111111111111111000110011;
    rom[1832] = 25'b1111111111111111000110011;
    rom[1833] = 25'b1111111111111111000110011;
    rom[1834] = 25'b1111111111111111000110011;
    rom[1835] = 25'b1111111111111111000110011;
    rom[1836] = 25'b1111111111111111000110011;
    rom[1837] = 25'b1111111111111111000110011;
    rom[1838] = 25'b1111111111111111000110011;
    rom[1839] = 25'b1111111111111111000110100;
    rom[1840] = 25'b1111111111111111000110100;
    rom[1841] = 25'b1111111111111111000110100;
    rom[1842] = 25'b1111111111111111000110100;
    rom[1843] = 25'b1111111111111111000110101;
    rom[1844] = 25'b1111111111111111000110101;
    rom[1845] = 25'b1111111111111111000110101;
    rom[1846] = 25'b1111111111111111000110101;
    rom[1847] = 25'b1111111111111111000110101;
    rom[1848] = 25'b1111111111111111000110110;
    rom[1849] = 25'b1111111111111111000110110;
    rom[1850] = 25'b1111111111111111000110110;
    rom[1851] = 25'b1111111111111111000110110;
    rom[1852] = 25'b1111111111111111000110110;
    rom[1853] = 25'b1111111111111111000110110;
    rom[1854] = 25'b1111111111111111000110110;
    rom[1855] = 25'b1111111111111111000110110;
    rom[1856] = 25'b1111111111111111000110111;
    rom[1857] = 25'b1111111111111111000110111;
    rom[1858] = 25'b1111111111111111000110111;
    rom[1859] = 25'b1111111111111111000110111;
    rom[1860] = 25'b1111111111111111000111000;
    rom[1861] = 25'b1111111111111111000111000;
    rom[1862] = 25'b1111111111111111000111000;
    rom[1863] = 25'b1111111111111111000111001;
    rom[1864] = 25'b1111111111111111000111001;
    rom[1865] = 25'b1111111111111111000111001;
    rom[1866] = 25'b1111111111111111000111001;
    rom[1867] = 25'b1111111111111111000111001;
    rom[1868] = 25'b1111111111111111000111001;
    rom[1869] = 25'b1111111111111111000111001;
    rom[1870] = 25'b1111111111111111000111001;
    rom[1871] = 25'b1111111111111111000111010;
    rom[1872] = 25'b1111111111111111000111010;
    rom[1873] = 25'b1111111111111111000111010;
    rom[1874] = 25'b1111111111111111000111011;
    rom[1875] = 25'b1111111111111111000111011;
    rom[1876] = 25'b1111111111111111000111011;
    rom[1877] = 25'b1111111111111111000111011;
    rom[1878] = 25'b1111111111111111000111100;
    rom[1879] = 25'b1111111111111111000111100;
    rom[1880] = 25'b1111111111111111000111100;
    rom[1881] = 25'b1111111111111111000111100;
    rom[1882] = 25'b1111111111111111000111100;
    rom[1883] = 25'b1111111111111111000111100;
    rom[1884] = 25'b1111111111111111000111100;
    rom[1885] = 25'b1111111111111111000111101;
    rom[1886] = 25'b1111111111111111000111101;
    rom[1887] = 25'b1111111111111111000111101;
    rom[1888] = 25'b1111111111111111000111110;
    rom[1889] = 25'b1111111111111111000111110;
    rom[1890] = 25'b1111111111111111000111110;
    rom[1891] = 25'b1111111111111111000111110;
    rom[1892] = 25'b1111111111111111000111110;
    rom[1893] = 25'b1111111111111111000111110;
    rom[1894] = 25'b1111111111111111000111110;
    rom[1895] = 25'b1111111111111111000111111;
    rom[1896] = 25'b1111111111111111000111111;
    rom[1897] = 25'b1111111111111111000111111;
    rom[1898] = 25'b1111111111111111001000000;
    rom[1899] = 25'b1111111111111111001000000;
    rom[1900] = 25'b1111111111111111001000000;
    rom[1901] = 25'b1111111111111111001000001;
    rom[1902] = 25'b1111111111111111001000001;
    rom[1903] = 25'b1111111111111111001000001;
    rom[1904] = 25'b1111111111111111001000001;
    rom[1905] = 25'b1111111111111111001000001;
    rom[1906] = 25'b1111111111111111001000001;
    rom[1907] = 25'b1111111111111111001000010;
    rom[1908] = 25'b1111111111111111001000010;
    rom[1909] = 25'b1111111111111111001000010;
    rom[1910] = 25'b1111111111111111001000011;
    rom[1911] = 25'b1111111111111111001000011;
    rom[1912] = 25'b1111111111111111001000011;
    rom[1913] = 25'b1111111111111111001000100;
    rom[1914] = 25'b1111111111111111001000100;
    rom[1915] = 25'b1111111111111111001000100;
    rom[1916] = 25'b1111111111111111001000100;
    rom[1917] = 25'b1111111111111111001000100;
    rom[1918] = 25'b1111111111111111001000100;
    rom[1919] = 25'b1111111111111111001000101;
    rom[1920] = 25'b1111111111111111001000101;
    rom[1921] = 25'b1111111111111111001000101;
    rom[1922] = 25'b1111111111111111001000110;
    rom[1923] = 25'b1111111111111111001000110;
    rom[1924] = 25'b1111111111111111001000110;
    rom[1925] = 25'b1111111111111111001000111;
    rom[1926] = 25'b1111111111111111001000111;
    rom[1927] = 25'b1111111111111111001000111;
    rom[1928] = 25'b1111111111111111001000111;
    rom[1929] = 25'b1111111111111111001000111;
    rom[1930] = 25'b1111111111111111001001000;
    rom[1931] = 25'b1111111111111111001001000;
    rom[1932] = 25'b1111111111111111001001000;
    rom[1933] = 25'b1111111111111111001001001;
    rom[1934] = 25'b1111111111111111001001001;
    rom[1935] = 25'b1111111111111111001001001;
    rom[1936] = 25'b1111111111111111001001010;
    rom[1937] = 25'b1111111111111111001001010;
    rom[1938] = 25'b1111111111111111001001010;
    rom[1939] = 25'b1111111111111111001001010;
    rom[1940] = 25'b1111111111111111001001010;
    rom[1941] = 25'b1111111111111111001001011;
    rom[1942] = 25'b1111111111111111001001011;
    rom[1943] = 25'b1111111111111111001001011;
    rom[1944] = 25'b1111111111111111001001100;
    rom[1945] = 25'b1111111111111111001001100;
    rom[1946] = 25'b1111111111111111001001101;
    rom[1947] = 25'b1111111111111111001001101;
    rom[1948] = 25'b1111111111111111001001101;
    rom[1949] = 25'b1111111111111111001001101;
    rom[1950] = 25'b1111111111111111001001101;
    rom[1951] = 25'b1111111111111111001001110;
    rom[1952] = 25'b1111111111111111001001110;
    rom[1953] = 25'b1111111111111111001001110;
    rom[1954] = 25'b1111111111111111001001111;
    rom[1955] = 25'b1111111111111111001001111;
    rom[1956] = 25'b1111111111111111001010000;
    rom[1957] = 25'b1111111111111111001010000;
    rom[1958] = 25'b1111111111111111001010000;
    rom[1959] = 25'b1111111111111111001010000;
    rom[1960] = 25'b1111111111111111001010000;
    rom[1961] = 25'b1111111111111111001010001;
    rom[1962] = 25'b1111111111111111001010001;
    rom[1963] = 25'b1111111111111111001010001;
    rom[1964] = 25'b1111111111111111001010010;
    rom[1965] = 25'b1111111111111111001010010;
    rom[1966] = 25'b1111111111111111001010011;
    rom[1967] = 25'b1111111111111111001010011;
    rom[1968] = 25'b1111111111111111001010011;
    rom[1969] = 25'b1111111111111111001010011;
    rom[1970] = 25'b1111111111111111001010011;
    rom[1971] = 25'b1111111111111111001010100;
    rom[1972] = 25'b1111111111111111001010100;
    rom[1973] = 25'b1111111111111111001010101;
    rom[1974] = 25'b1111111111111111001010101;
    rom[1975] = 25'b1111111111111111001010101;
    rom[1976] = 25'b1111111111111111001010110;
    rom[1977] = 25'b1111111111111111001010110;
    rom[1978] = 25'b1111111111111111001010110;
    rom[1979] = 25'b1111111111111111001010110;
    rom[1980] = 25'b1111111111111111001010111;
    rom[1981] = 25'b1111111111111111001010111;
    rom[1982] = 25'b1111111111111111001011000;
    rom[1983] = 25'b1111111111111111001011000;
    rom[1984] = 25'b1111111111111111001011000;
    rom[1985] = 25'b1111111111111111001011001;
    rom[1986] = 25'b1111111111111111001011001;
    rom[1987] = 25'b1111111111111111001011001;
    rom[1988] = 25'b1111111111111111001011001;
    rom[1989] = 25'b1111111111111111001011010;
    rom[1990] = 25'b1111111111111111001011010;
    rom[1991] = 25'b1111111111111111001011011;
    rom[1992] = 25'b1111111111111111001011011;
    rom[1993] = 25'b1111111111111111001011100;
    rom[1994] = 25'b1111111111111111001011100;
    rom[1995] = 25'b1111111111111111001011100;
    rom[1996] = 25'b1111111111111111001011100;
    rom[1997] = 25'b1111111111111111001011100;
    rom[1998] = 25'b1111111111111111001011101;
    rom[1999] = 25'b1111111111111111001011101;
    rom[2000] = 25'b1111111111111111001011110;
    rom[2001] = 25'b1111111111111111001011110;
    rom[2002] = 25'b1111111111111111001011111;
    rom[2003] = 25'b1111111111111111001011111;
    rom[2004] = 25'b1111111111111111001011111;
    rom[2005] = 25'b1111111111111111001011111;
    rom[2006] = 25'b1111111111111111001100000;
    rom[2007] = 25'b1111111111111111001100000;
    rom[2008] = 25'b1111111111111111001100001;
    rom[2009] = 25'b1111111111111111001100001;
    rom[2010] = 25'b1111111111111111001100010;
    rom[2011] = 25'b1111111111111111001100010;
    rom[2012] = 25'b1111111111111111001100010;
    rom[2013] = 25'b1111111111111111001100010;
    rom[2014] = 25'b1111111111111111001100011;
    rom[2015] = 25'b1111111111111111001100011;
    rom[2016] = 25'b1111111111111111001100100;
    rom[2017] = 25'b1111111111111111001100100;
    rom[2018] = 25'b1111111111111111001100101;
    rom[2019] = 25'b1111111111111111001100101;
    rom[2020] = 25'b1111111111111111001100101;
    rom[2021] = 25'b1111111111111111001100101;
    rom[2022] = 25'b1111111111111111001100110;
    rom[2023] = 25'b1111111111111111001100110;
    rom[2024] = 25'b1111111111111111001100111;
    rom[2025] = 25'b1111111111111111001100111;
    rom[2026] = 25'b1111111111111111001101000;
    rom[2027] = 25'b1111111111111111001101000;
    rom[2028] = 25'b1111111111111111001101000;
    rom[2029] = 25'b1111111111111111001101000;
    rom[2030] = 25'b1111111111111111001101001;
    rom[2031] = 25'b1111111111111111001101001;
    rom[2032] = 25'b1111111111111111001101010;
    rom[2033] = 25'b1111111111111111001101010;
    rom[2034] = 25'b1111111111111111001101011;
    rom[2035] = 25'b1111111111111111001101011;
    rom[2036] = 25'b1111111111111111001101011;
    rom[2037] = 25'b1111111111111111001101011;
    rom[2038] = 25'b1111111111111111001101100;
    rom[2039] = 25'b1111111111111111001101100;
    rom[2040] = 25'b1111111111111111001101101;
    rom[2041] = 25'b1111111111111111001101110;
    rom[2042] = 25'b1111111111111111001101110;
    rom[2043] = 25'b1111111111111111001101110;
    rom[2044] = 25'b1111111111111111001101110;
    rom[2045] = 25'b1111111111111111001101111;
    rom[2046] = 25'b1111111111111111001101111;
    rom[2047] = 25'b1111111111111111001110000;
    rom[2048] = 25'b1111111111111111001110000;
    rom[2049] = 25'b1111111111111111001110001;
    rom[2050] = 25'b1111111111111111001110001;
    rom[2051] = 25'b1111111111111111001110001;
    rom[2052] = 25'b1111111111111111001110010;
    rom[2053] = 25'b1111111111111111001110010;
    rom[2054] = 25'b1111111111111111001110011;
    rom[2055] = 25'b1111111111111111001110011;
    rom[2056] = 25'b1111111111111111001110100;
    rom[2057] = 25'b1111111111111111001110100;
    rom[2058] = 25'b1111111111111111001110100;
    rom[2059] = 25'b1111111111111111001110100;
    rom[2060] = 25'b1111111111111111001110101;
    rom[2061] = 25'b1111111111111111001110110;
    rom[2062] = 25'b1111111111111111001110110;
    rom[2063] = 25'b1111111111111111001110111;
    rom[2064] = 25'b1111111111111111001110111;
    rom[2065] = 25'b1111111111111111001110111;
    rom[2066] = 25'b1111111111111111001110111;
    rom[2067] = 25'b1111111111111111001111000;
    rom[2068] = 25'b1111111111111111001111001;
    rom[2069] = 25'b1111111111111111001111001;
    rom[2070] = 25'b1111111111111111001111010;
    rom[2071] = 25'b1111111111111111001111010;
    rom[2072] = 25'b1111111111111111001111010;
    rom[2073] = 25'b1111111111111111001111011;
    rom[2074] = 25'b1111111111111111001111011;
    rom[2075] = 25'b1111111111111111001111100;
    rom[2076] = 25'b1111111111111111001111100;
    rom[2077] = 25'b1111111111111111001111101;
    rom[2078] = 25'b1111111111111111001111101;
    rom[2079] = 25'b1111111111111111001111101;
    rom[2080] = 25'b1111111111111111001111110;
    rom[2081] = 25'b1111111111111111001111110;
    rom[2082] = 25'b1111111111111111001111111;
    rom[2083] = 25'b1111111111111111001111111;
    rom[2084] = 25'b1111111111111111001111111;
    rom[2085] = 25'b1111111111111111010000000;
    rom[2086] = 25'b1111111111111111010000000;
    rom[2087] = 25'b1111111111111111010000001;
    rom[2088] = 25'b1111111111111111010000010;
    rom[2089] = 25'b1111111111111111010000010;
    rom[2090] = 25'b1111111111111111010000010;
    rom[2091] = 25'b1111111111111111010000010;
    rom[2092] = 25'b1111111111111111010000011;
    rom[2093] = 25'b1111111111111111010000100;
    rom[2094] = 25'b1111111111111111010000100;
    rom[2095] = 25'b1111111111111111010000101;
    rom[2096] = 25'b1111111111111111010000101;
    rom[2097] = 25'b1111111111111111010000101;
    rom[2098] = 25'b1111111111111111010000110;
    rom[2099] = 25'b1111111111111111010000110;
    rom[2100] = 25'b1111111111111111010000111;
    rom[2101] = 25'b1111111111111111010001000;
    rom[2102] = 25'b1111111111111111010001000;
    rom[2103] = 25'b1111111111111111010001000;
    rom[2104] = 25'b1111111111111111010001001;
    rom[2105] = 25'b1111111111111111010001001;
    rom[2106] = 25'b1111111111111111010001010;
    rom[2107] = 25'b1111111111111111010001011;
    rom[2108] = 25'b1111111111111111010001011;
    rom[2109] = 25'b1111111111111111010001011;
    rom[2110] = 25'b1111111111111111010001011;
    rom[2111] = 25'b1111111111111111010001100;
    rom[2112] = 25'b1111111111111111010001101;
    rom[2113] = 25'b1111111111111111010001101;
    rom[2114] = 25'b1111111111111111010001110;
    rom[2115] = 25'b1111111111111111010001110;
    rom[2116] = 25'b1111111111111111010001110;
    rom[2117] = 25'b1111111111111111010001111;
    rom[2118] = 25'b1111111111111111010010000;
    rom[2119] = 25'b1111111111111111010010000;
    rom[2120] = 25'b1111111111111111010010001;
    rom[2121] = 25'b1111111111111111010010001;
    rom[2122] = 25'b1111111111111111010010001;
    rom[2123] = 25'b1111111111111111010010010;
    rom[2124] = 25'b1111111111111111010010011;
    rom[2125] = 25'b1111111111111111010010011;
    rom[2126] = 25'b1111111111111111010010100;
    rom[2127] = 25'b1111111111111111010010100;
    rom[2128] = 25'b1111111111111111010010100;
    rom[2129] = 25'b1111111111111111010010101;
    rom[2130] = 25'b1111111111111111010010110;
    rom[2131] = 25'b1111111111111111010010110;
    rom[2132] = 25'b1111111111111111010010111;
    rom[2133] = 25'b1111111111111111010010111;
    rom[2134] = 25'b1111111111111111010011000;
    rom[2135] = 25'b1111111111111111010011000;
    rom[2136] = 25'b1111111111111111010011001;
    rom[2137] = 25'b1111111111111111010011010;
    rom[2138] = 25'b1111111111111111010011010;
    rom[2139] = 25'b1111111111111111010011010;
    rom[2140] = 25'b1111111111111111010011011;
    rom[2141] = 25'b1111111111111111010011011;
    rom[2142] = 25'b1111111111111111010011100;
    rom[2143] = 25'b1111111111111111010011101;
    rom[2144] = 25'b1111111111111111010011101;
    rom[2145] = 25'b1111111111111111010011101;
    rom[2146] = 25'b1111111111111111010011110;
    rom[2147] = 25'b1111111111111111010011111;
    rom[2148] = 25'b1111111111111111010011111;
    rom[2149] = 25'b1111111111111111010100000;
    rom[2150] = 25'b1111111111111111010100000;
    rom[2151] = 25'b1111111111111111010100000;
    rom[2152] = 25'b1111111111111111010100001;
    rom[2153] = 25'b1111111111111111010100010;
    rom[2154] = 25'b1111111111111111010100011;
    rom[2155] = 25'b1111111111111111010100011;
    rom[2156] = 25'b1111111111111111010100011;
    rom[2157] = 25'b1111111111111111010100100;
    rom[2158] = 25'b1111111111111111010100101;
    rom[2159] = 25'b1111111111111111010100101;
    rom[2160] = 25'b1111111111111111010100110;
    rom[2161] = 25'b1111111111111111010100110;
    rom[2162] = 25'b1111111111111111010100110;
    rom[2163] = 25'b1111111111111111010100111;
    rom[2164] = 25'b1111111111111111010101000;
    rom[2165] = 25'b1111111111111111010101001;
    rom[2166] = 25'b1111111111111111010101001;
    rom[2167] = 25'b1111111111111111010101001;
    rom[2168] = 25'b1111111111111111010101010;
    rom[2169] = 25'b1111111111111111010101011;
    rom[2170] = 25'b1111111111111111010101011;
    rom[2171] = 25'b1111111111111111010101100;
    rom[2172] = 25'b1111111111111111010101100;
    rom[2173] = 25'b1111111111111111010101101;
    rom[2174] = 25'b1111111111111111010101101;
    rom[2175] = 25'b1111111111111111010101110;
    rom[2176] = 25'b1111111111111111010101111;
    rom[2177] = 25'b1111111111111111010101111;
    rom[2178] = 25'b1111111111111111010101111;
    rom[2179] = 25'b1111111111111111010110000;
    rom[2180] = 25'b1111111111111111010110001;
    rom[2181] = 25'b1111111111111111010110010;
    rom[2182] = 25'b1111111111111111010110010;
    rom[2183] = 25'b1111111111111111010110010;
    rom[2184] = 25'b1111111111111111010110011;
    rom[2185] = 25'b1111111111111111010110100;
    rom[2186] = 25'b1111111111111111010110101;
    rom[2187] = 25'b1111111111111111010110101;
    rom[2188] = 25'b1111111111111111010110101;
    rom[2189] = 25'b1111111111111111010110110;
    rom[2190] = 25'b1111111111111111010110111;
    rom[2191] = 25'b1111111111111111010110111;
    rom[2192] = 25'b1111111111111111010111000;
    rom[2193] = 25'b1111111111111111010111000;
    rom[2194] = 25'b1111111111111111010111001;
    rom[2195] = 25'b1111111111111111010111010;
    rom[2196] = 25'b1111111111111111010111010;
    rom[2197] = 25'b1111111111111111010111011;
    rom[2198] = 25'b1111111111111111010111011;
    rom[2199] = 25'b1111111111111111010111100;
    rom[2200] = 25'b1111111111111111010111101;
    rom[2201] = 25'b1111111111111111010111101;
    rom[2202] = 25'b1111111111111111010111110;
    rom[2203] = 25'b1111111111111111010111110;
    rom[2204] = 25'b1111111111111111010111111;
    rom[2205] = 25'b1111111111111111011000000;
    rom[2206] = 25'b1111111111111111011000000;
    rom[2207] = 25'b1111111111111111011000000;
    rom[2208] = 25'b1111111111111111011000001;
    rom[2209] = 25'b1111111111111111011000010;
    rom[2210] = 25'b1111111111111111011000011;
    rom[2211] = 25'b1111111111111111011000011;
    rom[2212] = 25'b1111111111111111011000011;
    rom[2213] = 25'b1111111111111111011000100;
    rom[2214] = 25'b1111111111111111011000101;
    rom[2215] = 25'b1111111111111111011000110;
    rom[2216] = 25'b1111111111111111011000110;
    rom[2217] = 25'b1111111111111111011000110;
    rom[2218] = 25'b1111111111111111011000111;
    rom[2219] = 25'b1111111111111111011001000;
    rom[2220] = 25'b1111111111111111011001001;
    rom[2221] = 25'b1111111111111111011001001;
    rom[2222] = 25'b1111111111111111011001010;
    rom[2223] = 25'b1111111111111111011001010;
    rom[2224] = 25'b1111111111111111011001011;
    rom[2225] = 25'b1111111111111111011001100;
    rom[2226] = 25'b1111111111111111011001100;
    rom[2227] = 25'b1111111111111111011001101;
    rom[2228] = 25'b1111111111111111011001110;
    rom[2229] = 25'b1111111111111111011001110;
    rom[2230] = 25'b1111111111111111011001111;
    rom[2231] = 25'b1111111111111111011001111;
    rom[2232] = 25'b1111111111111111011010000;
    rom[2233] = 25'b1111111111111111011010001;
    rom[2234] = 25'b1111111111111111011010010;
    rom[2235] = 25'b1111111111111111011010010;
    rom[2236] = 25'b1111111111111111011010010;
    rom[2237] = 25'b1111111111111111011010011;
    rom[2238] = 25'b1111111111111111011010100;
    rom[2239] = 25'b1111111111111111011010101;
    rom[2240] = 25'b1111111111111111011010101;
    rom[2241] = 25'b1111111111111111011010110;
    rom[2242] = 25'b1111111111111111011010111;
    rom[2243] = 25'b1111111111111111011010111;
    rom[2244] = 25'b1111111111111111011011000;
    rom[2245] = 25'b1111111111111111011011000;
    rom[2246] = 25'b1111111111111111011011001;
    rom[2247] = 25'b1111111111111111011011010;
    rom[2248] = 25'b1111111111111111011011011;
    rom[2249] = 25'b1111111111111111011011011;
    rom[2250] = 25'b1111111111111111011011100;
    rom[2251] = 25'b1111111111111111011011101;
    rom[2252] = 25'b1111111111111111011011101;
    rom[2253] = 25'b1111111111111111011011110;
    rom[2254] = 25'b1111111111111111011011110;
    rom[2255] = 25'b1111111111111111011011111;
    rom[2256] = 25'b1111111111111111011100000;
    rom[2257] = 25'b1111111111111111011100001;
    rom[2258] = 25'b1111111111111111011100001;
    rom[2259] = 25'b1111111111111111011100010;
    rom[2260] = 25'b1111111111111111011100011;
    rom[2261] = 25'b1111111111111111011100011;
    rom[2262] = 25'b1111111111111111011100100;
    rom[2263] = 25'b1111111111111111011100100;
    rom[2264] = 25'b1111111111111111011100101;
    rom[2265] = 25'b1111111111111111011100110;
    rom[2266] = 25'b1111111111111111011100111;
    rom[2267] = 25'b1111111111111111011100111;
    rom[2268] = 25'b1111111111111111011101000;
    rom[2269] = 25'b1111111111111111011101001;
    rom[2270] = 25'b1111111111111111011101010;
    rom[2271] = 25'b1111111111111111011101010;
    rom[2272] = 25'b1111111111111111011101010;
    rom[2273] = 25'b1111111111111111011101011;
    rom[2274] = 25'b1111111111111111011101100;
    rom[2275] = 25'b1111111111111111011101101;
    rom[2276] = 25'b1111111111111111011101101;
    rom[2277] = 25'b1111111111111111011101110;
    rom[2278] = 25'b1111111111111111011101111;
    rom[2279] = 25'b1111111111111111011110000;
    rom[2280] = 25'b1111111111111111011110000;
    rom[2281] = 25'b1111111111111111011110001;
    rom[2282] = 25'b1111111111111111011110010;
    rom[2283] = 25'b1111111111111111011110011;
    rom[2284] = 25'b1111111111111111011110011;
    rom[2285] = 25'b1111111111111111011110100;
    rom[2286] = 25'b1111111111111111011110100;
    rom[2287] = 25'b1111111111111111011110101;
    rom[2288] = 25'b1111111111111111011110110;
    rom[2289] = 25'b1111111111111111011110110;
    rom[2290] = 25'b1111111111111111011110111;
    rom[2291] = 25'b1111111111111111011111000;
    rom[2292] = 25'b1111111111111111011111001;
    rom[2293] = 25'b1111111111111111011111001;
    rom[2294] = 25'b1111111111111111011111010;
    rom[2295] = 25'b1111111111111111011111011;
    rom[2296] = 25'b1111111111111111011111100;
    rom[2297] = 25'b1111111111111111011111100;
    rom[2298] = 25'b1111111111111111011111101;
    rom[2299] = 25'b1111111111111111011111110;
    rom[2300] = 25'b1111111111111111011111110;
    rom[2301] = 25'b1111111111111111011111111;
    rom[2302] = 25'b1111111111111111100000000;
    rom[2303] = 25'b1111111111111111100000001;
    rom[2304] = 25'b1111111111111111100000001;
    rom[2305] = 25'b1111111111111111100000010;
    rom[2306] = 25'b1111111111111111100000011;
    rom[2307] = 25'b1111111111111111100000100;
    rom[2308] = 25'b1111111111111111100000100;
    rom[2309] = 25'b1111111111111111100000101;
    rom[2310] = 25'b1111111111111111100000110;
    rom[2311] = 25'b1111111111111111100000111;
    rom[2312] = 25'b1111111111111111100000111;
    rom[2313] = 25'b1111111111111111100001000;
    rom[2314] = 25'b1111111111111111100001001;
    rom[2315] = 25'b1111111111111111100001010;
    rom[2316] = 25'b1111111111111111100001010;
    rom[2317] = 25'b1111111111111111100001011;
    rom[2318] = 25'b1111111111111111100001011;
    rom[2319] = 25'b1111111111111111100001100;
    rom[2320] = 25'b1111111111111111100001101;
    rom[2321] = 25'b1111111111111111100001101;
    rom[2322] = 25'b1111111111111111100001110;
    rom[2323] = 25'b1111111111111111100001111;
    rom[2324] = 25'b1111111111111111100010000;
    rom[2325] = 25'b1111111111111111100010001;
    rom[2326] = 25'b1111111111111111100010010;
    rom[2327] = 25'b1111111111111111100010011;
    rom[2328] = 25'b1111111111111111100010011;
    rom[2329] = 25'b1111111111111111100010100;
    rom[2330] = 25'b1111111111111111100010101;
    rom[2331] = 25'b1111111111111111100010110;
    rom[2332] = 25'b1111111111111111100010110;
    rom[2333] = 25'b1111111111111111100010111;
    rom[2334] = 25'b1111111111111111100011000;
    rom[2335] = 25'b1111111111111111100011001;
    rom[2336] = 25'b1111111111111111100011001;
    rom[2337] = 25'b1111111111111111100011010;
    rom[2338] = 25'b1111111111111111100011011;
    rom[2339] = 25'b1111111111111111100011100;
    rom[2340] = 25'b1111111111111111100011100;
    rom[2341] = 25'b1111111111111111100011101;
    rom[2342] = 25'b1111111111111111100011110;
    rom[2343] = 25'b1111111111111111100011111;
    rom[2344] = 25'b1111111111111111100011111;
    rom[2345] = 25'b1111111111111111100100000;
    rom[2346] = 25'b1111111111111111100100001;
    rom[2347] = 25'b1111111111111111100100010;
    rom[2348] = 25'b1111111111111111100100010;
    rom[2349] = 25'b1111111111111111100100011;
    rom[2350] = 25'b1111111111111111100100100;
    rom[2351] = 25'b1111111111111111100100101;
    rom[2352] = 25'b1111111111111111100100101;
    rom[2353] = 25'b1111111111111111100100110;
    rom[2354] = 25'b1111111111111111100100111;
    rom[2355] = 25'b1111111111111111100101000;
    rom[2356] = 25'b1111111111111111100101001;
    rom[2357] = 25'b1111111111111111100101010;
    rom[2358] = 25'b1111111111111111100101011;
    rom[2359] = 25'b1111111111111111100101011;
    rom[2360] = 25'b1111111111111111100101100;
    rom[2361] = 25'b1111111111111111100101101;
    rom[2362] = 25'b1111111111111111100101110;
    rom[2363] = 25'b1111111111111111100101110;
    rom[2364] = 25'b1111111111111111100101111;
    rom[2365] = 25'b1111111111111111100110000;
    rom[2366] = 25'b1111111111111111100110001;
    rom[2367] = 25'b1111111111111111100110001;
    rom[2368] = 25'b1111111111111111100110010;
    rom[2369] = 25'b1111111111111111100110011;
    rom[2370] = 25'b1111111111111111100110100;
    rom[2371] = 25'b1111111111111111100110101;
    rom[2372] = 25'b1111111111111111100110110;
    rom[2373] = 25'b1111111111111111100110111;
    rom[2374] = 25'b1111111111111111100110111;
    rom[2375] = 25'b1111111111111111100111000;
    rom[2376] = 25'b1111111111111111100111001;
    rom[2377] = 25'b1111111111111111100111010;
    rom[2378] = 25'b1111111111111111100111010;
    rom[2379] = 25'b1111111111111111100111011;
    rom[2380] = 25'b1111111111111111100111100;
    rom[2381] = 25'b1111111111111111100111101;
    rom[2382] = 25'b1111111111111111100111110;
    rom[2383] = 25'b1111111111111111100111111;
    rom[2384] = 25'b1111111111111111100111111;
    rom[2385] = 25'b1111111111111111101000000;
    rom[2386] = 25'b1111111111111111101000001;
    rom[2387] = 25'b1111111111111111101000010;
    rom[2388] = 25'b1111111111111111101000010;
    rom[2389] = 25'b1111111111111111101000011;
    rom[2390] = 25'b1111111111111111101000101;
    rom[2391] = 25'b1111111111111111101000101;
    rom[2392] = 25'b1111111111111111101000110;
    rom[2393] = 25'b1111111111111111101000111;
    rom[2394] = 25'b1111111111111111101001000;
    rom[2395] = 25'b1111111111111111101001000;
    rom[2396] = 25'b1111111111111111101001001;
    rom[2397] = 25'b1111111111111111101001010;
    rom[2398] = 25'b1111111111111111101001011;
    rom[2399] = 25'b1111111111111111101001100;
    rom[2400] = 25'b1111111111111111101001101;
    rom[2401] = 25'b1111111111111111101001110;
    rom[2402] = 25'b1111111111111111101001110;
    rom[2403] = 25'b1111111111111111101001111;
    rom[2404] = 25'b1111111111111111101010000;
    rom[2405] = 25'b1111111111111111101010001;
    rom[2406] = 25'b1111111111111111101010010;
    rom[2407] = 25'b1111111111111111101010011;
    rom[2408] = 25'b1111111111111111101010100;
    rom[2409] = 25'b1111111111111111101010100;
    rom[2410] = 25'b1111111111111111101010101;
    rom[2411] = 25'b1111111111111111101010110;
    rom[2412] = 25'b1111111111111111101010111;
    rom[2413] = 25'b1111111111111111101011000;
    rom[2414] = 25'b1111111111111111101011001;
    rom[2415] = 25'b1111111111111111101011010;
    rom[2416] = 25'b1111111111111111101011010;
    rom[2417] = 25'b1111111111111111101011011;
    rom[2418] = 25'b1111111111111111101011100;
    rom[2419] = 25'b1111111111111111101011101;
    rom[2420] = 25'b1111111111111111101011110;
    rom[2421] = 25'b1111111111111111101011111;
    rom[2422] = 25'b1111111111111111101100000;
    rom[2423] = 25'b1111111111111111101100000;
    rom[2424] = 25'b1111111111111111101100001;
    rom[2425] = 25'b1111111111111111101100011;
    rom[2426] = 25'b1111111111111111101100011;
    rom[2427] = 25'b1111111111111111101100100;
    rom[2428] = 25'b1111111111111111101100101;
    rom[2429] = 25'b1111111111111111101100110;
    rom[2430] = 25'b1111111111111111101100110;
    rom[2431] = 25'b1111111111111111101101000;
    rom[2432] = 25'b1111111111111111101101001;
    rom[2433] = 25'b1111111111111111101101001;
    rom[2434] = 25'b1111111111111111101101010;
    rom[2435] = 25'b1111111111111111101101011;
    rom[2436] = 25'b1111111111111111101101100;
    rom[2437] = 25'b1111111111111111101101101;
    rom[2438] = 25'b1111111111111111101101110;
    rom[2439] = 25'b1111111111111111101101111;
    rom[2440] = 25'b1111111111111111101101111;
    rom[2441] = 25'b1111111111111111101110001;
    rom[2442] = 25'b1111111111111111101110010;
    rom[2443] = 25'b1111111111111111101110010;
    rom[2444] = 25'b1111111111111111101110011;
    rom[2445] = 25'b1111111111111111101110100;
    rom[2446] = 25'b1111111111111111101110101;
    rom[2447] = 25'b1111111111111111101110110;
    rom[2448] = 25'b1111111111111111101110111;
    rom[2449] = 25'b1111111111111111101111000;
    rom[2450] = 25'b1111111111111111101111000;
    rom[2451] = 25'b1111111111111111101111010;
    rom[2452] = 25'b1111111111111111101111011;
    rom[2453] = 25'b1111111111111111101111011;
    rom[2454] = 25'b1111111111111111101111100;
    rom[2455] = 25'b1111111111111111101111110;
    rom[2456] = 25'b1111111111111111101111110;
    rom[2457] = 25'b1111111111111111101111111;
    rom[2458] = 25'b1111111111111111110000000;
    rom[2459] = 25'b1111111111111111110000000;
    rom[2460] = 25'b1111111111111111110000010;
    rom[2461] = 25'b1111111111111111110000011;
    rom[2462] = 25'b1111111111111111110000011;
    rom[2463] = 25'b1111111111111111110000100;
    rom[2464] = 25'b1111111111111111110000110;
    rom[2465] = 25'b1111111111111111110000110;
    rom[2466] = 25'b1111111111111111110000111;
    rom[2467] = 25'b1111111111111111110001000;
    rom[2468] = 25'b1111111111111111110001001;
    rom[2469] = 25'b1111111111111111110001010;
    rom[2470] = 25'b1111111111111111110001011;
    rom[2471] = 25'b1111111111111111110001100;
    rom[2472] = 25'b1111111111111111110001101;
    rom[2473] = 25'b1111111111111111110001110;
    rom[2474] = 25'b1111111111111111110001111;
    rom[2475] = 25'b1111111111111111110001111;
    rom[2476] = 25'b1111111111111111110010001;
    rom[2477] = 25'b1111111111111111110010010;
    rom[2478] = 25'b1111111111111111110010010;
    rom[2479] = 25'b1111111111111111110010011;
    rom[2480] = 25'b1111111111111111110010101;
    rom[2481] = 25'b1111111111111111110010101;
    rom[2482] = 25'b1111111111111111110010110;
    rom[2483] = 25'b1111111111111111110010111;
    rom[2484] = 25'b1111111111111111110011000;
    rom[2485] = 25'b1111111111111111110011001;
    rom[2486] = 25'b1111111111111111110011010;
    rom[2487] = 25'b1111111111111111110011011;
    rom[2488] = 25'b1111111111111111110011100;
    rom[2489] = 25'b1111111111111111110011101;
    rom[2490] = 25'b1111111111111111110011110;
    rom[2491] = 25'b1111111111111111110011111;
    rom[2492] = 25'b1111111111111111110100000;
    rom[2493] = 25'b1111111111111111110100001;
    rom[2494] = 25'b1111111111111111110100001;
    rom[2495] = 25'b1111111111111111110100011;
    rom[2496] = 25'b1111111111111111110100100;
    rom[2497] = 25'b1111111111111111110100100;
    rom[2498] = 25'b1111111111111111110100110;
    rom[2499] = 25'b1111111111111111110100111;
    rom[2500] = 25'b1111111111111111110100111;
    rom[2501] = 25'b1111111111111111110101000;
    rom[2502] = 25'b1111111111111111110101010;
    rom[2503] = 25'b1111111111111111110101010;
    rom[2504] = 25'b1111111111111111110101011;
    rom[2505] = 25'b1111111111111111110101101;
    rom[2506] = 25'b1111111111111111110101101;
    rom[2507] = 25'b1111111111111111110101110;
    rom[2508] = 25'b1111111111111111110110000;
    rom[2509] = 25'b1111111111111111110110000;
    rom[2510] = 25'b1111111111111111110110001;
    rom[2511] = 25'b1111111111111111110110010;
    rom[2512] = 25'b1111111111111111110110011;
    rom[2513] = 25'b1111111111111111110110100;
    rom[2514] = 25'b1111111111111111110110101;
    rom[2515] = 25'b1111111111111111110110110;
    rom[2516] = 25'b1111111111111111110110111;
    rom[2517] = 25'b1111111111111111110111000;
    rom[2518] = 25'b1111111111111111110111001;
    rom[2519] = 25'b1111111111111111110111010;
    rom[2520] = 25'b1111111111111111110111011;
    rom[2521] = 25'b1111111111111111110111100;
    rom[2522] = 25'b1111111111111111110111101;
    rom[2523] = 25'b1111111111111111110111110;
    rom[2524] = 25'b1111111111111111110111111;
    rom[2525] = 25'b1111111111111111111000000;
    rom[2526] = 25'b1111111111111111111000001;
    rom[2527] = 25'b1111111111111111111000010;
    rom[2528] = 25'b1111111111111111111000011;
    rom[2529] = 25'b1111111111111111111000100;
    rom[2530] = 25'b1111111111111111111000101;
    rom[2531] = 25'b1111111111111111111000110;
    rom[2532] = 25'b1111111111111111111000111;
    rom[2533] = 25'b1111111111111111111001000;
    rom[2534] = 25'b1111111111111111111001001;
    rom[2535] = 25'b1111111111111111111001010;
    rom[2536] = 25'b1111111111111111111001011;
    rom[2537] = 25'b1111111111111111111001100;
    rom[2538] = 25'b1111111111111111111001101;
    rom[2539] = 25'b1111111111111111111001110;
    rom[2540] = 25'b1111111111111111111001111;
    rom[2541] = 25'b1111111111111111111010000;
    rom[2542] = 25'b1111111111111111111010001;
    rom[2543] = 25'b1111111111111111111010010;
    rom[2544] = 25'b1111111111111111111010011;
    rom[2545] = 25'b1111111111111111111010100;
    rom[2546] = 25'b1111111111111111111010101;
    rom[2547] = 25'b1111111111111111111010110;
    rom[2548] = 25'b1111111111111111111010111;
    rom[2549] = 25'b1111111111111111111011000;
    rom[2550] = 25'b1111111111111111111011001;
    rom[2551] = 25'b1111111111111111111011010;
    rom[2552] = 25'b1111111111111111111011100;
    rom[2553] = 25'b1111111111111111111011100;
    rom[2554] = 25'b1111111111111111111011101;
    rom[2555] = 25'b1111111111111111111011111;
    rom[2556] = 25'b1111111111111111111011111;
    rom[2557] = 25'b1111111111111111111100000;
    rom[2558] = 25'b1111111111111111111100010;
    rom[2559] = 25'b1111111111111111111100010;
    rom[2560] = 25'b1111111111111111111100100;
    rom[2561] = 25'b1111111111111111111100101;
    rom[2562] = 25'b1111111111111111111100101;
    rom[2563] = 25'b1111111111111111111100111;
    rom[2564] = 25'b1111111111111111111101000;
    rom[2565] = 25'b1111111111111111111101001;
    rom[2566] = 25'b1111111111111111111101010;
    rom[2567] = 25'b1111111111111111111101011;
    rom[2568] = 25'b1111111111111111111101100;
    rom[2569] = 25'b1111111111111111111101101;
    rom[2570] = 25'b1111111111111111111101110;
    rom[2571] = 25'b1111111111111111111101111;
    rom[2572] = 25'b1111111111111111111110000;
    rom[2573] = 25'b1111111111111111111110001;
    rom[2574] = 25'b1111111111111111111110010;
    rom[2575] = 25'b1111111111111111111110100;
    rom[2576] = 25'b1111111111111111111110100;
    rom[2577] = 25'b1111111111111111111110101;
    rom[2578] = 25'b1111111111111111111110111;
    rom[2579] = 25'b1111111111111111111110111;
    rom[2580] = 25'b1111111111111111111111001;
    rom[2581] = 25'b1111111111111111111111010;
    rom[2582] = 25'b1111111111111111111111010;
    rom[2583] = 25'b1111111111111111111111100;
    rom[2584] = 25'b1111111111111111111111101;
    rom[2585] = 25'b1111111111111111111111110;
    rom[2586] = 25'b1111111111111111111111111;
    rom[2587] = 25'b0000000000000000000000000;
    rom[2588] = 25'b0000000000000000000000000;
    rom[2589] = 25'b0000000000000000000000001;
    rom[2590] = 25'b0000000000000000000000010;
    rom[2591] = 25'b0000000000000000000000011;
    rom[2592] = 25'b0000000000000000000000101;
    rom[2593] = 25'b0000000000000000000000101;
    rom[2594] = 25'b0000000000000000000000111;
    rom[2595] = 25'b0000000000000000000001000;
    rom[2596] = 25'b0000000000000000000001000;
    rom[2597] = 25'b0000000000000000000001010;
    rom[2598] = 25'b0000000000000000000001011;
    rom[2599] = 25'b0000000000000000000001100;
    rom[2600] = 25'b0000000000000000000001101;
    rom[2601] = 25'b0000000000000000000001110;
    rom[2602] = 25'b0000000000000000000001111;
    rom[2603] = 25'b0000000000000000000010001;
    rom[2604] = 25'b0000000000000000000010001;
    rom[2605] = 25'b0000000000000000000010011;
    rom[2606] = 25'b0000000000000000000010100;
    rom[2607] = 25'b0000000000000000000010100;
    rom[2608] = 25'b0000000000000000000010110;
    rom[2609] = 25'b0000000000000000000010111;
    rom[2610] = 25'b0000000000000000000011000;
    rom[2611] = 25'b0000000000000000000011001;
    rom[2612] = 25'b0000000000000000000011010;
    rom[2613] = 25'b0000000000000000000011011;
    rom[2614] = 25'b0000000000000000000011101;
    rom[2615] = 25'b0000000000000000000011101;
    rom[2616] = 25'b0000000000000000000011111;
    rom[2617] = 25'b0000000000000000000100000;
    rom[2618] = 25'b0000000000000000000100001;
    rom[2619] = 25'b0000000000000000000100010;
    rom[2620] = 25'b0000000000000000000100011;
    rom[2621] = 25'b0000000000000000000100100;
    rom[2622] = 25'b0000000000000000000100101;
    rom[2623] = 25'b0000000000000000000100110;
    rom[2624] = 25'b0000000000000000000100111;
    rom[2625] = 25'b0000000000000000000101001;
    rom[2626] = 25'b0000000000000000000101001;
    rom[2627] = 25'b0000000000000000000101011;
    rom[2628] = 25'b0000000000000000000101100;
    rom[2629] = 25'b0000000000000000000101101;
    rom[2630] = 25'b0000000000000000000101110;
    rom[2631] = 25'b0000000000000000000101111;
    rom[2632] = 25'b0000000000000000000110000;
    rom[2633] = 25'b0000000000000000000110010;
    rom[2634] = 25'b0000000000000000000110010;
    rom[2635] = 25'b0000000000000000000110100;
    rom[2636] = 25'b0000000000000000000110101;
    rom[2637] = 25'b0000000000000000000110110;
    rom[2638] = 25'b0000000000000000000110111;
    rom[2639] = 25'b0000000000000000000111000;
    rom[2640] = 25'b0000000000000000000111001;
    rom[2641] = 25'b0000000000000000000111011;
    rom[2642] = 25'b0000000000000000000111011;
    rom[2643] = 25'b0000000000000000000111101;
    rom[2644] = 25'b0000000000000000000111110;
    rom[2645] = 25'b0000000000000000000111111;
    rom[2646] = 25'b0000000000000000001000000;
    rom[2647] = 25'b0000000000000000001000001;
    rom[2648] = 25'b0000000000000000001000010;
    rom[2649] = 25'b0000000000000000001000011;
    rom[2650] = 25'b0000000000000000001000101;
    rom[2651] = 25'b0000000000000000001000110;
    rom[2652] = 25'b0000000000000000001000111;
    rom[2653] = 25'b0000000000000000001001000;
    rom[2654] = 25'b0000000000000000001001001;
    rom[2655] = 25'b0000000000000000001001010;
    rom[2656] = 25'b0000000000000000001001100;
    rom[2657] = 25'b0000000000000000001001100;
    rom[2658] = 25'b0000000000000000001001110;
    rom[2659] = 25'b0000000000000000001001111;
    rom[2660] = 25'b0000000000000000001010000;
    rom[2661] = 25'b0000000000000000001010001;
    rom[2662] = 25'b0000000000000000001010010;
    rom[2663] = 25'b0000000000000000001010011;
    rom[2664] = 25'b0000000000000000001010101;
    rom[2665] = 25'b0000000000000000001010101;
    rom[2666] = 25'b0000000000000000001010111;
    rom[2667] = 25'b0000000000000000001011000;
    rom[2668] = 25'b0000000000000000001011001;
    rom[2669] = 25'b0000000000000000001011011;
    rom[2670] = 25'b0000000000000000001011011;
    rom[2671] = 25'b0000000000000000001011101;
    rom[2672] = 25'b0000000000000000001011110;
    rom[2673] = 25'b0000000000000000001011111;
    rom[2674] = 25'b0000000000000000001100000;
    rom[2675] = 25'b0000000000000000001100001;
    rom[2676] = 25'b0000000000000000001100011;
    rom[2677] = 25'b0000000000000000001100100;
    rom[2678] = 25'b0000000000000000001100101;
    rom[2679] = 25'b0000000000000000001100110;
    rom[2680] = 25'b0000000000000000001100111;
    rom[2681] = 25'b0000000000000000001101000;
    rom[2682] = 25'b0000000000000000001101010;
    rom[2683] = 25'b0000000000000000001101010;
    rom[2684] = 25'b0000000000000000001101100;
    rom[2685] = 25'b0000000000000000001101101;
    rom[2686] = 25'b0000000000000000001101110;
    rom[2687] = 25'b0000000000000000001110000;
    rom[2688] = 25'b0000000000000000001110000;
    rom[2689] = 25'b0000000000000000001110010;
    rom[2690] = 25'b0000000000000000001110011;
    rom[2691] = 25'b0000000000000000001110100;
    rom[2692] = 25'b0000000000000000001110110;
    rom[2693] = 25'b0000000000000000001110110;
    rom[2694] = 25'b0000000000000000001111000;
    rom[2695] = 25'b0000000000000000001111001;
    rom[2696] = 25'b0000000000000000001111010;
    rom[2697] = 25'b0000000000000000001111100;
    rom[2698] = 25'b0000000000000000001111100;
    rom[2699] = 25'b0000000000000000001111110;
    rom[2700] = 25'b0000000000000000001111111;
    rom[2701] = 25'b0000000000000000010000000;
    rom[2702] = 25'b0000000000000000010000001;
    rom[2703] = 25'b0000000000000000010000010;
    rom[2704] = 25'b0000000000000000010000100;
    rom[2705] = 25'b0000000000000000010000100;
    rom[2706] = 25'b0000000000000000010000110;
    rom[2707] = 25'b0000000000000000010000111;
    rom[2708] = 25'b0000000000000000010001000;
    rom[2709] = 25'b0000000000000000010001010;
    rom[2710] = 25'b0000000000000000010001010;
    rom[2711] = 25'b0000000000000000010001100;
    rom[2712] = 25'b0000000000000000010001101;
    rom[2713] = 25'b0000000000000000010001110;
    rom[2714] = 25'b0000000000000000010010000;
    rom[2715] = 25'b0000000000000000010010000;
    rom[2716] = 25'b0000000000000000010010010;
    rom[2717] = 25'b0000000000000000010010011;
    rom[2718] = 25'b0000000000000000010010100;
    rom[2719] = 25'b0000000000000000010010110;
    rom[2720] = 25'b0000000000000000010010110;
    rom[2721] = 25'b0000000000000000010011000;
    rom[2722] = 25'b0000000000000000010011001;
    rom[2723] = 25'b0000000000000000010011010;
    rom[2724] = 25'b0000000000000000010011100;
    rom[2725] = 25'b0000000000000000010011100;
    rom[2726] = 25'b0000000000000000010011110;
    rom[2727] = 25'b0000000000000000010011111;
    rom[2728] = 25'b0000000000000000010100000;
    rom[2729] = 25'b0000000000000000010100010;
    rom[2730] = 25'b0000000000000000010100011;
    rom[2731] = 25'b0000000000000000010100100;
    rom[2732] = 25'b0000000000000000010100101;
    rom[2733] = 25'b0000000000000000010100111;
    rom[2734] = 25'b0000000000000000010101000;
    rom[2735] = 25'b0000000000000000010101001;
    rom[2736] = 25'b0000000000000000010101010;
    rom[2737] = 25'b0000000000000000010101011;
    rom[2738] = 25'b0000000000000000010101101;
    rom[2739] = 25'b0000000000000000010101110;
    rom[2740] = 25'b0000000000000000010101111;
    rom[2741] = 25'b0000000000000000010110001;
    rom[2742] = 25'b0000000000000000010110001;
    rom[2743] = 25'b0000000000000000010110011;
    rom[2744] = 25'b0000000000000000010110100;
    rom[2745] = 25'b0000000000000000010110101;
    rom[2746] = 25'b0000000000000000010110111;
    rom[2747] = 25'b0000000000000000010111000;
    rom[2748] = 25'b0000000000000000010111001;
    rom[2749] = 25'b0000000000000000010111010;
    rom[2750] = 25'b0000000000000000010111100;
    rom[2751] = 25'b0000000000000000010111101;
    rom[2752] = 25'b0000000000000000010111110;
    rom[2753] = 25'b0000000000000000010111111;
    rom[2754] = 25'b0000000000000000011000000;
    rom[2755] = 25'b0000000000000000011000010;
    rom[2756] = 25'b0000000000000000011000010;
    rom[2757] = 25'b0000000000000000011000100;
    rom[2758] = 25'b0000000000000000011000101;
    rom[2759] = 25'b0000000000000000011000110;
    rom[2760] = 25'b0000000000000000011001000;
    rom[2761] = 25'b0000000000000000011001001;
    rom[2762] = 25'b0000000000000000011001010;
    rom[2763] = 25'b0000000000000000011001011;
    rom[2764] = 25'b0000000000000000011001101;
    rom[2765] = 25'b0000000000000000011001110;
    rom[2766] = 25'b0000000000000000011001111;
    rom[2767] = 25'b0000000000000000011010001;
    rom[2768] = 25'b0000000000000000011010010;
    rom[2769] = 25'b0000000000000000011010011;
    rom[2770] = 25'b0000000000000000011010100;
    rom[2771] = 25'b0000000000000000011010110;
    rom[2772] = 25'b0000000000000000011010111;
    rom[2773] = 25'b0000000000000000011011000;
    rom[2774] = 25'b0000000000000000011011010;
    rom[2775] = 25'b0000000000000000011011010;
    rom[2776] = 25'b0000000000000000011011100;
    rom[2777] = 25'b0000000000000000011011101;
    rom[2778] = 25'b0000000000000000011011110;
    rom[2779] = 25'b0000000000000000011100000;
    rom[2780] = 25'b0000000000000000011100001;
    rom[2781] = 25'b0000000000000000011100010;
    rom[2782] = 25'b0000000000000000011100011;
    rom[2783] = 25'b0000000000000000011100101;
    rom[2784] = 25'b0000000000000000011100110;
    rom[2785] = 25'b0000000000000000011100111;
    rom[2786] = 25'b0000000000000000011101001;
    rom[2787] = 25'b0000000000000000011101010;
    rom[2788] = 25'b0000000000000000011101011;
    rom[2789] = 25'b0000000000000000011101100;
    rom[2790] = 25'b0000000000000000011101110;
    rom[2791] = 25'b0000000000000000011101111;
    rom[2792] = 25'b0000000000000000011110000;
    rom[2793] = 25'b0000000000000000011110010;
    rom[2794] = 25'b0000000000000000011110011;
    rom[2795] = 25'b0000000000000000011110100;
    rom[2796] = 25'b0000000000000000011110101;
    rom[2797] = 25'b0000000000000000011110111;
    rom[2798] = 25'b0000000000000000011111000;
    rom[2799] = 25'b0000000000000000011111001;
    rom[2800] = 25'b0000000000000000011111011;
    rom[2801] = 25'b0000000000000000011111100;
    rom[2802] = 25'b0000000000000000011111101;
    rom[2803] = 25'b0000000000000000011111110;
    rom[2804] = 25'b0000000000000000100000000;
    rom[2805] = 25'b0000000000000000100000001;
    rom[2806] = 25'b0000000000000000100000010;
    rom[2807] = 25'b0000000000000000100000011;
    rom[2808] = 25'b0000000000000000100000101;
    rom[2809] = 25'b0000000000000000100000110;
    rom[2810] = 25'b0000000000000000100000111;
    rom[2811] = 25'b0000000000000000100001001;
    rom[2812] = 25'b0000000000000000100001010;
    rom[2813] = 25'b0000000000000000100001011;
    rom[2814] = 25'b0000000000000000100001100;
    rom[2815] = 25'b0000000000000000100001110;
    rom[2816] = 25'b0000000000000000100001111;
    rom[2817] = 25'b0000000000000000100010000;
    rom[2818] = 25'b0000000000000000100010010;
    rom[2819] = 25'b0000000000000000100010011;
    rom[2820] = 25'b0000000000000000100010101;
    rom[2821] = 25'b0000000000000000100010101;
    rom[2822] = 25'b0000000000000000100010111;
    rom[2823] = 25'b0000000000000000100011000;
    rom[2824] = 25'b0000000000000000100011001;
    rom[2825] = 25'b0000000000000000100011011;
    rom[2826] = 25'b0000000000000000100011100;
    rom[2827] = 25'b0000000000000000100011110;
    rom[2828] = 25'b0000000000000000100011110;
    rom[2829] = 25'b0000000000000000100100000;
    rom[2830] = 25'b0000000000000000100100001;
    rom[2831] = 25'b0000000000000000100100011;
    rom[2832] = 25'b0000000000000000100100100;
    rom[2833] = 25'b0000000000000000100100101;
    rom[2834] = 25'b0000000000000000100100111;
    rom[2835] = 25'b0000000000000000100101000;
    rom[2836] = 25'b0000000000000000100101010;
    rom[2837] = 25'b0000000000000000100101010;
    rom[2838] = 25'b0000000000000000100101100;
    rom[2839] = 25'b0000000000000000100101101;
    rom[2840] = 25'b0000000000000000100101111;
    rom[2841] = 25'b0000000000000000100110000;
    rom[2842] = 25'b0000000000000000100110001;
    rom[2843] = 25'b0000000000000000100110011;
    rom[2844] = 25'b0000000000000000100110100;
    rom[2845] = 25'b0000000000000000100110101;
    rom[2846] = 25'b0000000000000000100110110;
    rom[2847] = 25'b0000000000000000100111000;
    rom[2848] = 25'b0000000000000000100111001;
    rom[2849] = 25'b0000000000000000100111011;
    rom[2850] = 25'b0000000000000000100111100;
    rom[2851] = 25'b0000000000000000100111101;
    rom[2852] = 25'b0000000000000000100111111;
    rom[2853] = 25'b0000000000000000101000000;
    rom[2854] = 25'b0000000000000000101000001;
    rom[2855] = 25'b0000000000000000101000010;
    rom[2856] = 25'b0000000000000000101000100;
    rom[2857] = 25'b0000000000000000101000101;
    rom[2858] = 25'b0000000000000000101000111;
    rom[2859] = 25'b0000000000000000101000111;
    rom[2860] = 25'b0000000000000000101001001;
    rom[2861] = 25'b0000000000000000101001010;
    rom[2862] = 25'b0000000000000000101001100;
    rom[2863] = 25'b0000000000000000101001101;
    rom[2864] = 25'b0000000000000000101001110;
    rom[2865] = 25'b0000000000000000101010000;
    rom[2866] = 25'b0000000000000000101010001;
    rom[2867] = 25'b0000000000000000101010011;
    rom[2868] = 25'b0000000000000000101010011;
    rom[2869] = 25'b0000000000000000101010101;
    rom[2870] = 25'b0000000000000000101010110;
    rom[2871] = 25'b0000000000000000101011000;
    rom[2872] = 25'b0000000000000000101011001;
    rom[2873] = 25'b0000000000000000101011010;
    rom[2874] = 25'b0000000000000000101011100;
    rom[2875] = 25'b0000000000000000101011101;
    rom[2876] = 25'b0000000000000000101011111;
    rom[2877] = 25'b0000000000000000101100000;
    rom[2878] = 25'b0000000000000000101100001;
    rom[2879] = 25'b0000000000000000101100010;
    rom[2880] = 25'b0000000000000000101100100;
    rom[2881] = 25'b0000000000000000101100101;
    rom[2882] = 25'b0000000000000000101100111;
    rom[2883] = 25'b0000000000000000101101000;
    rom[2884] = 25'b0000000000000000101101001;
    rom[2885] = 25'b0000000000000000101101011;
    rom[2886] = 25'b0000000000000000101101100;
    rom[2887] = 25'b0000000000000000101101110;
    rom[2888] = 25'b0000000000000000101101111;
    rom[2889] = 25'b0000000000000000101110000;
    rom[2890] = 25'b0000000000000000101110001;
    rom[2891] = 25'b0000000000000000101110011;
    rom[2892] = 25'b0000000000000000101110100;
    rom[2893] = 25'b0000000000000000101110110;
    rom[2894] = 25'b0000000000000000101110111;
    rom[2895] = 25'b0000000000000000101111000;
    rom[2896] = 25'b0000000000000000101111010;
    rom[2897] = 25'b0000000000000000101111011;
    rom[2898] = 25'b0000000000000000101111101;
    rom[2899] = 25'b0000000000000000101111110;
    rom[2900] = 25'b0000000000000000101111111;
    rom[2901] = 25'b0000000000000000110000000;
    rom[2902] = 25'b0000000000000000110000010;
    rom[2903] = 25'b0000000000000000110000011;
    rom[2904] = 25'b0000000000000000110000101;
    rom[2905] = 25'b0000000000000000110000110;
    rom[2906] = 25'b0000000000000000110000111;
    rom[2907] = 25'b0000000000000000110001000;
    rom[2908] = 25'b0000000000000000110001010;
    rom[2909] = 25'b0000000000000000110001011;
    rom[2910] = 25'b0000000000000000110001101;
    rom[2911] = 25'b0000000000000000110001110;
    rom[2912] = 25'b0000000000000000110001111;
    rom[2913] = 25'b0000000000000000110010001;
    rom[2914] = 25'b0000000000000000110010010;
    rom[2915] = 25'b0000000000000000110010100;
    rom[2916] = 25'b0000000000000000110010101;
    rom[2917] = 25'b0000000000000000110010111;
    rom[2918] = 25'b0000000000000000110010111;
    rom[2919] = 25'b0000000000000000110011001;
    rom[2920] = 25'b0000000000000000110011010;
    rom[2921] = 25'b0000000000000000110011100;
    rom[2922] = 25'b0000000000000000110011101;
    rom[2923] = 25'b0000000000000000110011111;
    rom[2924] = 25'b0000000000000000110100000;
    rom[2925] = 25'b0000000000000000110100001;
    rom[2926] = 25'b0000000000000000110100011;
    rom[2927] = 25'b0000000000000000110100100;
    rom[2928] = 25'b0000000000000000110100110;
    rom[2929] = 25'b0000000000000000110100111;
    rom[2930] = 25'b0000000000000000110101001;
    rom[2931] = 25'b0000000000000000110101010;
    rom[2932] = 25'b0000000000000000110101011;
    rom[2933] = 25'b0000000000000000110101100;
    rom[2934] = 25'b0000000000000000110101110;
    rom[2935] = 25'b0000000000000000110101111;
    rom[2936] = 25'b0000000000000000110110001;
    rom[2937] = 25'b0000000000000000110110010;
    rom[2938] = 25'b0000000000000000110110100;
    rom[2939] = 25'b0000000000000000110110101;
    rom[2940] = 25'b0000000000000000110110110;
    rom[2941] = 25'b0000000000000000110111000;
    rom[2942] = 25'b0000000000000000110111001;
    rom[2943] = 25'b0000000000000000110111011;
    rom[2944] = 25'b0000000000000000110111100;
    rom[2945] = 25'b0000000000000000110111110;
    rom[2946] = 25'b0000000000000000110111111;
    rom[2947] = 25'b0000000000000000111000000;
    rom[2948] = 25'b0000000000000000111000001;
    rom[2949] = 25'b0000000000000000111000011;
    rom[2950] = 25'b0000000000000000111000100;
    rom[2951] = 25'b0000000000000000111000110;
    rom[2952] = 25'b0000000000000000111000111;
    rom[2953] = 25'b0000000000000000111001001;
    rom[2954] = 25'b0000000000000000111001010;
    rom[2955] = 25'b0000000000000000111001011;
    rom[2956] = 25'b0000000000000000111001100;
    rom[2957] = 25'b0000000000000000111001110;
    rom[2958] = 25'b0000000000000000111001111;
    rom[2959] = 25'b0000000000000000111010001;
    rom[2960] = 25'b0000000000000000111010010;
    rom[2961] = 25'b0000000000000000111010100;
    rom[2962] = 25'b0000000000000000111010101;
    rom[2963] = 25'b0000000000000000111010110;
    rom[2964] = 25'b0000000000000000111011000;
    rom[2965] = 25'b0000000000000000111011001;
    rom[2966] = 25'b0000000000000000111011011;
    rom[2967] = 25'b0000000000000000111011100;
    rom[2968] = 25'b0000000000000000111011110;
    rom[2969] = 25'b0000000000000000111011111;
    rom[2970] = 25'b0000000000000000111100001;
    rom[2971] = 25'b0000000000000000111100010;
    rom[2972] = 25'b0000000000000000111100011;
    rom[2973] = 25'b0000000000000000111100100;
    rom[2974] = 25'b0000000000000000111100110;
    rom[2975] = 25'b0000000000000000111100111;
    rom[2976] = 25'b0000000000000000111101001;
    rom[2977] = 25'b0000000000000000111101010;
    rom[2978] = 25'b0000000000000000111101100;
    rom[2979] = 25'b0000000000000000111101101;
    rom[2980] = 25'b0000000000000000111101111;
    rom[2981] = 25'b0000000000000000111110000;
    rom[2982] = 25'b0000000000000000111110001;
    rom[2983] = 25'b0000000000000000111110011;
    rom[2984] = 25'b0000000000000000111110100;
    rom[2985] = 25'b0000000000000000111110110;
    rom[2986] = 25'b0000000000000000111110111;
    rom[2987] = 25'b0000000000000000111111001;
    rom[2988] = 25'b0000000000000000111111010;
    rom[2989] = 25'b0000000000000000111111100;
    rom[2990] = 25'b0000000000000000111111101;
    rom[2991] = 25'b0000000000000000111111111;
    rom[2992] = 25'b0000000000000000111111111;
    rom[2993] = 25'b0000000000000001000000001;
    rom[2994] = 25'b0000000000000001000000010;
    rom[2995] = 25'b0000000000000001000000100;
    rom[2996] = 25'b0000000000000001000000101;
    rom[2997] = 25'b0000000000000001000000111;
    rom[2998] = 25'b0000000000000001000001000;
    rom[2999] = 25'b0000000000000001000001010;
    rom[3000] = 25'b0000000000000001000001011;
    rom[3001] = 25'b0000000000000001000001101;
    rom[3002] = 25'b0000000000000001000001110;
    rom[3003] = 25'b0000000000000001000010000;
    rom[3004] = 25'b0000000000000001000010000;
    rom[3005] = 25'b0000000000000001000010010;
    rom[3006] = 25'b0000000000000001000010011;
    rom[3007] = 25'b0000000000000001000010101;
    rom[3008] = 25'b0000000000000001000010110;
    rom[3009] = 25'b0000000000000001000011000;
    rom[3010] = 25'b0000000000000001000011001;
    rom[3011] = 25'b0000000000000001000011011;
    rom[3012] = 25'b0000000000000001000011100;
    rom[3013] = 25'b0000000000000001000011110;
    rom[3014] = 25'b0000000000000001000011111;
    rom[3015] = 25'b0000000000000001000100001;
    rom[3016] = 25'b0000000000000001000100010;
    rom[3017] = 25'b0000000000000001000100011;
    rom[3018] = 25'b0000000000000001000100101;
    rom[3019] = 25'b0000000000000001000100110;
    rom[3020] = 25'b0000000000000001000101000;
    rom[3021] = 25'b0000000000000001000101001;
    rom[3022] = 25'b0000000000000001000101011;
    rom[3023] = 25'b0000000000000001000101100;
    rom[3024] = 25'b0000000000000001000101110;
    rom[3025] = 25'b0000000000000001000101111;
    rom[3026] = 25'b0000000000000001000110001;
    rom[3027] = 25'b0000000000000001000110010;
    rom[3028] = 25'b0000000000000001000110100;
    rom[3029] = 25'b0000000000000001000110101;
    rom[3030] = 25'b0000000000000001000110111;
    rom[3031] = 25'b0000000000000001000111000;
    rom[3032] = 25'b0000000000000001000111001;
    rom[3033] = 25'b0000000000000001000111010;
    rom[3034] = 25'b0000000000000001000111100;
    rom[3035] = 25'b0000000000000001000111101;
    rom[3036] = 25'b0000000000000001000111111;
    rom[3037] = 25'b0000000000000001001000000;
    rom[3038] = 25'b0000000000000001001000010;
    rom[3039] = 25'b0000000000000001001000011;
    rom[3040] = 25'b0000000000000001001000101;
    rom[3041] = 25'b0000000000000001001000110;
    rom[3042] = 25'b0000000000000001001001000;
    rom[3043] = 25'b0000000000000001001001001;
    rom[3044] = 25'b0000000000000001001001011;
    rom[3045] = 25'b0000000000000001001001100;
    rom[3046] = 25'b0000000000000001001001110;
    rom[3047] = 25'b0000000000000001001001111;
    rom[3048] = 25'b0000000000000001001010001;
    rom[3049] = 25'b0000000000000001001010010;
    rom[3050] = 25'b0000000000000001001010011;
    rom[3051] = 25'b0000000000000001001010100;
    rom[3052] = 25'b0000000000000001001010110;
    rom[3053] = 25'b0000000000000001001010111;
    rom[3054] = 25'b0000000000000001001011001;
    rom[3055] = 25'b0000000000000001001011010;
    rom[3056] = 25'b0000000000000001001011100;
    rom[3057] = 25'b0000000000000001001011101;
    rom[3058] = 25'b0000000000000001001011111;
    rom[3059] = 25'b0000000000000001001100000;
    rom[3060] = 25'b0000000000000001001100010;
    rom[3061] = 25'b0000000000000001001100011;
    rom[3062] = 25'b0000000000000001001100101;
    rom[3063] = 25'b0000000000000001001100110;
    rom[3064] = 25'b0000000000000001001101000;
    rom[3065] = 25'b0000000000000001001101001;
    rom[3066] = 25'b0000000000000001001101011;
    rom[3067] = 25'b0000000000000001001101100;
    rom[3068] = 25'b0000000000000001001101110;
    rom[3069] = 25'b0000000000000001001101111;
    rom[3070] = 25'b0000000000000001001110001;
    rom[3071] = 25'b0000000000000001001110010;
    rom[3072] = 25'b0000000000000001001110100;
    rom[3073] = 25'b0000000000000001001110101;
    rom[3074] = 25'b0000000000000001001110110;
    rom[3075] = 25'b0000000000000001001111000;
    rom[3076] = 25'b0000000000000001001111001;
    rom[3077] = 25'b0000000000000001001111011;
    rom[3078] = 25'b0000000000000001001111100;
    rom[3079] = 25'b0000000000000001001111110;
    rom[3080] = 25'b0000000000000001001111111;
    rom[3081] = 25'b0000000000000001010000001;
    rom[3082] = 25'b0000000000000001010000010;
    rom[3083] = 25'b0000000000000001010000011;
    rom[3084] = 25'b0000000000000001010000101;
    rom[3085] = 25'b0000000000000001010000110;
    rom[3086] = 25'b0000000000000001010001000;
    rom[3087] = 25'b0000000000000001010001001;
    rom[3088] = 25'b0000000000000001010001011;
    rom[3089] = 25'b0000000000000001010001100;
    rom[3090] = 25'b0000000000000001010001110;
    rom[3091] = 25'b0000000000000001010001111;
    rom[3092] = 25'b0000000000000001010010001;
    rom[3093] = 25'b0000000000000001010010010;
    rom[3094] = 25'b0000000000000001010010100;
    rom[3095] = 25'b0000000000000001010010101;
    rom[3096] = 25'b0000000000000001010010111;
    rom[3097] = 25'b0000000000000001010011000;
    rom[3098] = 25'b0000000000000001010011010;
    rom[3099] = 25'b0000000000000001010011011;
    rom[3100] = 25'b0000000000000001010011101;
    rom[3101] = 25'b0000000000000001010011110;
    rom[3102] = 25'b0000000000000001010100000;
    rom[3103] = 25'b0000000000000001010100001;
    rom[3104] = 25'b0000000000000001010100011;
    rom[3105] = 25'b0000000000000001010100100;
    rom[3106] = 25'b0000000000000001010100110;
    rom[3107] = 25'b0000000000000001010100111;
    rom[3108] = 25'b0000000000000001010101001;
    rom[3109] = 25'b0000000000000001010101010;
    rom[3110] = 25'b0000000000000001010101100;
    rom[3111] = 25'b0000000000000001010101101;
    rom[3112] = 25'b0000000000000001010101111;
    rom[3113] = 25'b0000000000000001010110000;
    rom[3114] = 25'b0000000000000001010110001;
    rom[3115] = 25'b0000000000000001010110011;
    rom[3116] = 25'b0000000000000001010110100;
    rom[3117] = 25'b0000000000000001010110110;
    rom[3118] = 25'b0000000000000001010110111;
    rom[3119] = 25'b0000000000000001010111001;
    rom[3120] = 25'b0000000000000001010111010;
    rom[3121] = 25'b0000000000000001010111100;
    rom[3122] = 25'b0000000000000001010111101;
    rom[3123] = 25'b0000000000000001010111111;
    rom[3124] = 25'b0000000000000001011000000;
    rom[3125] = 25'b0000000000000001011000010;
    rom[3126] = 25'b0000000000000001011000011;
    rom[3127] = 25'b0000000000000001011000100;
    rom[3128] = 25'b0000000000000001011000110;
    rom[3129] = 25'b0000000000000001011000111;
    rom[3130] = 25'b0000000000000001011001001;
    rom[3131] = 25'b0000000000000001011001010;
    rom[3132] = 25'b0000000000000001011001100;
    rom[3133] = 25'b0000000000000001011001101;
    rom[3134] = 25'b0000000000000001011001111;
    rom[3135] = 25'b0000000000000001011010000;
    rom[3136] = 25'b0000000000000001011010010;
    rom[3137] = 25'b0000000000000001011010011;
    rom[3138] = 25'b0000000000000001011010101;
    rom[3139] = 25'b0000000000000001011010110;
    rom[3140] = 25'b0000000000000001011011000;
    rom[3141] = 25'b0000000000000001011011001;
    rom[3142] = 25'b0000000000000001011011011;
    rom[3143] = 25'b0000000000000001011011100;
    rom[3144] = 25'b0000000000000001011011110;
    rom[3145] = 25'b0000000000000001011011111;
    rom[3146] = 25'b0000000000000001011100001;
    rom[3147] = 25'b0000000000000001011100010;
    rom[3148] = 25'b0000000000000001011100100;
    rom[3149] = 25'b0000000000000001011100101;
    rom[3150] = 25'b0000000000000001011100111;
    rom[3151] = 25'b0000000000000001011101000;
    rom[3152] = 25'b0000000000000001011101010;
    rom[3153] = 25'b0000000000000001011101011;
    rom[3154] = 25'b0000000000000001011101101;
    rom[3155] = 25'b0000000000000001011101110;
    rom[3156] = 25'b0000000000000001011110000;
    rom[3157] = 25'b0000000000000001011110001;
    rom[3158] = 25'b0000000000000001011110011;
    rom[3159] = 25'b0000000000000001011110100;
    rom[3160] = 25'b0000000000000001011110110;
    rom[3161] = 25'b0000000000000001011110111;
    rom[3162] = 25'b0000000000000001011111001;
    rom[3163] = 25'b0000000000000001011111010;
    rom[3164] = 25'b0000000000000001011111100;
    rom[3165] = 25'b0000000000000001011111101;
    rom[3166] = 25'b0000000000000001011111111;
    rom[3167] = 25'b0000000000000001100000000;
    rom[3168] = 25'b0000000000000001100000010;
    rom[3169] = 25'b0000000000000001100000011;
    rom[3170] = 25'b0000000000000001100000101;
    rom[3171] = 25'b0000000000000001100000110;
    rom[3172] = 25'b0000000000000001100001000;
    rom[3173] = 25'b0000000000000001100001001;
    rom[3174] = 25'b0000000000000001100001011;
    rom[3175] = 25'b0000000000000001100001100;
    rom[3176] = 25'b0000000000000001100001110;
    rom[3177] = 25'b0000000000000001100001111;
    rom[3178] = 25'b0000000000000001100010001;
    rom[3179] = 25'b0000000000000001100010010;
    rom[3180] = 25'b0000000000000001100010100;
    rom[3181] = 25'b0000000000000001100010101;
    rom[3182] = 25'b0000000000000001100010111;
    rom[3183] = 25'b0000000000000001100011000;
    rom[3184] = 25'b0000000000000001100011010;
    rom[3185] = 25'b0000000000000001100011011;
    rom[3186] = 25'b0000000000000001100011101;
    rom[3187] = 25'b0000000000000001100011110;
    rom[3188] = 25'b0000000000000001100100000;
    rom[3189] = 25'b0000000000000001100100001;
    rom[3190] = 25'b0000000000000001100100011;
    rom[3191] = 25'b0000000000000001100100100;
    rom[3192] = 25'b0000000000000001100100110;
    rom[3193] = 25'b0000000000000001100100111;
    rom[3194] = 25'b0000000000000001100101001;
    rom[3195] = 25'b0000000000000001100101010;
    rom[3196] = 25'b0000000000000001100101100;
    rom[3197] = 25'b0000000000000001100101101;
    rom[3198] = 25'b0000000000000001100101111;
    rom[3199] = 25'b0000000000000001100110001;
    rom[3200] = 25'b0000000000000001100110010;
    rom[3201] = 25'b0000000000000001100110100;
    rom[3202] = 25'b0000000000000001100110101;
    rom[3203] = 25'b0000000000000001100110111;
    rom[3204] = 25'b0000000000000001100111000;
    rom[3205] = 25'b0000000000000001100111010;
    rom[3206] = 25'b0000000000000001100111011;
    rom[3207] = 25'b0000000000000001100111101;
    rom[3208] = 25'b0000000000000001100111110;
    rom[3209] = 25'b0000000000000001101000000;
    rom[3210] = 25'b0000000000000001101000001;
    rom[3211] = 25'b0000000000000001101000011;
    rom[3212] = 25'b0000000000000001101000100;
    rom[3213] = 25'b0000000000000001101000110;
    rom[3214] = 25'b0000000000000001101000111;
    rom[3215] = 25'b0000000000000001101001001;
    rom[3216] = 25'b0000000000000001101001010;
    rom[3217] = 25'b0000000000000001101001100;
    rom[3218] = 25'b0000000000000001101001101;
    rom[3219] = 25'b0000000000000001101001111;
    rom[3220] = 25'b0000000000000001101010000;
    rom[3221] = 25'b0000000000000001101010010;
    rom[3222] = 25'b0000000000000001101010011;
    rom[3223] = 25'b0000000000000001101010101;
    rom[3224] = 25'b0000000000000001101010110;
    rom[3225] = 25'b0000000000000001101011000;
    rom[3226] = 25'b0000000000000001101011001;
    rom[3227] = 25'b0000000000000001101011011;
    rom[3228] = 25'b0000000000000001101011100;
    rom[3229] = 25'b0000000000000001101011110;
    rom[3230] = 25'b0000000000000001101011111;
    rom[3231] = 25'b0000000000000001101100001;
    rom[3232] = 25'b0000000000000001101100010;
    rom[3233] = 25'b0000000000000001101100100;
    rom[3234] = 25'b0000000000000001101100101;
    rom[3235] = 25'b0000000000000001101100111;
    rom[3236] = 25'b0000000000000001101101000;
    rom[3237] = 25'b0000000000000001101101010;
    rom[3238] = 25'b0000000000000001101101011;
    rom[3239] = 25'b0000000000000001101101101;
    rom[3240] = 25'b0000000000000001101101110;
    rom[3241] = 25'b0000000000000001101110000;
    rom[3242] = 25'b0000000000000001101110001;
    rom[3243] = 25'b0000000000000001101110011;
    rom[3244] = 25'b0000000000000001101110100;
    rom[3245] = 25'b0000000000000001101110110;
    rom[3246] = 25'b0000000000000001101110111;
    rom[3247] = 25'b0000000000000001101111001;
    rom[3248] = 25'b0000000000000001101111010;
    rom[3249] = 25'b0000000000000001101111100;
    rom[3250] = 25'b0000000000000001101111101;
    rom[3251] = 25'b0000000000000001101111111;
    rom[3252] = 25'b0000000000000001110000000;
    rom[3253] = 25'b0000000000000001110000010;
    rom[3254] = 25'b0000000000000001110000011;
    rom[3255] = 25'b0000000000000001110000100;
    rom[3256] = 25'b0000000000000001110000110;
    rom[3257] = 25'b0000000000000001110000111;
    rom[3258] = 25'b0000000000000001110001001;
    rom[3259] = 25'b0000000000000001110001010;
    rom[3260] = 25'b0000000000000001110001100;
    rom[3261] = 25'b0000000000000001110001110;
    rom[3262] = 25'b0000000000000001110010000;
    rom[3263] = 25'b0000000000000001110010001;
    rom[3264] = 25'b0000000000000001110010011;
    rom[3265] = 25'b0000000000000001110010100;
    rom[3266] = 25'b0000000000000001110010110;
    rom[3267] = 25'b0000000000000001110010111;
    rom[3268] = 25'b0000000000000001110011001;
    rom[3269] = 25'b0000000000000001110011010;
    rom[3270] = 25'b0000000000000001110011100;
    rom[3271] = 25'b0000000000000001110011101;
    rom[3272] = 25'b0000000000000001110011111;
    rom[3273] = 25'b0000000000000001110100000;
    rom[3274] = 25'b0000000000000001110100010;
    rom[3275] = 25'b0000000000000001110100011;
    rom[3276] = 25'b0000000000000001110100101;
    rom[3277] = 25'b0000000000000001110100110;
    rom[3278] = 25'b0000000000000001110101000;
    rom[3279] = 25'b0000000000000001110101001;
    rom[3280] = 25'b0000000000000001110101011;
    rom[3281] = 25'b0000000000000001110101100;
    rom[3282] = 25'b0000000000000001110101110;
    rom[3283] = 25'b0000000000000001110101111;
    rom[3284] = 25'b0000000000000001110110001;
    rom[3285] = 25'b0000000000000001110110010;
    rom[3286] = 25'b0000000000000001110110100;
    rom[3287] = 25'b0000000000000001110110101;
    rom[3288] = 25'b0000000000000001110110111;
    rom[3289] = 25'b0000000000000001110111000;
    rom[3290] = 25'b0000000000000001110111010;
    rom[3291] = 25'b0000000000000001110111011;
    rom[3292] = 25'b0000000000000001110111101;
    rom[3293] = 25'b0000000000000001110111110;
    rom[3294] = 25'b0000000000000001111000000;
    rom[3295] = 25'b0000000000000001111000001;
    rom[3296] = 25'b0000000000000001111000011;
    rom[3297] = 25'b0000000000000001111000100;
    rom[3298] = 25'b0000000000000001111000101;
    rom[3299] = 25'b0000000000000001111000111;
    rom[3300] = 25'b0000000000000001111001000;
    rom[3301] = 25'b0000000000000001111001010;
    rom[3302] = 25'b0000000000000001111001011;
    rom[3303] = 25'b0000000000000001111001101;
    rom[3304] = 25'b0000000000000001111001110;
    rom[3305] = 25'b0000000000000001111010000;
    rom[3306] = 25'b0000000000000001111010001;
    rom[3307] = 25'b0000000000000001111010011;
    rom[3308] = 25'b0000000000000001111010100;
    rom[3309] = 25'b0000000000000001111010110;
    rom[3310] = 25'b0000000000000001111010111;
    rom[3311] = 25'b0000000000000001111011001;
    rom[3312] = 25'b0000000000000001111011010;
    rom[3313] = 25'b0000000000000001111011100;
    rom[3314] = 25'b0000000000000001111011101;
    rom[3315] = 25'b0000000000000001111011111;
    rom[3316] = 25'b0000000000000001111100000;
    rom[3317] = 25'b0000000000000001111100010;
    rom[3318] = 25'b0000000000000001111100011;
    rom[3319] = 25'b0000000000000001111100101;
    rom[3320] = 25'b0000000000000001111100110;
    rom[3321] = 25'b0000000000000001111101000;
    rom[3322] = 25'b0000000000000001111101001;
    rom[3323] = 25'b0000000000000001111101011;
    rom[3324] = 25'b0000000000000001111101100;
    rom[3325] = 25'b0000000000000001111101110;
    rom[3326] = 25'b0000000000000001111101111;
    rom[3327] = 25'b0000000000000001111110001;
    rom[3328] = 25'b0000000000000001111110011;
    rom[3329] = 25'b0000000000000001111110101;
    rom[3330] = 25'b0000000000000001111110110;
    rom[3331] = 25'b0000000000000001111111000;
    rom[3332] = 25'b0000000000000001111111001;
    rom[3333] = 25'b0000000000000001111111011;
    rom[3334] = 25'b0000000000000001111111100;
    rom[3335] = 25'b0000000000000001111111110;
    rom[3336] = 25'b0000000000000001111111111;
    rom[3337] = 25'b0000000000000010000000001;
    rom[3338] = 25'b0000000000000010000000010;
    rom[3339] = 25'b0000000000000010000000100;
    rom[3340] = 25'b0000000000000010000000101;
    rom[3341] = 25'b0000000000000010000000110;
    rom[3342] = 25'b0000000000000010000001000;
    rom[3343] = 25'b0000000000000010000001001;
    rom[3344] = 25'b0000000000000010000001011;
    rom[3345] = 25'b0000000000000010000001100;
    rom[3346] = 25'b0000000000000010000001110;
    rom[3347] = 25'b0000000000000010000001111;
    rom[3348] = 25'b0000000000000010000010001;
    rom[3349] = 25'b0000000000000010000010010;
    rom[3350] = 25'b0000000000000010000010100;
    rom[3351] = 25'b0000000000000010000010101;
    rom[3352] = 25'b0000000000000010000010111;
    rom[3353] = 25'b0000000000000010000011000;
    rom[3354] = 25'b0000000000000010000011010;
    rom[3355] = 25'b0000000000000010000011011;
    rom[3356] = 25'b0000000000000010000011101;
    rom[3357] = 25'b0000000000000010000011110;
    rom[3358] = 25'b0000000000000010000100000;
    rom[3359] = 25'b0000000000000010000100001;
    rom[3360] = 25'b0000000000000010000100011;
    rom[3361] = 25'b0000000000000010000100100;
    rom[3362] = 25'b0000000000000010000100110;
    rom[3363] = 25'b0000000000000010000100111;
    rom[3364] = 25'b0000000000000010000101001;
    rom[3365] = 25'b0000000000000010000101010;
    rom[3366] = 25'b0000000000000010000101100;
    rom[3367] = 25'b0000000000000010000101101;
    rom[3368] = 25'b0000000000000010000101111;
    rom[3369] = 25'b0000000000000010000110000;
    rom[3370] = 25'b0000000000000010000110010;
    rom[3371] = 25'b0000000000000010000110011;
    rom[3372] = 25'b0000000000000010000110101;
    rom[3373] = 25'b0000000000000010000110110;
    rom[3374] = 25'b0000000000000010000111000;
    rom[3375] = 25'b0000000000000010000111001;
    rom[3376] = 25'b0000000000000010000111011;
    rom[3377] = 25'b0000000000000010000111100;
    rom[3378] = 25'b0000000000000010000111110;
    rom[3379] = 25'b0000000000000010000111111;
    rom[3380] = 25'b0000000000000010001000001;
    rom[3381] = 25'b0000000000000010001000010;
    rom[3382] = 25'b0000000000000010001000100;
    rom[3383] = 25'b0000000000000010001000101;
    rom[3384] = 25'b0000000000000010001000111;
    rom[3385] = 25'b0000000000000010001001000;
    rom[3386] = 25'b0000000000000010001001010;
    rom[3387] = 25'b0000000000000010001001011;
    rom[3388] = 25'b0000000000000010001001101;
    rom[3389] = 25'b0000000000000010001001110;
    rom[3390] = 25'b0000000000000010001010000;
    rom[3391] = 25'b0000000000000010001010000;
    rom[3392] = 25'b0000000000000010001010010;
    rom[3393] = 25'b0000000000000010001010011;
    rom[3394] = 25'b0000000000000010001010101;
    rom[3395] = 25'b0000000000000010001010110;
    rom[3396] = 25'b0000000000000010001011000;
    rom[3397] = 25'b0000000000000010001011001;
    rom[3398] = 25'b0000000000000010001011011;
    rom[3399] = 25'b0000000000000010001011100;
    rom[3400] = 25'b0000000000000010001011110;
    rom[3401] = 25'b0000000000000010001011111;
    rom[3402] = 25'b0000000000000010001100001;
    rom[3403] = 25'b0000000000000010001100010;
    rom[3404] = 25'b0000000000000010001100100;
    rom[3405] = 25'b0000000000000010001100101;
    rom[3406] = 25'b0000000000000010001100111;
    rom[3407] = 25'b0000000000000010001101000;
    rom[3408] = 25'b0000000000000010001101010;
    rom[3409] = 25'b0000000000000010001101011;
    rom[3410] = 25'b0000000000000010001101101;
    rom[3411] = 25'b0000000000000010001101110;
    rom[3412] = 25'b0000000000000010001110000;
    rom[3413] = 25'b0000000000000010001110001;
    rom[3414] = 25'b0000000000000010001110011;
    rom[3415] = 25'b0000000000000010001110100;
    rom[3416] = 25'b0000000000000010001110110;
    rom[3417] = 25'b0000000000000010001110111;
    rom[3418] = 25'b0000000000000010001111001;
    rom[3419] = 25'b0000000000000010001111010;
    rom[3420] = 25'b0000000000000010001111100;
    rom[3421] = 25'b0000000000000010001111101;
    rom[3422] = 25'b0000000000000010001111111;
    rom[3423] = 25'b0000000000000010010000000;
    rom[3424] = 25'b0000000000000010010000010;
    rom[3425] = 25'b0000000000000010010000011;
    rom[3426] = 25'b0000000000000010010000101;
    rom[3427] = 25'b0000000000000010010000110;
    rom[3428] = 25'b0000000000000010010001000;
    rom[3429] = 25'b0000000000000010010001001;
    rom[3430] = 25'b0000000000000010010001011;
    rom[3431] = 25'b0000000000000010010001100;
    rom[3432] = 25'b0000000000000010010001110;
    rom[3433] = 25'b0000000000000010010001111;
    rom[3434] = 25'b0000000000000010010010000;
    rom[3435] = 25'b0000000000000010010010001;
    rom[3436] = 25'b0000000000000010010010011;
    rom[3437] = 25'b0000000000000010010010100;
    rom[3438] = 25'b0000000000000010010010110;
    rom[3439] = 25'b0000000000000010010010111;
    rom[3440] = 25'b0000000000000010010011001;
    rom[3441] = 25'b0000000000000010010011010;
    rom[3442] = 25'b0000000000000010010011100;
    rom[3443] = 25'b0000000000000010010011101;
    rom[3444] = 25'b0000000000000010010011111;
    rom[3445] = 25'b0000000000000010010100000;
    rom[3446] = 25'b0000000000000010010100010;
    rom[3447] = 25'b0000000000000010010100011;
    rom[3448] = 25'b0000000000000010010100101;
    rom[3449] = 25'b0000000000000010010100110;
    rom[3450] = 25'b0000000000000010010101000;
    rom[3451] = 25'b0000000000000010010101001;
    rom[3452] = 25'b0000000000000010010101011;
    rom[3453] = 25'b0000000000000010010101100;
    rom[3454] = 25'b0000000000000010010101110;
    rom[3455] = 25'b0000000000000010010101111;
    rom[3456] = 25'b0000000000000010010110001;
    rom[3457] = 25'b0000000000000010010110010;
    rom[3458] = 25'b0000000000000010010110011;
    rom[3459] = 25'b0000000000000010010110101;
    rom[3460] = 25'b0000000000000010010110110;
    rom[3461] = 25'b0000000000000010010111000;
    rom[3462] = 25'b0000000000000010010111001;
    rom[3463] = 25'b0000000000000010010111011;
    rom[3464] = 25'b0000000000000010010111100;
    rom[3465] = 25'b0000000000000010010111110;
    rom[3466] = 25'b0000000000000010010111111;
    rom[3467] = 25'b0000000000000010011000001;
    rom[3468] = 25'b0000000000000010011000010;
    rom[3469] = 25'b0000000000000010011000100;
    rom[3470] = 25'b0000000000000010011000101;
    rom[3471] = 25'b0000000000000010011000110;
    rom[3472] = 25'b0000000000000010011001000;
    rom[3473] = 25'b0000000000000010011001001;
    rom[3474] = 25'b0000000000000010011001011;
    rom[3475] = 25'b0000000000000010011001100;
    rom[3476] = 25'b0000000000000010011001101;
    rom[3477] = 25'b0000000000000010011001111;
    rom[3478] = 25'b0000000000000010011010000;
    rom[3479] = 25'b0000000000000010011010010;
    rom[3480] = 25'b0000000000000010011010011;
    rom[3481] = 25'b0000000000000010011010101;
    rom[3482] = 25'b0000000000000010011010110;
    rom[3483] = 25'b0000000000000010011011000;
    rom[3484] = 25'b0000000000000010011011001;
    rom[3485] = 25'b0000000000000010011011011;
    rom[3486] = 25'b0000000000000010011011100;
    rom[3487] = 25'b0000000000000010011011110;
    rom[3488] = 25'b0000000000000010011011111;
    rom[3489] = 25'b0000000000000010011100000;
    rom[3490] = 25'b0000000000000010011100001;
    rom[3491] = 25'b0000000000000010011100011;
    rom[3492] = 25'b0000000000000010011100100;
    rom[3493] = 25'b0000000000000010011100110;
    rom[3494] = 25'b0000000000000010011100111;
    rom[3495] = 25'b0000000000000010011101001;
    rom[3496] = 25'b0000000000000010011101010;
    rom[3497] = 25'b0000000000000010011101100;
    rom[3498] = 25'b0000000000000010011101101;
    rom[3499] = 25'b0000000000000010011101111;
    rom[3500] = 25'b0000000000000010011110000;
    rom[3501] = 25'b0000000000000010011110010;
    rom[3502] = 25'b0000000000000010011110011;
    rom[3503] = 25'b0000000000000010011110100;
    rom[3504] = 25'b0000000000000010011110110;
    rom[3505] = 25'b0000000000000010011110111;
    rom[3506] = 25'b0000000000000010011111001;
    rom[3507] = 25'b0000000000000010011111010;
    rom[3508] = 25'b0000000000000010011111100;
    rom[3509] = 25'b0000000000000010011111101;
    rom[3510] = 25'b0000000000000010011111111;
    rom[3511] = 25'b0000000000000010100000000;
    rom[3512] = 25'b0000000000000010100000010;
    rom[3513] = 25'b0000000000000010100000010;
    rom[3514] = 25'b0000000000000010100000100;
    rom[3515] = 25'b0000000000000010100000101;
    rom[3516] = 25'b0000000000000010100000111;
    rom[3517] = 25'b0000000000000010100001000;
    rom[3518] = 25'b0000000000000010100001010;
    rom[3519] = 25'b0000000000000010100001011;
    rom[3520] = 25'b0000000000000010100001101;
    rom[3521] = 25'b0000000000000010100001110;
    rom[3522] = 25'b0000000000000010100010000;
    rom[3523] = 25'b0000000000000010100010000;
    rom[3524] = 25'b0000000000000010100010010;
    rom[3525] = 25'b0000000000000010100010011;
    rom[3526] = 25'b0000000000000010100010101;
    rom[3527] = 25'b0000000000000010100010110;
    rom[3528] = 25'b0000000000000010100011000;
    rom[3529] = 25'b0000000000000010100011001;
    rom[3530] = 25'b0000000000000010100011011;
    rom[3531] = 25'b0000000000000010100011100;
    rom[3532] = 25'b0000000000000010100011101;
    rom[3533] = 25'b0000000000000010100011111;
    rom[3534] = 25'b0000000000000010100100000;
    rom[3535] = 25'b0000000000000010100100010;
    rom[3536] = 25'b0000000000000010100100011;
    rom[3537] = 25'b0000000000000010100100101;
    rom[3538] = 25'b0000000000000010100100110;
    rom[3539] = 25'b0000000000000010100101000;
    rom[3540] = 25'b0000000000000010100101000;
    rom[3541] = 25'b0000000000000010100101010;
    rom[3542] = 25'b0000000000000010100101011;
    rom[3543] = 25'b0000000000000010100101101;
    rom[3544] = 25'b0000000000000010100101110;
    rom[3545] = 25'b0000000000000010100110000;
    rom[3546] = 25'b0000000000000010100110001;
    rom[3547] = 25'b0000000000000010100110011;
    rom[3548] = 25'b0000000000000010100110100;
    rom[3549] = 25'b0000000000000010100110101;
    rom[3550] = 25'b0000000000000010100110111;
    rom[3551] = 25'b0000000000000010100111000;
    rom[3552] = 25'b0000000000000010100111010;
    rom[3553] = 25'b0000000000000010100111011;
    rom[3554] = 25'b0000000000000010100111101;
    rom[3555] = 25'b0000000000000010100111110;
    rom[3556] = 25'b0000000000000010100111111;
    rom[3557] = 25'b0000000000000010101000000;
    rom[3558] = 25'b0000000000000010101000010;
    rom[3559] = 25'b0000000000000010101000011;
    rom[3560] = 25'b0000000000000010101000101;
    rom[3561] = 25'b0000000000000010101000110;
    rom[3562] = 25'b0000000000000010101001000;
    rom[3563] = 25'b0000000000000010101001000;
    rom[3564] = 25'b0000000000000010101001010;
    rom[3565] = 25'b0000000000000010101001011;
    rom[3566] = 25'b0000000000000010101001101;
    rom[3567] = 25'b0000000000000010101001110;
    rom[3568] = 25'b0000000000000010101010000;
    rom[3569] = 25'b0000000000000010101010001;
    rom[3570] = 25'b0000000000000010101010010;
    rom[3571] = 25'b0000000000000010101010100;
    rom[3572] = 25'b0000000000000010101010101;
    rom[3573] = 25'b0000000000000010101010111;
    rom[3574] = 25'b0000000000000010101011000;
    rom[3575] = 25'b0000000000000010101011010;
    rom[3576] = 25'b0000000000000010101011010;
    rom[3577] = 25'b0000000000000010101011100;
    rom[3578] = 25'b0000000000000010101011101;
    rom[3579] = 25'b0000000000000010101011111;
    rom[3580] = 25'b0000000000000010101100000;
    rom[3581] = 25'b0000000000000010101100010;
    rom[3582] = 25'b0000000000000010101100011;
    rom[3583] = 25'b0000000000000010101100100;
    rom[3584] = 25'b0000000000000010101100110;
    rom[3585] = 25'b0000000000000010101100111;
    rom[3586] = 25'b0000000000000010101101001;
    rom[3587] = 25'b0000000000000010101101010;
    rom[3588] = 25'b0000000000000010101101011;
    rom[3589] = 25'b0000000000000010101101100;
    rom[3590] = 25'b0000000000000010101101110;
    rom[3591] = 25'b0000000000000010101101111;
    rom[3592] = 25'b0000000000000010101110001;
    rom[3593] = 25'b0000000000000010101110010;
    rom[3594] = 25'b0000000000000010101110011;
    rom[3595] = 25'b0000000000000010101110101;
    rom[3596] = 25'b0000000000000010101110110;
    rom[3597] = 25'b0000000000000010101111000;
    rom[3598] = 25'b0000000000000010101111001;
    rom[3599] = 25'b0000000000000010101111010;
    rom[3600] = 25'b0000000000000010101111011;
    rom[3601] = 25'b0000000000000010101111101;
    rom[3602] = 25'b0000000000000010101111110;
    rom[3603] = 25'b0000000000000010110000000;
    rom[3604] = 25'b0000000000000010110000001;
    rom[3605] = 25'b0000000000000010110000010;
    rom[3606] = 25'b0000000000000010110000100;
    rom[3607] = 25'b0000000000000010110000101;
    rom[3608] = 25'b0000000000000010110000111;
    rom[3609] = 25'b0000000000000010110000111;
    rom[3610] = 25'b0000000000000010110001001;
    rom[3611] = 25'b0000000000000010110001010;
    rom[3612] = 25'b0000000000000010110001100;
    rom[3613] = 25'b0000000000000010110001101;
    rom[3614] = 25'b0000000000000010110001110;
    rom[3615] = 25'b0000000000000010110001111;
    rom[3616] = 25'b0000000000000010110010001;
    rom[3617] = 25'b0000000000000010110010010;
    rom[3618] = 25'b0000000000000010110010011;
    rom[3619] = 25'b0000000000000010110010101;
    rom[3620] = 25'b0000000000000010110010110;
    rom[3621] = 25'b0000000000000010110011000;
    rom[3622] = 25'b0000000000000010110011001;
    rom[3623] = 25'b0000000000000010110011010;
    rom[3624] = 25'b0000000000000010110011011;
    rom[3625] = 25'b0000000000000010110011101;
    rom[3626] = 25'b0000000000000010110011110;
    rom[3627] = 25'b0000000000000010110011111;
    rom[3628] = 25'b0000000000000010110100001;
    rom[3629] = 25'b0000000000000010110100010;
    rom[3630] = 25'b0000000000000010110100100;
    rom[3631] = 25'b0000000000000010110100101;
    rom[3632] = 25'b0000000000000010110100110;
    rom[3633] = 25'b0000000000000010110100111;
    rom[3634] = 25'b0000000000000010110101001;
    rom[3635] = 25'b0000000000000010110101010;
    rom[3636] = 25'b0000000000000010110101011;
    rom[3637] = 25'b0000000000000010110101101;
    rom[3638] = 25'b0000000000000010110101110;
    rom[3639] = 25'b0000000000000010110110000;
    rom[3640] = 25'b0000000000000010110110000;
    rom[3641] = 25'b0000000000000010110110010;
    rom[3642] = 25'b0000000000000010110110011;
    rom[3643] = 25'b0000000000000010110110101;
    rom[3644] = 25'b0000000000000010110110110;
    rom[3645] = 25'b0000000000000010110110111;
    rom[3646] = 25'b0000000000000010110111001;
    rom[3647] = 25'b0000000000000010110111010;
    rom[3648] = 25'b0000000000000010110111011;
    rom[3649] = 25'b0000000000000010110111100;
    rom[3650] = 25'b0000000000000010110111110;
    rom[3651] = 25'b0000000000000010110111111;
    rom[3652] = 25'b0000000000000010111000000;
    rom[3653] = 25'b0000000000000010111000010;
    rom[3654] = 25'b0000000000000010111000011;
    rom[3655] = 25'b0000000000000010111000101;
    rom[3656] = 25'b0000000000000010111000101;
    rom[3657] = 25'b0000000000000010111000111;
    rom[3658] = 25'b0000000000000010111001000;
    rom[3659] = 25'b0000000000000010111001010;
    rom[3660] = 25'b0000000000000010111001010;
    rom[3661] = 25'b0000000000000010111001100;
    rom[3662] = 25'b0000000000000010111001101;
    rom[3663] = 25'b0000000000000010111001110;
    rom[3664] = 25'b0000000000000010111010000;
    rom[3665] = 25'b0000000000000010111010001;
    rom[3666] = 25'b0000000000000010111010011;
    rom[3667] = 25'b0000000000000010111010011;
    rom[3668] = 25'b0000000000000010111010101;
    rom[3669] = 25'b0000000000000010111010110;
    rom[3670] = 25'b0000000000000010111010111;
    rom[3671] = 25'b0000000000000010111011001;
    rom[3672] = 25'b0000000000000010111011010;
    rom[3673] = 25'b0000000000000010111011100;
    rom[3674] = 25'b0000000000000010111011100;
    rom[3675] = 25'b0000000000000010111011110;
    rom[3676] = 25'b0000000000000010111011111;
    rom[3677] = 25'b0000000000000010111100000;
    rom[3678] = 25'b0000000000000010111100010;
    rom[3679] = 25'b0000000000000010111100011;
    rom[3680] = 25'b0000000000000010111100100;
    rom[3681] = 25'b0000000000000010111100101;
    rom[3682] = 25'b0000000000000010111100111;
    rom[3683] = 25'b0000000000000010111101000;
    rom[3684] = 25'b0000000000000010111101001;
    rom[3685] = 25'b0000000000000010111101011;
    rom[3686] = 25'b0000000000000010111101100;
    rom[3687] = 25'b0000000000000010111101101;
    rom[3688] = 25'b0000000000000010111101110;
    rom[3689] = 25'b0000000000000010111110000;
    rom[3690] = 25'b0000000000000010111110001;
    rom[3691] = 25'b0000000000000010111110010;
    rom[3692] = 25'b0000000000000010111110100;
    rom[3693] = 25'b0000000000000010111110100;
    rom[3694] = 25'b0000000000000010111110110;
    rom[3695] = 25'b0000000000000010111110111;
    rom[3696] = 25'b0000000000000010111111000;
    rom[3697] = 25'b0000000000000010111111010;
    rom[3698] = 25'b0000000000000010111111011;
    rom[3699] = 25'b0000000000000010111111100;
    rom[3700] = 25'b0000000000000010111111101;
    rom[3701] = 25'b0000000000000010111111111;
    rom[3702] = 25'b0000000000000011000000000;
    rom[3703] = 25'b0000000000000011000000001;
    rom[3704] = 25'b0000000000000011000000011;
    rom[3705] = 25'b0000000000000011000000011;
    rom[3706] = 25'b0000000000000011000000101;
    rom[3707] = 25'b0000000000000011000000110;
    rom[3708] = 25'b0000000000000011000000111;
    rom[3709] = 25'b0000000000000011000001000;
    rom[3710] = 25'b0000000000000011000001010;
    rom[3711] = 25'b0000000000000011000001011;
    rom[3712] = 25'b0000000000000011000001100;
    rom[3713] = 25'b0000000000000011000001110;
    rom[3714] = 25'b0000000000000011000001110;
    rom[3715] = 25'b0000000000000011000010000;
    rom[3716] = 25'b0000000000000011000010001;
    rom[3717] = 25'b0000000000000011000010010;
    rom[3718] = 25'b0000000000000011000010100;
    rom[3719] = 25'b0000000000000011000010100;
    rom[3720] = 25'b0000000000000011000010110;
    rom[3721] = 25'b0000000000000011000010111;
    rom[3722] = 25'b0000000000000011000011000;
    rom[3723] = 25'b0000000000000011000011010;
    rom[3724] = 25'b0000000000000011000011010;
    rom[3725] = 25'b0000000000000011000011100;
    rom[3726] = 25'b0000000000000011000011101;
    rom[3727] = 25'b0000000000000011000011110;
    rom[3728] = 25'b0000000000000011000100000;
    rom[3729] = 25'b0000000000000011000100001;
    rom[3730] = 25'b0000000000000011000100010;
    rom[3731] = 25'b0000000000000011000100011;
    rom[3732] = 25'b0000000000000011000100100;
    rom[3733] = 25'b0000000000000011000100110;
    rom[3734] = 25'b0000000000000011000100111;
    rom[3735] = 25'b0000000000000011000101000;
    rom[3736] = 25'b0000000000000011000101001;
    rom[3737] = 25'b0000000000000011000101010;
    rom[3738] = 25'b0000000000000011000101100;
    rom[3739] = 25'b0000000000000011000101101;
    rom[3740] = 25'b0000000000000011000101110;
    rom[3741] = 25'b0000000000000011000101111;
    rom[3742] = 25'b0000000000000011000110000;
    rom[3743] = 25'b0000000000000011000110010;
    rom[3744] = 25'b0000000000000011000110011;
    rom[3745] = 25'b0000000000000011000110100;
    rom[3746] = 25'b0000000000000011000110101;
    rom[3747] = 25'b0000000000000011000110110;
    rom[3748] = 25'b0000000000000011000111000;
    rom[3749] = 25'b0000000000000011000111000;
    rom[3750] = 25'b0000000000000011000111010;
    rom[3751] = 25'b0000000000000011000111011;
    rom[3752] = 25'b0000000000000011000111100;
    rom[3753] = 25'b0000000000000011000111110;
    rom[3754] = 25'b0000000000000011000111110;
    rom[3755] = 25'b0000000000000011001000000;
    rom[3756] = 25'b0000000000000011001000001;
    rom[3757] = 25'b0000000000000011001000010;
    rom[3758] = 25'b0000000000000011001000100;
    rom[3759] = 25'b0000000000000011001000100;
    rom[3760] = 25'b0000000000000011001000110;
    rom[3761] = 25'b0000000000000011001000111;
    rom[3762] = 25'b0000000000000011001001000;
    rom[3763] = 25'b0000000000000011001001001;
    rom[3764] = 25'b0000000000000011001001010;
    rom[3765] = 25'b0000000000000011001001011;
    rom[3766] = 25'b0000000000000011001001100;
    rom[3767] = 25'b0000000000000011001001101;
    rom[3768] = 25'b0000000000000011001001111;
    rom[3769] = 25'b0000000000000011001010000;
    rom[3770] = 25'b0000000000000011001010001;
    rom[3771] = 25'b0000000000000011001010010;
    rom[3772] = 25'b0000000000000011001010011;
    rom[3773] = 25'b0000000000000011001010101;
    rom[3774] = 25'b0000000000000011001010101;
    rom[3775] = 25'b0000000000000011001010111;
    rom[3776] = 25'b0000000000000011001011000;
    rom[3777] = 25'b0000000000000011001011001;
    rom[3778] = 25'b0000000000000011001011010;
    rom[3779] = 25'b0000000000000011001011011;
    rom[3780] = 25'b0000000000000011001011100;
    rom[3781] = 25'b0000000000000011001011110;
    rom[3782] = 25'b0000000000000011001011110;
    rom[3783] = 25'b0000000000000011001100000;
    rom[3784] = 25'b0000000000000011001100001;
    rom[3785] = 25'b0000000000000011001100010;
    rom[3786] = 25'b0000000000000011001100011;
    rom[3787] = 25'b0000000000000011001100100;
    rom[3788] = 25'b0000000000000011001100101;
    rom[3789] = 25'b0000000000000011001100111;
    rom[3790] = 25'b0000000000000011001100111;
    rom[3791] = 25'b0000000000000011001101001;
    rom[3792] = 25'b0000000000000011001101010;
    rom[3793] = 25'b0000000000000011001101011;
    rom[3794] = 25'b0000000000000011001101100;
    rom[3795] = 25'b0000000000000011001101101;
    rom[3796] = 25'b0000000000000011001101110;
    rom[3797] = 25'b0000000000000011001110000;
    rom[3798] = 25'b0000000000000011001110000;
    rom[3799] = 25'b0000000000000011001110010;
    rom[3800] = 25'b0000000000000011001110011;
    rom[3801] = 25'b0000000000000011001110100;
    rom[3802] = 25'b0000000000000011001110101;
    rom[3803] = 25'b0000000000000011001110110;
    rom[3804] = 25'b0000000000000011001110111;
    rom[3805] = 25'b0000000000000011001111001;
    rom[3806] = 25'b0000000000000011001111001;
    rom[3807] = 25'b0000000000000011001111011;
    rom[3808] = 25'b0000000000000011001111100;
    rom[3809] = 25'b0000000000000011001111100;
    rom[3810] = 25'b0000000000000011001111110;
    rom[3811] = 25'b0000000000000011001111111;
    rom[3812] = 25'b0000000000000011010000000;
    rom[3813] = 25'b0000000000000011010000001;
    rom[3814] = 25'b0000000000000011010000010;
    rom[3815] = 25'b0000000000000011010000011;
    rom[3816] = 25'b0000000000000011010000101;
    rom[3817] = 25'b0000000000000011010000101;
    rom[3818] = 25'b0000000000000011010000111;
    rom[3819] = 25'b0000000000000011010001000;
    rom[3820] = 25'b0000000000000011010001000;
    rom[3821] = 25'b0000000000000011010001010;
    rom[3822] = 25'b0000000000000011010001010;
    rom[3823] = 25'b0000000000000011010001100;
    rom[3824] = 25'b0000000000000011010001101;
    rom[3825] = 25'b0000000000000011010001110;
    rom[3826] = 25'b0000000000000011010001111;
    rom[3827] = 25'b0000000000000011010010000;
    rom[3828] = 25'b0000000000000011010010001;
    rom[3829] = 25'b0000000000000011010010010;
    rom[3830] = 25'b0000000000000011010010011;
    rom[3831] = 25'b0000000000000011010010100;
    rom[3832] = 25'b0000000000000011010010101;
    rom[3833] = 25'b0000000000000011010010110;
    rom[3834] = 25'b0000000000000011010010111;
    rom[3835] = 25'b0000000000000011010011001;
    rom[3836] = 25'b0000000000000011010011001;
    rom[3837] = 25'b0000000000000011010011010;
    rom[3838] = 25'b0000000000000011010011100;
    rom[3839] = 25'b0000000000000011010011100;
    rom[3840] = 25'b0000000000000011010011110;
    rom[3841] = 25'b0000000000000011010011111;
    rom[3842] = 25'b0000000000000011010011111;
    rom[3843] = 25'b0000000000000011010100001;
    rom[3844] = 25'b0000000000000011010100010;
    rom[3845] = 25'b0000000000000011010100011;
    rom[3846] = 25'b0000000000000011010100100;
    rom[3847] = 25'b0000000000000011010100101;
    rom[3848] = 25'b0000000000000011010100110;
    rom[3849] = 25'b0000000000000011010100111;
    rom[3850] = 25'b0000000000000011010101000;
    rom[3851] = 25'b0000000000000011010101001;
    rom[3852] = 25'b0000000000000011010101010;
    rom[3853] = 25'b0000000000000011010101011;
    rom[3854] = 25'b0000000000000011010101100;
    rom[3855] = 25'b0000000000000011010101101;
    rom[3856] = 25'b0000000000000011010101110;
    rom[3857] = 25'b0000000000000011010101111;
    rom[3858] = 25'b0000000000000011010110000;
    rom[3859] = 25'b0000000000000011010110001;
    rom[3860] = 25'b0000000000000011010110010;
    rom[3861] = 25'b0000000000000011010110011;
    rom[3862] = 25'b0000000000000011010110100;
    rom[3863] = 25'b0000000000000011010110101;
    rom[3864] = 25'b0000000000000011010110110;
    rom[3865] = 25'b0000000000000011010110111;
    rom[3866] = 25'b0000000000000011010111000;
    rom[3867] = 25'b0000000000000011010111001;
    rom[3868] = 25'b0000000000000011010111010;
    rom[3869] = 25'b0000000000000011010111011;
    rom[3870] = 25'b0000000000000011010111100;
    rom[3871] = 25'b0000000000000011010111101;
    rom[3872] = 25'b0000000000000011010111110;
    rom[3873] = 25'b0000000000000011010111111;
    rom[3874] = 25'b0000000000000011011000000;
    rom[3875] = 25'b0000000000000011011000001;
    rom[3876] = 25'b0000000000000011011000010;
    rom[3877] = 25'b0000000000000011011000011;
    rom[3878] = 25'b0000000000000011011000100;
    rom[3879] = 25'b0000000000000011011000101;
    rom[3880] = 25'b0000000000000011011000110;
    rom[3881] = 25'b0000000000000011011000111;
    rom[3882] = 25'b0000000000000011011001000;
    rom[3883] = 25'b0000000000000011011001000;
    rom[3884] = 25'b0000000000000011011001010;
    rom[3885] = 25'b0000000000000011011001011;
    rom[3886] = 25'b0000000000000011011001011;
    rom[3887] = 25'b0000000000000011011001100;
    rom[3888] = 25'b0000000000000011011001110;
    rom[3889] = 25'b0000000000000011011001110;
    rom[3890] = 25'b0000000000000011011001111;
    rom[3891] = 25'b0000000000000011011010000;
    rom[3892] = 25'b0000000000000011011010001;
    rom[3893] = 25'b0000000000000011011010010;
    rom[3894] = 25'b0000000000000011011010011;
    rom[3895] = 25'b0000000000000011011010100;
    rom[3896] = 25'b0000000000000011011010101;
    rom[3897] = 25'b0000000000000011011010110;
    rom[3898] = 25'b0000000000000011011010111;
    rom[3899] = 25'b0000000000000011011011000;
    rom[3900] = 25'b0000000000000011011011001;
    rom[3901] = 25'b0000000000000011011011010;
    rom[3902] = 25'b0000000000000011011011010;
    rom[3903] = 25'b0000000000000011011011100;
    rom[3904] = 25'b0000000000000011011011101;
    rom[3905] = 25'b0000000000000011011011101;
    rom[3906] = 25'b0000000000000011011011110;
    rom[3907] = 25'b0000000000000011011011111;
    rom[3908] = 25'b0000000000000011011100000;
    rom[3909] = 25'b0000000000000011011100001;
    rom[3910] = 25'b0000000000000011011100010;
    rom[3911] = 25'b0000000000000011011100011;
    rom[3912] = 25'b0000000000000011011100100;
    rom[3913] = 25'b0000000000000011011100101;
    rom[3914] = 25'b0000000000000011011100110;
    rom[3915] = 25'b0000000000000011011100110;
    rom[3916] = 25'b0000000000000011011100111;
    rom[3917] = 25'b0000000000000011011101001;
    rom[3918] = 25'b0000000000000011011101001;
    rom[3919] = 25'b0000000000000011011101010;
    rom[3920] = 25'b0000000000000011011101011;
    rom[3921] = 25'b0000000000000011011101100;
    rom[3922] = 25'b0000000000000011011101101;
    rom[3923] = 25'b0000000000000011011101110;
    rom[3924] = 25'b0000000000000011011101111;
    rom[3925] = 25'b0000000000000011011101111;
    rom[3926] = 25'b0000000000000011011110000;
    rom[3927] = 25'b0000000000000011011110010;
    rom[3928] = 25'b0000000000000011011110010;
    rom[3929] = 25'b0000000000000011011110011;
    rom[3930] = 25'b0000000000000011011110100;
    rom[3931] = 25'b0000000000000011011110101;
    rom[3932] = 25'b0000000000000011011110101;
    rom[3933] = 25'b0000000000000011011110111;
    rom[3934] = 25'b0000000000000011011111000;
    rom[3935] = 25'b0000000000000011011111000;
    rom[3936] = 25'b0000000000000011011111001;
    rom[3937] = 25'b0000000000000011011111010;
    rom[3938] = 25'b0000000000000011011111011;
    rom[3939] = 25'b0000000000000011011111100;
    rom[3940] = 25'b0000000000000011011111101;
    rom[3941] = 25'b0000000000000011011111110;
    rom[3942] = 25'b0000000000000011011111110;
    rom[3943] = 25'b0000000000000011011111111;
    rom[3944] = 25'b0000000000000011100000000;
    rom[3945] = 25'b0000000000000011100000001;
    rom[3946] = 25'b0000000000000011100000001;
    rom[3947] = 25'b0000000000000011100000011;
    rom[3948] = 25'b0000000000000011100000100;
    rom[3949] = 25'b0000000000000011100000100;
    rom[3950] = 25'b0000000000000011100000101;
    rom[3951] = 25'b0000000000000011100000110;
    rom[3952] = 25'b0000000000000011100000111;
    rom[3953] = 25'b0000000000000011100000111;
    rom[3954] = 25'b0000000000000011100001000;
    rom[3955] = 25'b0000000000000011100001001;
    rom[3956] = 25'b0000000000000011100001010;
    rom[3957] = 25'b0000000000000011100001011;
    rom[3958] = 25'b0000000000000011100001100;
    rom[3959] = 25'b0000000000000011100001100;
    rom[3960] = 25'b0000000000000011100001101;
    rom[3961] = 25'b0000000000000011100001110;
    rom[3962] = 25'b0000000000000011100001111;
    rom[3963] = 25'b0000000000000011100001111;
    rom[3964] = 25'b0000000000000011100010000;
    rom[3965] = 25'b0000000000000011100010001;
    rom[3966] = 25'b0000000000000011100010010;
    rom[3967] = 25'b0000000000000011100010011;
    rom[3968] = 25'b0000000000000011100010100;
    rom[3969] = 25'b0000000000000011100010101;
    rom[3970] = 25'b0000000000000011100010101;
    rom[3971] = 25'b0000000000000011100010110;
    rom[3972] = 25'b0000000000000011100010111;
    rom[3973] = 25'b0000000000000011100011000;
    rom[3974] = 25'b0000000000000011100011000;
    rom[3975] = 25'b0000000000000011100011001;
    rom[3976] = 25'b0000000000000011100011010;
    rom[3977] = 25'b0000000000000011100011011;
    rom[3978] = 25'b0000000000000011100011011;
    rom[3979] = 25'b0000000000000011100011100;
    rom[3980] = 25'b0000000000000011100011101;
    rom[3981] = 25'b0000000000000011100011110;
    rom[3982] = 25'b0000000000000011100011110;
    rom[3983] = 25'b0000000000000011100011111;
    rom[3984] = 25'b0000000000000011100100000;
    rom[3985] = 25'b0000000000000011100100001;
    rom[3986] = 25'b0000000000000011100100001;
    rom[3987] = 25'b0000000000000011100100011;
    rom[3988] = 25'b0000000000000011100100100;
    rom[3989] = 25'b0000000000000011100100100;
    rom[3990] = 25'b0000000000000011100100101;
    rom[3991] = 25'b0000000000000011100100110;
    rom[3992] = 25'b0000000000000011100100111;
    rom[3993] = 25'b0000000000000011100100111;
    rom[3994] = 25'b0000000000000011100101000;
    rom[3995] = 25'b0000000000000011100101001;
    rom[3996] = 25'b0000000000000011100101010;
    rom[3997] = 25'b0000000000000011100101010;
    rom[3998] = 25'b0000000000000011100101011;
    rom[3999] = 25'b0000000000000011100101100;
    rom[4000] = 25'b0000000000000011100101100;
    rom[4001] = 25'b0000000000000011100101101;
    rom[4002] = 25'b0000000000000011100101101;
    rom[4003] = 25'b0000000000000011100101110;
    rom[4004] = 25'b0000000000000011100101111;
    rom[4005] = 25'b0000000000000011100110000;
    rom[4006] = 25'b0000000000000011100110000;
    rom[4007] = 25'b0000000000000011100110001;
    rom[4008] = 25'b0000000000000011100110010;
    rom[4009] = 25'b0000000000000011100110011;
    rom[4010] = 25'b0000000000000011100110011;
    rom[4011] = 25'b0000000000000011100110100;
    rom[4012] = 25'b0000000000000011100110101;
    rom[4013] = 25'b0000000000000011100110110;
    rom[4014] = 25'b0000000000000011100110110;
    rom[4015] = 25'b0000000000000011100110111;
    rom[4016] = 25'b0000000000000011100111000;
    rom[4017] = 25'b0000000000000011100111001;
    rom[4018] = 25'b0000000000000011100111001;
    rom[4019] = 25'b0000000000000011100111010;
    rom[4020] = 25'b0000000000000011100111010;
    rom[4021] = 25'b0000000000000011100111011;
    rom[4022] = 25'b0000000000000011100111100;
    rom[4023] = 25'b0000000000000011100111100;
    rom[4024] = 25'b0000000000000011100111101;
    rom[4025] = 25'b0000000000000011100111110;
    rom[4026] = 25'b0000000000000011100111111;
    rom[4027] = 25'b0000000000000011100111111;
    rom[4028] = 25'b0000000000000011101000000;
    rom[4029] = 25'b0000000000000011101000001;
    rom[4030] = 25'b0000000000000011101000010;
    rom[4031] = 25'b0000000000000011101000010;
    rom[4032] = 25'b0000000000000011101000010;
    rom[4033] = 25'b0000000000000011101000011;
    rom[4034] = 25'b0000000000000011101000100;
    rom[4035] = 25'b0000000000000011101000101;
    rom[4036] = 25'b0000000000000011101000101;
    rom[4037] = 25'b0000000000000011101000110;
    rom[4038] = 25'b0000000000000011101000111;
    rom[4039] = 25'b0000000000000011101000111;
    rom[4040] = 25'b0000000000000011101001000;
    rom[4041] = 25'b0000000000000011101001000;
    rom[4042] = 25'b0000000000000011101001001;
    rom[4043] = 25'b0000000000000011101001010;
    rom[4044] = 25'b0000000000000011101001010;
    rom[4045] = 25'b0000000000000011101001011;
    rom[4046] = 25'b0000000000000011101001011;
    rom[4047] = 25'b0000000000000011101001100;
    rom[4048] = 25'b0000000000000011101001101;
    rom[4049] = 25'b0000000000000011101001101;
    rom[4050] = 25'b0000000000000011101001110;
    rom[4051] = 25'b0000000000000011101001111;
    rom[4052] = 25'b0000000000000011101001111;
    rom[4053] = 25'b0000000000000011101010000;
    rom[4054] = 25'b0000000000000011101010000;
    rom[4055] = 25'b0000000000000011101010001;
    rom[4056] = 25'b0000000000000011101010010;
    rom[4057] = 25'b0000000000000011101010011;
    rom[4058] = 25'b0000000000000011101010011;
    rom[4059] = 25'b0000000000000011101010011;
    rom[4060] = 25'b0000000000000011101010100;
    rom[4061] = 25'b0000000000000011101010101;
    rom[4062] = 25'b0000000000000011101010110;
    rom[4063] = 25'b0000000000000011101010110;
    rom[4064] = 25'b0000000000000011101010110;
    rom[4065] = 25'b0000000000000011101010111;
    rom[4066] = 25'b0000000000000011101011000;
    rom[4067] = 25'b0000000000000011101011000;
    rom[4068] = 25'b0000000000000011101011001;
    rom[4069] = 25'b0000000000000011101011001;
    rom[4070] = 25'b0000000000000011101011010;
    rom[4071] = 25'b0000000000000011101011011;
    rom[4072] = 25'b0000000000000011101011011;
    rom[4073] = 25'b0000000000000011101011100;
    rom[4074] = 25'b0000000000000011101011100;
    rom[4075] = 25'b0000000000000011101011101;
    rom[4076] = 25'b0000000000000011101011101;
    rom[4077] = 25'b0000000000000011101011110;
    rom[4078] = 25'b0000000000000011101011111;
    rom[4079] = 25'b0000000000000011101011111;
    rom[4080] = 25'b0000000000000011101011111;
    rom[4081] = 25'b0000000000000011101100000;
    rom[4082] = 25'b0000000000000011101100001;
    rom[4083] = 25'b0000000000000011101100001;
    rom[4084] = 25'b0000000000000011101100010;
    rom[4085] = 25'b0000000000000011101100010;
    rom[4086] = 25'b0000000000000011101100011;
    rom[4087] = 25'b0000000000000011101100011;
    rom[4088] = 25'b0000000000000011101100100;
    rom[4089] = 25'b0000000000000011101100101;
    rom[4090] = 25'b0000000000000011101100101;
    rom[4091] = 25'b0000000000000011101100101;
    rom[4092] = 25'b0000000000000011101100110;
    rom[4093] = 25'b0000000000000011101100111;
    rom[4094] = 25'b0000000000000011101100111;
    rom[4095] = 25'b0000000000000011101101000;
    rom[4096] = 25'b0000000000000011101101000;
    rom[4097] = 25'b0000000000000011101101000;
    rom[4098] = 25'b0000000000000011101101001;
    rom[4099] = 25'b0000000000000011101101010;
    rom[4100] = 25'b0000000000000011101101010;
    rom[4101] = 25'b0000000000000011101101011;
    rom[4102] = 25'b0000000000000011101101011;
    rom[4103] = 25'b0000000000000011101101011;
    rom[4104] = 25'b0000000000000011101101100;
    rom[4105] = 25'b0000000000000011101101101;
    rom[4106] = 25'b0000000000000011101101101;
    rom[4107] = 25'b0000000000000011101101110;
    rom[4108] = 25'b0000000000000011101101110;
    rom[4109] = 25'b0000000000000011101101110;
    rom[4110] = 25'b0000000000000011101101111;
    rom[4111] = 25'b0000000000000011101110000;
    rom[4112] = 25'b0000000000000011101110000;
    rom[4113] = 25'b0000000000000011101110001;
    rom[4114] = 25'b0000000000000011101110001;
    rom[4115] = 25'b0000000000000011101110001;
    rom[4116] = 25'b0000000000000011101110010;
    rom[4117] = 25'b0000000000000011101110010;
    rom[4118] = 25'b0000000000000011101110011;
    rom[4119] = 25'b0000000000000011101110100;
    rom[4120] = 25'b0000000000000011101110100;
    rom[4121] = 25'b0000000000000011101110100;
    rom[4122] = 25'b0000000000000011101110100;
    rom[4123] = 25'b0000000000000011101110101;
    rom[4124] = 25'b0000000000000011101110110;
    rom[4125] = 25'b0000000000000011101110110;
    rom[4126] = 25'b0000000000000011101110111;
    rom[4127] = 25'b0000000000000011101110111;
    rom[4128] = 25'b0000000000000011101110111;
    rom[4129] = 25'b0000000000000011101110111;
    rom[4130] = 25'b0000000000000011101111000;
    rom[4131] = 25'b0000000000000011101111001;
    rom[4132] = 25'b0000000000000011101111001;
    rom[4133] = 25'b0000000000000011101111010;
    rom[4134] = 25'b0000000000000011101111010;
    rom[4135] = 25'b0000000000000011101111010;
    rom[4136] = 25'b0000000000000011101111010;
    rom[4137] = 25'b0000000000000011101111011;
    rom[4138] = 25'b0000000000000011101111011;
    rom[4139] = 25'b0000000000000011101111100;
    rom[4140] = 25'b0000000000000011101111101;
    rom[4141] = 25'b0000000000000011101111101;
    rom[4142] = 25'b0000000000000011101111101;
    rom[4143] = 25'b0000000000000011101111101;
    rom[4144] = 25'b0000000000000011101111110;
    rom[4145] = 25'b0000000000000011101111110;
    rom[4146] = 25'b0000000000000011101111111;
    rom[4147] = 25'b0000000000000011101111111;
    rom[4148] = 25'b0000000000000011110000000;
    rom[4149] = 25'b0000000000000011110000000;
    rom[4150] = 25'b0000000000000011110000000;
    rom[4151] = 25'b0000000000000011110000000;
    rom[4152] = 25'b0000000000000011110000001;
    rom[4153] = 25'b0000000000000011110000001;
    rom[4154] = 25'b0000000000000011110000010;
    rom[4155] = 25'b0000000000000011110000010;
    rom[4156] = 25'b0000000000000011110000011;
    rom[4157] = 25'b0000000000000011110000011;
    rom[4158] = 25'b0000000000000011110000011;
    rom[4159] = 25'b0000000000000011110000011;
    rom[4160] = 25'b0000000000000011110000100;
    rom[4161] = 25'b0000000000000011110000100;
    rom[4162] = 25'b0000000000000011110000101;
    rom[4163] = 25'b0000000000000011110000101;
    rom[4164] = 25'b0000000000000011110000101;
    rom[4165] = 25'b0000000000000011110000110;
    rom[4166] = 25'b0000000000000011110000110;
    rom[4167] = 25'b0000000000000011110000110;
    rom[4168] = 25'b0000000000000011110000110;
    rom[4169] = 25'b0000000000000011110000111;
    rom[4170] = 25'b0000000000000011110000111;
    rom[4171] = 25'b0000000000000011110001000;
    rom[4172] = 25'b0000000000000011110001000;
    rom[4173] = 25'b0000000000000011110001000;
    rom[4174] = 25'b0000000000000011110001001;
    rom[4175] = 25'b0000000000000011110001001;
    rom[4176] = 25'b0000000000000011110001001;
    rom[4177] = 25'b0000000000000011110001001;
    rom[4178] = 25'b0000000000000011110001001;
    rom[4179] = 25'b0000000000000011110001010;
    rom[4180] = 25'b0000000000000011110001010;
    rom[4181] = 25'b0000000000000011110001011;
    rom[4182] = 25'b0000000000000011110001011;
    rom[4183] = 25'b0000000000000011110001011;
    rom[4184] = 25'b0000000000000011110001011;
    rom[4185] = 25'b0000000000000011110001011;
    rom[4186] = 25'b0000000000000011110001100;
    rom[4187] = 25'b0000000000000011110001100;
    rom[4188] = 25'b0000000000000011110001100;
    rom[4189] = 25'b0000000000000011110001101;
    rom[4190] = 25'b0000000000000011110001101;
    rom[4191] = 25'b0000000000000011110001101;
    rom[4192] = 25'b0000000000000011110001110;
    rom[4193] = 25'b0000000000000011110001110;
    rom[4194] = 25'b0000000000000011110001110;
    rom[4195] = 25'b0000000000000011110001110;
    rom[4196] = 25'b0000000000000011110001110;
    rom[4197] = 25'b0000000000000011110001111;
    rom[4198] = 25'b0000000000000011110001111;
    rom[4199] = 25'b0000000000000011110001111;
    rom[4200] = 25'b0000000000000011110010000;
    rom[4201] = 25'b0000000000000011110010000;
    rom[4202] = 25'b0000000000000011110010000;
    rom[4203] = 25'b0000000000000011110010001;
    rom[4204] = 25'b0000000000000011110010001;
    rom[4205] = 25'b0000000000000011110010001;
    rom[4206] = 25'b0000000000000011110010001;
    rom[4207] = 25'b0000000000000011110010001;
    rom[4208] = 25'b0000000000000011110010001;
    rom[4209] = 25'b0000000000000011110010001;
    rom[4210] = 25'b0000000000000011110010010;
    rom[4211] = 25'b0000000000000011110010010;
    rom[4212] = 25'b0000000000000011110010010;
    rom[4213] = 25'b0000000000000011110010010;
    rom[4214] = 25'b0000000000000011110010011;
    rom[4215] = 25'b0000000000000011110010011;
    rom[4216] = 25'b0000000000000011110010011;
    rom[4217] = 25'b0000000000000011110010100;
    rom[4218] = 25'b0000000000000011110010100;
    rom[4219] = 25'b0000000000000011110010100;
    rom[4220] = 25'b0000000000000011110010100;
    rom[4221] = 25'b0000000000000011110010100;
    rom[4222] = 25'b0000000000000011110010100;
    rom[4223] = 25'b0000000000000011110010100;
    rom[4224] = 25'b0000000000000011110010100;
    rom[4225] = 25'b0000000000000011110010101;
    rom[4226] = 25'b0000000000000011110010101;
    rom[4227] = 25'b0000000000000011110010101;
    rom[4228] = 25'b0000000000000011110010101;
    rom[4229] = 25'b0000000000000011110010101;
    rom[4230] = 25'b0000000000000011110010110;
    rom[4231] = 25'b0000000000000011110010110;
    rom[4232] = 25'b0000000000000011110010110;
    rom[4233] = 25'b0000000000000011110010110;
    rom[4234] = 25'b0000000000000011110010111;
    rom[4235] = 25'b0000000000000011110010111;
    rom[4236] = 25'b0000000000000011110010111;
    rom[4237] = 25'b0000000000000011110010111;
    rom[4238] = 25'b0000000000000011110010111;
    rom[4239] = 25'b0000000000000011110010111;
    rom[4240] = 25'b0000000000000011110010111;
    rom[4241] = 25'b0000000000000011110010111;
    rom[4242] = 25'b0000000000000011110010111;
    rom[4243] = 25'b0000000000000011110010111;
    rom[4244] = 25'b0000000000000011110010111;
    rom[4245] = 25'b0000000000000011110010111;
    rom[4246] = 25'b0000000000000011110011000;
    rom[4247] = 25'b0000000000000011110011000;
    rom[4248] = 25'b0000000000000011110011000;
    rom[4249] = 25'b0000000000000011110011000;
    rom[4250] = 25'b0000000000000011110011000;
    rom[4251] = 25'b0000000000000011110011000;
    rom[4252] = 25'b0000000000000011110011001;
    rom[4253] = 25'b0000000000000011110011001;
    rom[4254] = 25'b0000000000000011110011001;
    rom[4255] = 25'b0000000000000011110011001;
    rom[4256] = 25'b0000000000000011110011001;
    rom[4257] = 25'b0000000000000011110011001;
    rom[4258] = 25'b0000000000000011110011001;
    rom[4259] = 25'b0000000000000011110011001;
    rom[4260] = 25'b0000000000000011110011001;
    rom[4261] = 25'b0000000000000011110011010;
    rom[4262] = 25'b0000000000000011110011010;
    rom[4263] = 25'b0000000000000011110011010;
    rom[4264] = 25'b0000000000000011110011010;
    rom[4265] = 25'b0000000000000011110011010;
    rom[4266] = 25'b0000000000000011110011010;
    rom[4267] = 25'b0000000000000011110011010;
    rom[4268] = 25'b0000000000000011110011010;
    rom[4269] = 25'b0000000000000011110011010;
    rom[4270] = 25'b0000000000000011110011010;
    rom[4271] = 25'b0000000000000011110011010;
    rom[4272] = 25'b0000000000000011110011010;
    rom[4273] = 25'b0000000000000011110011010;
    rom[4274] = 25'b0000000000000011110011010;
    rom[4275] = 25'b0000000000000011110011010;
    rom[4276] = 25'b0000000000000011110011010;
    rom[4277] = 25'b0000000000000011110011010;
    rom[4278] = 25'b0000000000000011110011010;
    rom[4279] = 25'b0000000000000011110011010;
    rom[4280] = 25'b0000000000000011110011010;
    rom[4281] = 25'b0000000000000011110011010;
    rom[4282] = 25'b0000000000000011110011010;
    rom[4283] = 25'b0000000000000011110011010;
    rom[4284] = 25'b0000000000000011110011010;
    rom[4285] = 25'b0000000000000011110011010;
    rom[4286] = 25'b0000000000000011110011010;
    rom[4287] = 25'b0000000000000011110011010;
    rom[4288] = 25'b0000000000000011110011010;
    rom[4289] = 25'b0000000000000011110011010;
    rom[4290] = 25'b0000000000000011110011010;
    rom[4291] = 25'b0000000000000011110011010;
    rom[4292] = 25'b0000000000000011110011010;
    rom[4293] = 25'b0000000000000011110011010;
    rom[4294] = 25'b0000000000000011110011010;
    rom[4295] = 25'b0000000000000011110011010;
    rom[4296] = 25'b0000000000000011110011010;
    rom[4297] = 25'b0000000000000011110011010;
    rom[4298] = 25'b0000000000000011110011010;
    rom[4299] = 25'b0000000000000011110011010;
    rom[4300] = 25'b0000000000000011110011010;
    rom[4301] = 25'b0000000000000011110011010;
    rom[4302] = 25'b0000000000000011110011010;
    rom[4303] = 25'b0000000000000011110011010;
    rom[4304] = 25'b0000000000000011110011010;
    rom[4305] = 25'b0000000000000011110011010;
    rom[4306] = 25'b0000000000000011110011010;
    rom[4307] = 25'b0000000000000011110011010;
    rom[4308] = 25'b0000000000000011110011010;
    rom[4309] = 25'b0000000000000011110011010;
    rom[4310] = 25'b0000000000000011110011010;
    rom[4311] = 25'b0000000000000011110011010;
    rom[4312] = 25'b0000000000000011110011001;
    rom[4313] = 25'b0000000000000011110011001;
    rom[4314] = 25'b0000000000000011110011001;
    rom[4315] = 25'b0000000000000011110011001;
    rom[4316] = 25'b0000000000000011110011001;
    rom[4317] = 25'b0000000000000011110011001;
    rom[4318] = 25'b0000000000000011110011001;
    rom[4319] = 25'b0000000000000011110011001;
    rom[4320] = 25'b0000000000000011110011001;
    rom[4321] = 25'b0000000000000011110011000;
    rom[4322] = 25'b0000000000000011110011000;
    rom[4323] = 25'b0000000000000011110011000;
    rom[4324] = 25'b0000000000000011110011000;
    rom[4325] = 25'b0000000000000011110011000;
    rom[4326] = 25'b0000000000000011110011000;
    rom[4327] = 25'b0000000000000011110010111;
    rom[4328] = 25'b0000000000000011110010111;
    rom[4329] = 25'b0000000000000011110010111;
    rom[4330] = 25'b0000000000000011110010111;
    rom[4331] = 25'b0000000000000011110010111;
    rom[4332] = 25'b0000000000000011110010111;
    rom[4333] = 25'b0000000000000011110010111;
    rom[4334] = 25'b0000000000000011110010111;
    rom[4335] = 25'b0000000000000011110010111;
    rom[4336] = 25'b0000000000000011110010111;
    rom[4337] = 25'b0000000000000011110010111;
    rom[4338] = 25'b0000000000000011110010110;
    rom[4339] = 25'b0000000000000011110010110;
    rom[4340] = 25'b0000000000000011110010110;
    rom[4341] = 25'b0000000000000011110010110;
    rom[4342] = 25'b0000000000000011110010110;
    rom[4343] = 25'b0000000000000011110010101;
    rom[4344] = 25'b0000000000000011110010101;
    rom[4345] = 25'b0000000000000011110010101;
    rom[4346] = 25'b0000000000000011110010101;
    rom[4347] = 25'b0000000000000011110010100;
    rom[4348] = 25'b0000000000000011110010100;
    rom[4349] = 25'b0000000000000011110010100;
    rom[4350] = 25'b0000000000000011110010100;
    rom[4351] = 25'b0000000000000011110010100;
    rom[4352] = 25'b0000000000000011110010100;
    rom[4353] = 25'b0000000000000011110010100;
    rom[4354] = 25'b0000000000000011110010100;
    rom[4355] = 25'b0000000000000011110010011;
    rom[4356] = 25'b0000000000000011110010011;
    rom[4357] = 25'b0000000000000011110010011;
    rom[4358] = 25'b0000000000000011110010010;
    rom[4359] = 25'b0000000000000011110010010;
    rom[4360] = 25'b0000000000000011110010010;
    rom[4361] = 25'b0000000000000011110010010;
    rom[4362] = 25'b0000000000000011110010001;
    rom[4363] = 25'b0000000000000011110010001;
    rom[4364] = 25'b0000000000000011110010001;
    rom[4365] = 25'b0000000000000011110010001;
    rom[4366] = 25'b0000000000000011110010001;
    rom[4367] = 25'b0000000000000011110010001;
    rom[4368] = 25'b0000000000000011110010000;
    rom[4369] = 25'b0000000000000011110010000;
    rom[4370] = 25'b0000000000000011110010000;
    rom[4371] = 25'b0000000000000011110001111;
    rom[4372] = 25'b0000000000000011110001111;
    rom[4373] = 25'b0000000000000011110001111;
    rom[4374] = 25'b0000000000000011110001110;
    rom[4375] = 25'b0000000000000011110001110;
    rom[4376] = 25'b0000000000000011110001110;
    rom[4377] = 25'b0000000000000011110001110;
    rom[4378] = 25'b0000000000000011110001110;
    rom[4379] = 25'b0000000000000011110001101;
    rom[4380] = 25'b0000000000000011110001101;
    rom[4381] = 25'b0000000000000011110001101;
    rom[4382] = 25'b0000000000000011110001100;
    rom[4383] = 25'b0000000000000011110001100;
    rom[4384] = 25'b0000000000000011110001100;
    rom[4385] = 25'b0000000000000011110001011;
    rom[4386] = 25'b0000000000000011110001011;
    rom[4387] = 25'b0000000000000011110001011;
    rom[4388] = 25'b0000000000000011110001011;
    rom[4389] = 25'b0000000000000011110001010;
    rom[4390] = 25'b0000000000000011110001010;
    rom[4391] = 25'b0000000000000011110001010;
    rom[4392] = 25'b0000000000000011110001001;
    rom[4393] = 25'b0000000000000011110001001;
    rom[4394] = 25'b0000000000000011110001001;
    rom[4395] = 25'b0000000000000011110001001;
    rom[4396] = 25'b0000000000000011110001000;
    rom[4397] = 25'b0000000000000011110001000;
    rom[4398] = 25'b0000000000000011110001000;
    rom[4399] = 25'b0000000000000011110000111;
    rom[4400] = 25'b0000000000000011110000111;
    rom[4401] = 25'b0000000000000011110000110;
    rom[4402] = 25'b0000000000000011110000110;
    rom[4403] = 25'b0000000000000011110000110;
    rom[4404] = 25'b0000000000000011110000110;
    rom[4405] = 25'b0000000000000011110000101;
    rom[4406] = 25'b0000000000000011110000101;
    rom[4407] = 25'b0000000000000011110000100;
    rom[4408] = 25'b0000000000000011110000100;
    rom[4409] = 25'b0000000000000011110000011;
    rom[4410] = 25'b0000000000000011110000011;
    rom[4411] = 25'b0000000000000011110000011;
    rom[4412] = 25'b0000000000000011110000011;
    rom[4413] = 25'b0000000000000011110000010;
    rom[4414] = 25'b0000000000000011110000010;
    rom[4415] = 25'b0000000000000011110000001;
    rom[4416] = 25'b0000000000000011110000001;
    rom[4417] = 25'b0000000000000011110000000;
    rom[4418] = 25'b0000000000000011110000000;
    rom[4419] = 25'b0000000000000011110000000;
    rom[4420] = 25'b0000000000000011101111111;
    rom[4421] = 25'b0000000000000011101111111;
    rom[4422] = 25'b0000000000000011101111110;
    rom[4423] = 25'b0000000000000011101111110;
    rom[4424] = 25'b0000000000000011101111101;
    rom[4425] = 25'b0000000000000011101111101;
    rom[4426] = 25'b0000000000000011101111101;
    rom[4427] = 25'b0000000000000011101111100;
    rom[4428] = 25'b0000000000000011101111100;
    rom[4429] = 25'b0000000000000011101111011;
    rom[4430] = 25'b0000000000000011101111011;
    rom[4431] = 25'b0000000000000011101111010;
    rom[4432] = 25'b0000000000000011101111010;
    rom[4433] = 25'b0000000000000011101111010;
    rom[4434] = 25'b0000000000000011101111001;
    rom[4435] = 25'b0000000000000011101111001;
    rom[4436] = 25'b0000000000000011101111000;
    rom[4437] = 25'b0000000000000011101110111;
    rom[4438] = 25'b0000000000000011101110111;
    rom[4439] = 25'b0000000000000011101110111;
    rom[4440] = 25'b0000000000000011101110111;
    rom[4441] = 25'b0000000000000011101110110;
    rom[4442] = 25'b0000000000000011101110101;
    rom[4443] = 25'b0000000000000011101110101;
    rom[4444] = 25'b0000000000000011101110100;
    rom[4445] = 25'b0000000000000011101110100;
    rom[4446] = 25'b0000000000000011101110100;
    rom[4447] = 25'b0000000000000011101110011;
    rom[4448] = 25'b0000000000000011101110010;
    rom[4449] = 25'b0000000000000011101110010;
    rom[4450] = 25'b0000000000000011101110001;
    rom[4451] = 25'b0000000000000011101110001;
    rom[4452] = 25'b0000000000000011101110001;
    rom[4453] = 25'b0000000000000011101110000;
    rom[4454] = 25'b0000000000000011101101111;
    rom[4455] = 25'b0000000000000011101101110;
    rom[4456] = 25'b0000000000000011101101110;
    rom[4457] = 25'b0000000000000011101101110;
    rom[4458] = 25'b0000000000000011101101101;
    rom[4459] = 25'b0000000000000011101101101;
    rom[4460] = 25'b0000000000000011101101100;
    rom[4461] = 25'b0000000000000011101101011;
    rom[4462] = 25'b0000000000000011101101011;
    rom[4463] = 25'b0000000000000011101101011;
    rom[4464] = 25'b0000000000000011101101010;
    rom[4465] = 25'b0000000000000011101101001;
    rom[4466] = 25'b0000000000000011101101000;
    rom[4467] = 25'b0000000000000011101101000;
    rom[4468] = 25'b0000000000000011101101000;
    rom[4469] = 25'b0000000000000011101100111;
    rom[4470] = 25'b0000000000000011101100110;
    rom[4471] = 25'b0000000000000011101100110;
    rom[4472] = 25'b0000000000000011101100101;
    rom[4473] = 25'b0000000000000011101100101;
    rom[4474] = 25'b0000000000000011101100100;
    rom[4475] = 25'b0000000000000011101100011;
    rom[4476] = 25'b0000000000000011101100011;
    rom[4477] = 25'b0000000000000011101100010;
    rom[4478] = 25'b0000000000000011101100010;
    rom[4479] = 25'b0000000000000011101100001;
    rom[4480] = 25'b0000000000000011101100000;
    rom[4481] = 25'b0000000000000011101100000;
    rom[4482] = 25'b0000000000000011101011111;
    rom[4483] = 25'b0000000000000011101011111;
    rom[4484] = 25'b0000000000000011101011110;
    rom[4485] = 25'b0000000000000011101011101;
    rom[4486] = 25'b0000000000000011101011100;
    rom[4487] = 25'b0000000000000011101011100;
    rom[4488] = 25'b0000000000000011101011100;
    rom[4489] = 25'b0000000000000011101011011;
    rom[4490] = 25'b0000000000000011101011010;
    rom[4491] = 25'b0000000000000011101011001;
    rom[4492] = 25'b0000000000000011101011001;
    rom[4493] = 25'b0000000000000011101011000;
    rom[4494] = 25'b0000000000000011101011000;
    rom[4495] = 25'b0000000000000011101010111;
    rom[4496] = 25'b0000000000000011101010110;
    rom[4497] = 25'b0000000000000011101010110;
    rom[4498] = 25'b0000000000000011101010101;
    rom[4499] = 25'b0000000000000011101010100;
    rom[4500] = 25'b0000000000000011101010011;
    rom[4501] = 25'b0000000000000011101010011;
    rom[4502] = 25'b0000000000000011101010010;
    rom[4503] = 25'b0000000000000011101010001;
    rom[4504] = 25'b0000000000000011101010001;
    rom[4505] = 25'b0000000000000011101010000;
    rom[4506] = 25'b0000000000000011101010000;
    rom[4507] = 25'b0000000000000011101001111;
    rom[4508] = 25'b0000000000000011101001110;
    rom[4509] = 25'b0000000000000011101001101;
    rom[4510] = 25'b0000000000000011101001101;
    rom[4511] = 25'b0000000000000011101001100;
    rom[4512] = 25'b0000000000000011101001011;
    rom[4513] = 25'b0000000000000011101001010;
    rom[4514] = 25'b0000000000000011101001010;
    rom[4515] = 25'b0000000000000011101001001;
    rom[4516] = 25'b0000000000000011101001000;
    rom[4517] = 25'b0000000000000011101001000;
    rom[4518] = 25'b0000000000000011101000111;
    rom[4519] = 25'b0000000000000011101000110;
    rom[4520] = 25'b0000000000000011101000101;
    rom[4521] = 25'b0000000000000011101000101;
    rom[4522] = 25'b0000000000000011101000100;
    rom[4523] = 25'b0000000000000011101000011;
    rom[4524] = 25'b0000000000000011101000010;
    rom[4525] = 25'b0000000000000011101000010;
    rom[4526] = 25'b0000000000000011101000001;
    rom[4527] = 25'b0000000000000011101000000;
    rom[4528] = 25'b0000000000000011100111111;
    rom[4529] = 25'b0000000000000011100111111;
    rom[4530] = 25'b0000000000000011100111110;
    rom[4531] = 25'b0000000000000011100111101;
    rom[4532] = 25'b0000000000000011100111100;
    rom[4533] = 25'b0000000000000011100111100;
    rom[4534] = 25'b0000000000000011100111011;
    rom[4535] = 25'b0000000000000011100111010;
    rom[4536] = 25'b0000000000000011100111001;
    rom[4537] = 25'b0000000000000011100111001;
    rom[4538] = 25'b0000000000000011100110111;
    rom[4539] = 25'b0000000000000011100110110;
    rom[4540] = 25'b0000000000000011100110110;
    rom[4541] = 25'b0000000000000011100110101;
    rom[4542] = 25'b0000000000000011100110100;
    rom[4543] = 25'b0000000000000011100110011;
    rom[4544] = 25'b0000000000000011100110011;
    rom[4545] = 25'b0000000000000011100110010;
    rom[4546] = 25'b0000000000000011100110001;
    rom[4547] = 25'b0000000000000011100110000;
    rom[4548] = 25'b0000000000000011100101111;
    rom[4549] = 25'b0000000000000011100101110;
    rom[4550] = 25'b0000000000000011100101101;
    rom[4551] = 25'b0000000000000011100101101;
    rom[4552] = 25'b0000000000000011100101100;
    rom[4553] = 25'b0000000000000011100101011;
    rom[4554] = 25'b0000000000000011100101010;
    rom[4555] = 25'b0000000000000011100101001;
    rom[4556] = 25'b0000000000000011100101000;
    rom[4557] = 25'b0000000000000011100100111;
    rom[4558] = 25'b0000000000000011100100111;
    rom[4559] = 25'b0000000000000011100100110;
    rom[4560] = 25'b0000000000000011100100101;
    rom[4561] = 25'b0000000000000011100100100;
    rom[4562] = 25'b0000000000000011100100011;
    rom[4563] = 25'b0000000000000011100100010;
    rom[4564] = 25'b0000000000000011100100001;
    rom[4565] = 25'b0000000000000011100100001;
    rom[4566] = 25'b0000000000000011100011111;
    rom[4567] = 25'b0000000000000011100011110;
    rom[4568] = 25'b0000000000000011100011110;
    rom[4569] = 25'b0000000000000011100011101;
    rom[4570] = 25'b0000000000000011100011100;
    rom[4571] = 25'b0000000000000011100011011;
    rom[4572] = 25'b0000000000000011100011010;
    rom[4573] = 25'b0000000000000011100011001;
    rom[4574] = 25'b0000000000000011100011000;
    rom[4575] = 25'b0000000000000011100010111;
    rom[4576] = 25'b0000000000000011100010110;
    rom[4577] = 25'b0000000000000011100010101;
    rom[4578] = 25'b0000000000000011100010101;
    rom[4579] = 25'b0000000000000011100010011;
    rom[4580] = 25'b0000000000000011100010010;
    rom[4581] = 25'b0000000000000011100010010;
    rom[4582] = 25'b0000000000000011100010000;
    rom[4583] = 25'b0000000000000011100001111;
    rom[4584] = 25'b0000000000000011100001111;
    rom[4585] = 25'b0000000000000011100001110;
    rom[4586] = 25'b0000000000000011100001100;
    rom[4587] = 25'b0000000000000011100001100;
    rom[4588] = 25'b0000000000000011100001011;
    rom[4589] = 25'b0000000000000011100001001;
    rom[4590] = 25'b0000000000000011100001001;
    rom[4591] = 25'b0000000000000011100001000;
    rom[4592] = 25'b0000000000000011100000111;
    rom[4593] = 25'b0000000000000011100000110;
    rom[4594] = 25'b0000000000000011100000101;
    rom[4595] = 25'b0000000000000011100000100;
    rom[4596] = 25'b0000000000000011100000011;
    rom[4597] = 25'b0000000000000011100000010;
    rom[4598] = 25'b0000000000000011100000001;
    rom[4599] = 25'b0000000000000011100000000;
    rom[4600] = 25'b0000000000000011011111111;
    rom[4601] = 25'b0000000000000011011111110;
    rom[4602] = 25'b0000000000000011011111101;
    rom[4603] = 25'b0000000000000011011111011;
    rom[4604] = 25'b0000000000000011011111011;
    rom[4605] = 25'b0000000000000011011111010;
    rom[4606] = 25'b0000000000000011011111000;
    rom[4607] = 25'b0000000000000011011111000;
    rom[4608] = 25'b0000000000000011011110110;
    rom[4609] = 25'b0000000000000011011110101;
    rom[4610] = 25'b0000000000000011011110101;
    rom[4611] = 25'b0000000000000011011110011;
    rom[4612] = 25'b0000000000000011011110010;
    rom[4613] = 25'b0000000000000011011110001;
    rom[4614] = 25'b0000000000000011011110000;
    rom[4615] = 25'b0000000000000011011101111;
    rom[4616] = 25'b0000000000000011011101110;
    rom[4617] = 25'b0000000000000011011101101;
    rom[4618] = 25'b0000000000000011011101100;
    rom[4619] = 25'b0000000000000011011101011;
    rom[4620] = 25'b0000000000000011011101001;
    rom[4621] = 25'b0000000000000011011101001;
    rom[4622] = 25'b0000000000000011011100111;
    rom[4623] = 25'b0000000000000011011100110;
    rom[4624] = 25'b0000000000000011011100101;
    rom[4625] = 25'b0000000000000011011100100;
    rom[4626] = 25'b0000000000000011011100011;
    rom[4627] = 25'b0000000000000011011100010;
    rom[4628] = 25'b0000000000000011011100000;
    rom[4629] = 25'b0000000000000011011100000;
    rom[4630] = 25'b0000000000000011011011110;
    rom[4631] = 25'b0000000000000011011011101;
    rom[4632] = 25'b0000000000000011011011100;
    rom[4633] = 25'b0000000000000011011011011;
    rom[4634] = 25'b0000000000000011011011010;
    rom[4635] = 25'b0000000000000011011011001;
    rom[4636] = 25'b0000000000000011011010111;
    rom[4637] = 25'b0000000000000011011010111;
    rom[4638] = 25'b0000000000000011011010101;
    rom[4639] = 25'b0000000000000011011010100;
    rom[4640] = 25'b0000000000000011011010011;
    rom[4641] = 25'b0000000000000011011010001;
    rom[4642] = 25'b0000000000000011011010001;
    rom[4643] = 25'b0000000000000011011001111;
    rom[4644] = 25'b0000000000000011011001110;
    rom[4645] = 25'b0000000000000011011001101;
    rom[4646] = 25'b0000000000000011011001100;
    rom[4647] = 25'b0000000000000011011001011;
    rom[4648] = 25'b0000000000000011011001001;
    rom[4649] = 25'b0000000000000011011001000;
    rom[4650] = 25'b0000000000000011011000111;
    rom[4651] = 25'b0000000000000011011000110;
    rom[4652] = 25'b0000000000000011011000101;
    rom[4653] = 25'b0000000000000011011000011;
    rom[4654] = 25'b0000000000000011011000011;
    rom[4655] = 25'b0000000000000011011000001;
    rom[4656] = 25'b0000000000000011011000000;
    rom[4657] = 25'b0000000000000011010111111;
    rom[4658] = 25'b0000000000000011010111101;
    rom[4659] = 25'b0000000000000011010111101;
    rom[4660] = 25'b0000000000000011010111011;
    rom[4661] = 25'b0000000000000011010111010;
    rom[4662] = 25'b0000000000000011010111001;
    rom[4663] = 25'b0000000000000011010110111;
    rom[4664] = 25'b0000000000000011010110110;
    rom[4665] = 25'b0000000000000011010110101;
    rom[4666] = 25'b0000000000000011010110100;
    rom[4667] = 25'b0000000000000011010110010;
    rom[4668] = 25'b0000000000000011010110001;
    rom[4669] = 25'b0000000000000011010110000;
    rom[4670] = 25'b0000000000000011010101110;
    rom[4671] = 25'b0000000000000011010101101;
    rom[4672] = 25'b0000000000000011010101100;
    rom[4673] = 25'b0000000000000011010101011;
    rom[4674] = 25'b0000000000000011010101001;
    rom[4675] = 25'b0000000000000011010101000;
    rom[4676] = 25'b0000000000000011010100111;
    rom[4677] = 25'b0000000000000011010100101;
    rom[4678] = 25'b0000000000000011010100100;
    rom[4679] = 25'b0000000000000011010100011;
    rom[4680] = 25'b0000000000000011010100010;
    rom[4681] = 25'b0000000000000011010100000;
    rom[4682] = 25'b0000000000000011010011111;
    rom[4683] = 25'b0000000000000011010011110;
    rom[4684] = 25'b0000000000000011010011100;
    rom[4685] = 25'b0000000000000011010011011;
    rom[4686] = 25'b0000000000000011010011001;
    rom[4687] = 25'b0000000000000011010011000;
    rom[4688] = 25'b0000000000000011010010111;
    rom[4689] = 25'b0000000000000011010010110;
    rom[4690] = 25'b0000000000000011010010100;
    rom[4691] = 25'b0000000000000011010010011;
    rom[4692] = 25'b0000000000000011010010001;
    rom[4693] = 25'b0000000000000011010010000;
    rom[4694] = 25'b0000000000000011010001111;
    rom[4695] = 25'b0000000000000011010001101;
    rom[4696] = 25'b0000000000000011010001100;
    rom[4697] = 25'b0000000000000011010001010;
    rom[4698] = 25'b0000000000000011010001010;
    rom[4699] = 25'b0000000000000011010001000;
    rom[4700] = 25'b0000000000000011010000111;
    rom[4701] = 25'b0000000000000011010000101;
    rom[4702] = 25'b0000000000000011010000100;
    rom[4703] = 25'b0000000000000011010000010;
    rom[4704] = 25'b0000000000000011010000001;
    rom[4705] = 25'b0000000000000011010000000;
    rom[4706] = 25'b0000000000000011001111111;
    rom[4707] = 25'b0000000000000011001111101;
    rom[4708] = 25'b0000000000000011001111100;
    rom[4709] = 25'b0000000000000011001111010;
    rom[4710] = 25'b0000000000000011001111001;
    rom[4711] = 25'b0000000000000011001110111;
    rom[4712] = 25'b0000000000000011001110110;
    rom[4713] = 25'b0000000000000011001110100;
    rom[4714] = 25'b0000000000000011001110011;
    rom[4715] = 25'b0000000000000011001110010;
    rom[4716] = 25'b0000000000000011001110000;
    rom[4717] = 25'b0000000000000011001101111;
    rom[4718] = 25'b0000000000000011001101101;
    rom[4719] = 25'b0000000000000011001101100;
    rom[4720] = 25'b0000000000000011001101010;
    rom[4721] = 25'b0000000000000011001101001;
    rom[4722] = 25'b0000000000000011001100111;
    rom[4723] = 25'b0000000000000011001100110;
    rom[4724] = 25'b0000000000000011001100100;
    rom[4725] = 25'b0000000000000011001100011;
    rom[4726] = 25'b0000000000000011001100001;
    rom[4727] = 25'b0000000000000011001100000;
    rom[4728] = 25'b0000000000000011001011110;
    rom[4729] = 25'b0000000000000011001011101;
    rom[4730] = 25'b0000000000000011001011011;
    rom[4731] = 25'b0000000000000011001011010;
    rom[4732] = 25'b0000000000000011001011000;
    rom[4733] = 25'b0000000000000011001010111;
    rom[4734] = 25'b0000000000000011001010101;
    rom[4735] = 25'b0000000000000011001010100;
    rom[4736] = 25'b0000000000000011001010010;
    rom[4737] = 25'b0000000000000011001010001;
    rom[4738] = 25'b0000000000000011001001111;
    rom[4739] = 25'b0000000000000011001001110;
    rom[4740] = 25'b0000000000000011001001100;
    rom[4741] = 25'b0000000000000011001001011;
    rom[4742] = 25'b0000000000000011001001001;
    rom[4743] = 25'b0000000000000011001001000;
    rom[4744] = 25'b0000000000000011001000111;
    rom[4745] = 25'b0000000000000011001000101;
    rom[4746] = 25'b0000000000000011001000100;
    rom[4747] = 25'b0000000000000011001000010;
    rom[4748] = 25'b0000000000000011001000000;
    rom[4749] = 25'b0000000000000011000111110;
    rom[4750] = 25'b0000000000000011000111101;
    rom[4751] = 25'b0000000000000011000111011;
    rom[4752] = 25'b0000000000000011000111010;
    rom[4753] = 25'b0000000000000011000111000;
    rom[4754] = 25'b0000000000000011000110111;
    rom[4755] = 25'b0000000000000011000110101;
    rom[4756] = 25'b0000000000000011000110100;
    rom[4757] = 25'b0000000000000011000110010;
    rom[4758] = 25'b0000000000000011000110000;
    rom[4759] = 25'b0000000000000011000101111;
    rom[4760] = 25'b0000000000000011000101101;
    rom[4761] = 25'b0000000000000011000101100;
    rom[4762] = 25'b0000000000000011000101010;
    rom[4763] = 25'b0000000000000011000101001;
    rom[4764] = 25'b0000000000000011000100111;
    rom[4765] = 25'b0000000000000011000100101;
    rom[4766] = 25'b0000000000000011000100011;
    rom[4767] = 25'b0000000000000011000100010;
    rom[4768] = 25'b0000000000000011000100000;
    rom[4769] = 25'b0000000000000011000011111;
    rom[4770] = 25'b0000000000000011000011101;
    rom[4771] = 25'b0000000000000011000011011;
    rom[4772] = 25'b0000000000000011000011010;
    rom[4773] = 25'b0000000000000011000011000;
    rom[4774] = 25'b0000000000000011000010111;
    rom[4775] = 25'b0000000000000011000010100;
    rom[4776] = 25'b0000000000000011000010011;
    rom[4777] = 25'b0000000000000011000010001;
    rom[4778] = 25'b0000000000000011000010000;
    rom[4779] = 25'b0000000000000011000001110;
    rom[4780] = 25'b0000000000000011000001100;
    rom[4781] = 25'b0000000000000011000001011;
    rom[4782] = 25'b0000000000000011000001001;
    rom[4783] = 25'b0000000000000011000001000;
    rom[4784] = 25'b0000000000000011000000110;
    rom[4785] = 25'b0000000000000011000000100;
    rom[4786] = 25'b0000000000000011000000011;
    rom[4787] = 25'b0000000000000011000000001;
    rom[4788] = 25'b0000000000000010111111111;
    rom[4789] = 25'b0000000000000010111111101;
    rom[4790] = 25'b0000000000000010111111100;
    rom[4791] = 25'b0000000000000010111111010;
    rom[4792] = 25'b0000000000000010111111000;
    rom[4793] = 25'b0000000000000010111110111;
    rom[4794] = 25'b0000000000000010111110100;
    rom[4795] = 25'b0000000000000010111110011;
    rom[4796] = 25'b0000000000000010111110001;
    rom[4797] = 25'b0000000000000010111110000;
    rom[4798] = 25'b0000000000000010111101110;
    rom[4799] = 25'b0000000000000010111101100;
    rom[4800] = 25'b0000000000000010111101011;
    rom[4801] = 25'b0000000000000010111101000;
    rom[4802] = 25'b0000000000000010111100111;
    rom[4803] = 25'b0000000000000010111100101;
    rom[4804] = 25'b0000000000000010111100011;
    rom[4805] = 25'b0000000000000010111100010;
    rom[4806] = 25'b0000000000000010111011111;
    rom[4807] = 25'b0000000000000010111011110;
    rom[4808] = 25'b0000000000000010111011100;
    rom[4809] = 25'b0000000000000010111011010;
    rom[4810] = 25'b0000000000000010111011001;
    rom[4811] = 25'b0000000000000010111010111;
    rom[4812] = 25'b0000000000000010111010101;
    rom[4813] = 25'b0000000000000010111010011;
    rom[4814] = 25'b0000000000000010111010001;
    rom[4815] = 25'b0000000000000010111010000;
    rom[4816] = 25'b0000000000000010111001101;
    rom[4817] = 25'b0000000000000010111001100;
    rom[4818] = 25'b0000000000000010111001010;
    rom[4819] = 25'b0000000000000010111001000;
    rom[4820] = 25'b0000000000000010111000111;
    rom[4821] = 25'b0000000000000010111000101;
    rom[4822] = 25'b0000000000000010111000011;
    rom[4823] = 25'b0000000000000010111000001;
    rom[4824] = 25'b0000000000000010110111111;
    rom[4825] = 25'b0000000000000010110111110;
    rom[4826] = 25'b0000000000000010110111100;
    rom[4827] = 25'b0000000000000010110111010;
    rom[4828] = 25'b0000000000000010110111000;
    rom[4829] = 25'b0000000000000010110110110;
    rom[4830] = 25'b0000000000000010110110100;
    rom[4831] = 25'b0000000000000010110110011;
    rom[4832] = 25'b0000000000000010110110000;
    rom[4833] = 25'b0000000000000010110101111;
    rom[4834] = 25'b0000000000000010110101101;
    rom[4835] = 25'b0000000000000010110101011;
    rom[4836] = 25'b0000000000000010110101001;
    rom[4837] = 25'b0000000000000010110100111;
    rom[4838] = 25'b0000000000000010110100101;
    rom[4839] = 25'b0000000000000010110100100;
    rom[4840] = 25'b0000000000000010110100001;
    rom[4841] = 25'b0000000000000010110011111;
    rom[4842] = 25'b0000000000000010110011110;
    rom[4843] = 25'b0000000000000010110011011;
    rom[4844] = 25'b0000000000000010110011010;
    rom[4845] = 25'b0000000000000010110011000;
    rom[4846] = 25'b0000000000000010110010110;
    rom[4847] = 25'b0000000000000010110010100;
    rom[4848] = 25'b0000000000000010110010010;
    rom[4849] = 25'b0000000000000010110010000;
    rom[4850] = 25'b0000000000000010110001110;
    rom[4851] = 25'b0000000000000010110001100;
    rom[4852] = 25'b0000000000000010110001010;
    rom[4853] = 25'b0000000000000010110001001;
    rom[4854] = 25'b0000000000000010110000111;
    rom[4855] = 25'b0000000000000010110000100;
    rom[4856] = 25'b0000000000000010110000011;
    rom[4857] = 25'b0000000000000010110000001;
    rom[4858] = 25'b0000000000000010101111111;
    rom[4859] = 25'b0000000000000010101111101;
    rom[4860] = 25'b0000000000000010101111011;
    rom[4861] = 25'b0000000000000010101111001;
    rom[4862] = 25'b0000000000000010101110111;
    rom[4863] = 25'b0000000000000010101110101;
    rom[4864] = 25'b0000000000000010101110011;
    rom[4865] = 25'b0000000000000010101110001;
    rom[4866] = 25'b0000000000000010101101111;
    rom[4867] = 25'b0000000000000010101101101;
    rom[4868] = 25'b0000000000000010101101011;
    rom[4869] = 25'b0000000000000010101101001;
    rom[4870] = 25'b0000000000000010101100111;
    rom[4871] = 25'b0000000000000010101100101;
    rom[4872] = 25'b0000000000000010101100011;
    rom[4873] = 25'b0000000000000010101100001;
    rom[4874] = 25'b0000000000000010101011111;
    rom[4875] = 25'b0000000000000010101011101;
    rom[4876] = 25'b0000000000000010101011011;
    rom[4877] = 25'b0000000000000010101011001;
    rom[4878] = 25'b0000000000000010101010111;
    rom[4879] = 25'b0000000000000010101010100;
    rom[4880] = 25'b0000000000000010101010011;
    rom[4881] = 25'b0000000000000010101010001;
    rom[4882] = 25'b0000000000000010101001110;
    rom[4883] = 25'b0000000000000010101001100;
    rom[4884] = 25'b0000000000000010101001011;
    rom[4885] = 25'b0000000000000010101001000;
    rom[4886] = 25'b0000000000000010101000110;
    rom[4887] = 25'b0000000000000010101000100;
    rom[4888] = 25'b0000000000000010101000011;
    rom[4889] = 25'b0000000000000010101000000;
    rom[4890] = 25'b0000000000000010100111110;
    rom[4891] = 25'b0000000000000010100111100;
    rom[4892] = 25'b0000000000000010100111010;
    rom[4893] = 25'b0000000000000010100111000;
    rom[4894] = 25'b0000000000000010100110110;
    rom[4895] = 25'b0000000000000010100110100;
    rom[4896] = 25'b0000000000000010100110001;
    rom[4897] = 25'b0000000000000010100101111;
    rom[4898] = 25'b0000000000000010100101110;
    rom[4899] = 25'b0000000000000010100101011;
    rom[4900] = 25'b0000000000000010100101001;
    rom[4901] = 25'b0000000000000010100100111;
    rom[4902] = 25'b0000000000000010100100101;
    rom[4903] = 25'b0000000000000010100100010;
    rom[4904] = 25'b0000000000000010100100001;
    rom[4905] = 25'b0000000000000010100011111;
    rom[4906] = 25'b0000000000000010100011100;
    rom[4907] = 25'b0000000000000010100011010;
    rom[4908] = 25'b0000000000000010100011000;
    rom[4909] = 25'b0000000000000010100010110;
    rom[4910] = 25'b0000000000000010100010011;
    rom[4911] = 25'b0000000000000010100010010;
    rom[4912] = 25'b0000000000000010100010000;
    rom[4913] = 25'b0000000000000010100001101;
    rom[4914] = 25'b0000000000000010100001011;
    rom[4915] = 25'b0000000000000010100001001;
    rom[4916] = 25'b0000000000000010100000111;
    rom[4917] = 25'b0000000000000010100000101;
    rom[4918] = 25'b0000000000000010100000010;
    rom[4919] = 25'b0000000000000010100000000;
    rom[4920] = 25'b0000000000000010011111110;
    rom[4921] = 25'b0000000000000010011111100;
    rom[4922] = 25'b0000000000000010011111001;
    rom[4923] = 25'b0000000000000010011111000;
    rom[4924] = 25'b0000000000000010011110110;
    rom[4925] = 25'b0000000000000010011110011;
    rom[4926] = 25'b0000000000000010011110001;
    rom[4927] = 25'b0000000000000010011101111;
    rom[4928] = 25'b0000000000000010011101101;
    rom[4929] = 25'b0000000000000010011101010;
    rom[4930] = 25'b0000000000000010011101000;
    rom[4931] = 25'b0000000000000010011100110;
    rom[4932] = 25'b0000000000000010011100100;
    rom[4933] = 25'b0000000000000010011100001;
    rom[4934] = 25'b0000000000000010011011111;
    rom[4935] = 25'b0000000000000010011011101;
    rom[4936] = 25'b0000000000000010011011011;
    rom[4937] = 25'b0000000000000010011011000;
    rom[4938] = 25'b0000000000000010011010110;
    rom[4939] = 25'b0000000000000010011010100;
    rom[4940] = 25'b0000000000000010011010010;
    rom[4941] = 25'b0000000000000010011001111;
    rom[4942] = 25'b0000000000000010011001101;
    rom[4943] = 25'b0000000000000010011001011;
    rom[4944] = 25'b0000000000000010011001001;
    rom[4945] = 25'b0000000000000010011000110;
    rom[4946] = 25'b0000000000000010011000100;
    rom[4947] = 25'b0000000000000010011000001;
    rom[4948] = 25'b0000000000000010010111111;
    rom[4949] = 25'b0000000000000010010111101;
    rom[4950] = 25'b0000000000000010010111011;
    rom[4951] = 25'b0000000000000010010111000;
    rom[4952] = 25'b0000000000000010010110110;
    rom[4953] = 25'b0000000000000010010110100;
    rom[4954] = 25'b0000000000000010010110010;
    rom[4955] = 25'b0000000000000010010101111;
    rom[4956] = 25'b0000000000000010010101101;
    rom[4957] = 25'b0000000000000010010101010;
    rom[4958] = 25'b0000000000000010010101000;
    rom[4959] = 25'b0000000000000010010100110;
    rom[4960] = 25'b0000000000000010010100011;
    rom[4961] = 25'b0000000000000010010100001;
    rom[4962] = 25'b0000000000000010010011111;
    rom[4963] = 25'b0000000000000010010011101;
    rom[4964] = 25'b0000000000000010010011010;
    rom[4965] = 25'b0000000000000010010010111;
    rom[4966] = 25'b0000000000000010010010101;
    rom[4967] = 25'b0000000000000010010010011;
    rom[4968] = 25'b0000000000000010010010001;
    rom[4969] = 25'b0000000000000010010001110;
    rom[4970] = 25'b0000000000000010010001100;
    rom[4971] = 25'b0000000000000010010001001;
    rom[4972] = 25'b0000000000000010010000111;
    rom[4973] = 25'b0000000000000010010000101;
    rom[4974] = 25'b0000000000000010010000011;
    rom[4975] = 25'b0000000000000010010000000;
    rom[4976] = 25'b0000000000000010001111101;
    rom[4977] = 25'b0000000000000010001111011;
    rom[4978] = 25'b0000000000000010001111001;
    rom[4979] = 25'b0000000000000010001110111;
    rom[4980] = 25'b0000000000000010001110100;
    rom[4981] = 25'b0000000000000010001110001;
    rom[4982] = 25'b0000000000000010001101111;
    rom[4983] = 25'b0000000000000010001101101;
    rom[4984] = 25'b0000000000000010001101011;
    rom[4985] = 25'b0000000000000010001101000;
    rom[4986] = 25'b0000000000000010001100101;
    rom[4987] = 25'b0000000000000010001100011;
    rom[4988] = 25'b0000000000000010001100001;
    rom[4989] = 25'b0000000000000010001011110;
    rom[4990] = 25'b0000000000000010001011100;
    rom[4991] = 25'b0000000000000010001011001;
    rom[4992] = 25'b0000000000000010001010111;
    rom[4993] = 25'b0000000000000010001010100;
    rom[4994] = 25'b0000000000000010001010010;
    rom[4995] = 25'b0000000000000010001010000;
    rom[4996] = 25'b0000000000000010001001101;
    rom[4997] = 25'b0000000000000010001001010;
    rom[4998] = 25'b0000000000000010001001000;
    rom[4999] = 25'b0000000000000010001000101;
    rom[5000] = 25'b0000000000000010001000011;
    rom[5001] = 25'b0000000000000010001000001;
    rom[5002] = 25'b0000000000000010000111110;
    rom[5003] = 25'b0000000000000010000111100;
    rom[5004] = 25'b0000000000000010000111001;
    rom[5005] = 25'b0000000000000010000110110;
    rom[5006] = 25'b0000000000000010000110100;
    rom[5007] = 25'b0000000000000010000110010;
    rom[5008] = 25'b0000000000000010000101111;
    rom[5009] = 25'b0000000000000010000101101;
    rom[5010] = 25'b0000000000000010000101010;
    rom[5011] = 25'b0000000000000010000100111;
    rom[5012] = 25'b0000000000000010000100101;
    rom[5013] = 25'b0000000000000010000100011;
    rom[5014] = 25'b0000000000000010000100000;
    rom[5015] = 25'b0000000000000010000011110;
    rom[5016] = 25'b0000000000000010000011011;
    rom[5017] = 25'b0000000000000010000011000;
    rom[5018] = 25'b0000000000000010000010110;
    rom[5019] = 25'b0000000000000010000010011;
    rom[5020] = 25'b0000000000000010000010001;
    rom[5021] = 25'b0000000000000010000001110;
    rom[5022] = 25'b0000000000000010000001100;
    rom[5023] = 25'b0000000000000010000001001;
    rom[5024] = 25'b0000000000000010000000110;
    rom[5025] = 25'b0000000000000010000000100;
    rom[5026] = 25'b0000000000000010000000001;
    rom[5027] = 25'b0000000000000001111111111;
    rom[5028] = 25'b0000000000000001111111100;
    rom[5029] = 25'b0000000000000001111111010;
    rom[5030] = 25'b0000000000000001111110111;
    rom[5031] = 25'b0000000000000001111110101;
    rom[5032] = 25'b0000000000000001111110010;
    rom[5033] = 25'b0000000000000001111101111;
    rom[5034] = 25'b0000000000000001111101100;
    rom[5035] = 25'b0000000000000001111101010;
    rom[5036] = 25'b0000000000000001111100111;
    rom[5037] = 25'b0000000000000001111100101;
    rom[5038] = 25'b0000000000000001111100010;
    rom[5039] = 25'b0000000000000001111100000;
    rom[5040] = 25'b0000000000000001111011101;
    rom[5041] = 25'b0000000000000001111011010;
    rom[5042] = 25'b0000000000000001111010111;
    rom[5043] = 25'b0000000000000001111010101;
    rom[5044] = 25'b0000000000000001111010010;
    rom[5045] = 25'b0000000000000001111010000;
    rom[5046] = 25'b0000000000000001111001101;
    rom[5047] = 25'b0000000000000001111001011;
    rom[5048] = 25'b0000000000000001111001000;
    rom[5049] = 25'b0000000000000001111000101;
    rom[5050] = 25'b0000000000000001111000011;
    rom[5051] = 25'b0000000000000001111000000;
    rom[5052] = 25'b0000000000000001110111101;
    rom[5053] = 25'b0000000000000001110111010;
    rom[5054] = 25'b0000000000000001110111000;
    rom[5055] = 25'b0000000000000001110110101;
    rom[5056] = 25'b0000000000000001110110010;
    rom[5057] = 25'b0000000000000001110110000;
    rom[5058] = 25'b0000000000000001110101101;
    rom[5059] = 25'b0000000000000001110101011;
    rom[5060] = 25'b0000000000000001110101000;
    rom[5061] = 25'b0000000000000001110100101;
    rom[5062] = 25'b0000000000000001110100010;
    rom[5063] = 25'b0000000000000001110011111;
    rom[5064] = 25'b0000000000000001110011101;
    rom[5065] = 25'b0000000000000001110011010;
    rom[5066] = 25'b0000000000000001110010111;
    rom[5067] = 25'b0000000000000001110010101;
    rom[5068] = 25'b0000000000000001110010010;
    rom[5069] = 25'b0000000000000001110001111;
    rom[5070] = 25'b0000000000000001110001101;
    rom[5071] = 25'b0000000000000001110001010;
    rom[5072] = 25'b0000000000000001110000111;
    rom[5073] = 25'b0000000000000001110000100;
    rom[5074] = 25'b0000000000000001110000010;
    rom[5075] = 25'b0000000000000001101111111;
    rom[5076] = 25'b0000000000000001101111100;
    rom[5077] = 25'b0000000000000001101111001;
    rom[5078] = 25'b0000000000000001101110110;
    rom[5079] = 25'b0000000000000001101110100;
    rom[5080] = 25'b0000000000000001101110001;
    rom[5081] = 25'b0000000000000001101101110;
    rom[5082] = 25'b0000000000000001101101011;
    rom[5083] = 25'b0000000000000001101101001;
    rom[5084] = 25'b0000000000000001101100110;
    rom[5085] = 25'b0000000000000001101100011;
    rom[5086] = 25'b0000000000000001101100001;
    rom[5087] = 25'b0000000000000001101011110;
    rom[5088] = 25'b0000000000000001101011011;
    rom[5089] = 25'b0000000000000001101011000;
    rom[5090] = 25'b0000000000000001101010101;
    rom[5091] = 25'b0000000000000001101010010;
    rom[5092] = 25'b0000000000000001101001111;
    rom[5093] = 25'b0000000000000001101001100;
    rom[5094] = 25'b0000000000000001101001010;
    rom[5095] = 25'b0000000000000001101000111;
    rom[5096] = 25'b0000000000000001101000100;
    rom[5097] = 25'b0000000000000001101000001;
    rom[5098] = 25'b0000000000000001100111110;
    rom[5099] = 25'b0000000000000001100111100;
    rom[5100] = 25'b0000000000000001100111001;
    rom[5101] = 25'b0000000000000001100110110;
    rom[5102] = 25'b0000000000000001100110011;
    rom[5103] = 25'b0000000000000001100110000;
    rom[5104] = 25'b0000000000000001100101110;
    rom[5105] = 25'b0000000000000001100101011;
    rom[5106] = 25'b0000000000000001100101000;
    rom[5107] = 25'b0000000000000001100100101;
    rom[5108] = 25'b0000000000000001100100010;
    rom[5109] = 25'b0000000000000001100011111;
    rom[5110] = 25'b0000000000000001100011101;
    rom[5111] = 25'b0000000000000001100011010;
    rom[5112] = 25'b0000000000000001100010111;
    rom[5113] = 25'b0000000000000001100010100;
    rom[5114] = 25'b0000000000000001100010001;
    rom[5115] = 25'b0000000000000001100001110;
    rom[5116] = 25'b0000000000000001100001011;
    rom[5117] = 25'b0000000000000001100001000;
    rom[5118] = 25'b0000000000000001100000101;
    rom[5119] = 25'b0000000000000001100000011;
    rom[5120] = 25'b0000000000000001100000000;
    rom[5121] = 25'b0000000000000001011111101;
    rom[5122] = 25'b0000000000000001011111010;
    rom[5123] = 25'b0000000000000001011110111;
    rom[5124] = 25'b0000000000000001011110100;
    rom[5125] = 25'b0000000000000001011110001;
    rom[5126] = 25'b0000000000000001011101110;
    rom[5127] = 25'b0000000000000001011101011;
    rom[5128] = 25'b0000000000000001011101000;
    rom[5129] = 25'b0000000000000001011100101;
    rom[5130] = 25'b0000000000000001011100010;
    rom[5131] = 25'b0000000000000001011011111;
    rom[5132] = 25'b0000000000000001011011100;
    rom[5133] = 25'b0000000000000001011011001;
    rom[5134] = 25'b0000000000000001011010110;
    rom[5135] = 25'b0000000000000001011010011;
    rom[5136] = 25'b0000000000000001011010000;
    rom[5137] = 25'b0000000000000001011001101;
    rom[5138] = 25'b0000000000000001011001010;
    rom[5139] = 25'b0000000000000001011000111;
    rom[5140] = 25'b0000000000000001011000100;
    rom[5141] = 25'b0000000000000001011000010;
    rom[5142] = 25'b0000000000000001010111111;
    rom[5143] = 25'b0000000000000001010111100;
    rom[5144] = 25'b0000000000000001010111001;
    rom[5145] = 25'b0000000000000001010110110;
    rom[5146] = 25'b0000000000000001010110011;
    rom[5147] = 25'b0000000000000001010110000;
    rom[5148] = 25'b0000000000000001010101101;
    rom[5149] = 25'b0000000000000001010101010;
    rom[5150] = 25'b0000000000000001010100111;
    rom[5151] = 25'b0000000000000001010100100;
    rom[5152] = 25'b0000000000000001010100001;
    rom[5153] = 25'b0000000000000001010011110;
    rom[5154] = 25'b0000000000000001010011011;
    rom[5155] = 25'b0000000000000001010011000;
    rom[5156] = 25'b0000000000000001010010101;
    rom[5157] = 25'b0000000000000001010010010;
    rom[5158] = 25'b0000000000000001010001111;
    rom[5159] = 25'b0000000000000001010001011;
    rom[5160] = 25'b0000000000000001010001000;
    rom[5161] = 25'b0000000000000001010000101;
    rom[5162] = 25'b0000000000000001010000010;
    rom[5163] = 25'b0000000000000001001111111;
    rom[5164] = 25'b0000000000000001001111100;
    rom[5165] = 25'b0000000000000001001111001;
    rom[5166] = 25'b0000000000000001001110110;
    rom[5167] = 25'b0000000000000001001110011;
    rom[5168] = 25'b0000000000000001001110000;
    rom[5169] = 25'b0000000000000001001101101;
    rom[5170] = 25'b0000000000000001001101001;
    rom[5171] = 25'b0000000000000001001100110;
    rom[5172] = 25'b0000000000000001001100011;
    rom[5173] = 25'b0000000000000001001100000;
    rom[5174] = 25'b0000000000000001001011101;
    rom[5175] = 25'b0000000000000001001011010;
    rom[5176] = 25'b0000000000000001001010111;
    rom[5177] = 25'b0000000000000001001010100;
    rom[5178] = 25'b0000000000000001001010001;
    rom[5179] = 25'b0000000000000001001001110;
    rom[5180] = 25'b0000000000000001001001011;
    rom[5181] = 25'b0000000000000001001001000;
    rom[5182] = 25'b0000000000000001001000101;
    rom[5183] = 25'b0000000000000001001000001;
    rom[5184] = 25'b0000000000000001000111110;
    rom[5185] = 25'b0000000000000001000111011;
    rom[5186] = 25'b0000000000000001000111000;
    rom[5187] = 25'b0000000000000001000110101;
    rom[5188] = 25'b0000000000000001000110001;
    rom[5189] = 25'b0000000000000001000101110;
    rom[5190] = 25'b0000000000000001000101011;
    rom[5191] = 25'b0000000000000001000101000;
    rom[5192] = 25'b0000000000000001000100101;
    rom[5193] = 25'b0000000000000001000100010;
    rom[5194] = 25'b0000000000000001000011111;
    rom[5195] = 25'b0000000000000001000011100;
    rom[5196] = 25'b0000000000000001000011001;
    rom[5197] = 25'b0000000000000001000010101;
    rom[5198] = 25'b0000000000000001000010010;
    rom[5199] = 25'b0000000000000001000001111;
    rom[5200] = 25'b0000000000000001000001100;
    rom[5201] = 25'b0000000000000001000001000;
    rom[5202] = 25'b0000000000000001000000101;
    rom[5203] = 25'b0000000000000001000000010;
    rom[5204] = 25'b0000000000000000111111111;
    rom[5205] = 25'b0000000000000000111111100;
    rom[5206] = 25'b0000000000000000111111001;
    rom[5207] = 25'b0000000000000000111110110;
    rom[5208] = 25'b0000000000000000111110010;
    rom[5209] = 25'b0000000000000000111101111;
    rom[5210] = 25'b0000000000000000111101100;
    rom[5211] = 25'b0000000000000000111101001;
    rom[5212] = 25'b0000000000000000111100101;
    rom[5213] = 25'b0000000000000000111100010;
    rom[5214] = 25'b0000000000000000111011111;
    rom[5215] = 25'b0000000000000000111011011;
    rom[5216] = 25'b0000000000000000111011000;
    rom[5217] = 25'b0000000000000000111010101;
    rom[5218] = 25'b0000000000000000111010010;
    rom[5219] = 25'b0000000000000000111001111;
    rom[5220] = 25'b0000000000000000111001100;
    rom[5221] = 25'b0000000000000000111001000;
    rom[5222] = 25'b0000000000000000111000101;
    rom[5223] = 25'b0000000000000000111000010;
    rom[5224] = 25'b0000000000000000110111110;
    rom[5225] = 25'b0000000000000000110111011;
    rom[5226] = 25'b0000000000000000110111000;
    rom[5227] = 25'b0000000000000000110110101;
    rom[5228] = 25'b0000000000000000110110010;
    rom[5229] = 25'b0000000000000000110101110;
    rom[5230] = 25'b0000000000000000110101011;
    rom[5231] = 25'b0000000000000000110101000;
    rom[5232] = 25'b0000000000000000110100100;
    rom[5233] = 25'b0000000000000000110100001;
    rom[5234] = 25'b0000000000000000110011101;
    rom[5235] = 25'b0000000000000000110011010;
    rom[5236] = 25'b0000000000000000110010111;
    rom[5237] = 25'b0000000000000000110010100;
    rom[5238] = 25'b0000000000000000110010001;
    rom[5239] = 25'b0000000000000000110001101;
    rom[5240] = 25'b0000000000000000110001010;
    rom[5241] = 25'b0000000000000000110000110;
    rom[5242] = 25'b0000000000000000110000011;
    rom[5243] = 25'b0000000000000000110000000;
    rom[5244] = 25'b0000000000000000101111101;
    rom[5245] = 25'b0000000000000000101111010;
    rom[5246] = 25'b0000000000000000101110110;
    rom[5247] = 25'b0000000000000000101110011;
    rom[5248] = 25'b0000000000000000101101111;
    rom[5249] = 25'b0000000000000000101101100;
    rom[5250] = 25'b0000000000000000101101000;
    rom[5251] = 25'b0000000000000000101100101;
    rom[5252] = 25'b0000000000000000101100010;
    rom[5253] = 25'b0000000000000000101011111;
    rom[5254] = 25'b0000000000000000101011011;
    rom[5255] = 25'b0000000000000000101011000;
    rom[5256] = 25'b0000000000000000101010100;
    rom[5257] = 25'b0000000000000000101010001;
    rom[5258] = 25'b0000000000000000101001101;
    rom[5259] = 25'b0000000000000000101001010;
    rom[5260] = 25'b0000000000000000101000111;
    rom[5261] = 25'b0000000000000000101000100;
    rom[5262] = 25'b0000000000000000101000000;
    rom[5263] = 25'b0000000000000000100111101;
    rom[5264] = 25'b0000000000000000100111001;
    rom[5265] = 25'b0000000000000000100110110;
    rom[5266] = 25'b0000000000000000100110011;
    rom[5267] = 25'b0000000000000000100110000;
    rom[5268] = 25'b0000000000000000100101100;
    rom[5269] = 25'b0000000000000000100101000;
    rom[5270] = 25'b0000000000000000100100101;
    rom[5271] = 25'b0000000000000000100100001;
    rom[5272] = 25'b0000000000000000100011110;
    rom[5273] = 25'b0000000000000000100011011;
    rom[5274] = 25'b0000000000000000100011000;
    rom[5275] = 25'b0000000000000000100010100;
    rom[5276] = 25'b0000000000000000100010000;
    rom[5277] = 25'b0000000000000000100001101;
    rom[5278] = 25'b0000000000000000100001001;
    rom[5279] = 25'b0000000000000000100000110;
    rom[5280] = 25'b0000000000000000100000011;
    rom[5281] = 25'b0000000000000000100000000;
    rom[5282] = 25'b0000000000000000011111100;
    rom[5283] = 25'b0000000000000000011111000;
    rom[5284] = 25'b0000000000000000011110101;
    rom[5285] = 25'b0000000000000000011110010;
    rom[5286] = 25'b0000000000000000011101110;
    rom[5287] = 25'b0000000000000000011101011;
    rom[5288] = 25'b0000000000000000011100111;
    rom[5289] = 25'b0000000000000000011100100;
    rom[5290] = 25'b0000000000000000011100000;
    rom[5291] = 25'b0000000000000000011011101;
    rom[5292] = 25'b0000000000000000011011010;
    rom[5293] = 25'b0000000000000000011010110;
    rom[5294] = 25'b0000000000000000011010010;
    rom[5295] = 25'b0000000000000000011001111;
    rom[5296] = 25'b0000000000000000011001011;
    rom[5297] = 25'b0000000000000000011001000;
    rom[5298] = 25'b0000000000000000011000101;
    rom[5299] = 25'b0000000000000000011000001;
    rom[5300] = 25'b0000000000000000010111101;
    rom[5301] = 25'b0000000000000000010111010;
    rom[5302] = 25'b0000000000000000010110111;
    rom[5303] = 25'b0000000000000000010110011;
    rom[5304] = 25'b0000000000000000010101111;
    rom[5305] = 25'b0000000000000000010101100;
    rom[5306] = 25'b0000000000000000010101000;
    rom[5307] = 25'b0000000000000000010100101;
    rom[5308] = 25'b0000000000000000010100010;
    rom[5309] = 25'b0000000000000000010011110;
    rom[5310] = 25'b0000000000000000010011010;
    rom[5311] = 25'b0000000000000000010010110;
    rom[5312] = 25'b0000000000000000010010011;
    rom[5313] = 25'b0000000000000000010010000;
    rom[5314] = 25'b0000000000000000010001100;
    rom[5315] = 25'b0000000000000000010001000;
    rom[5316] = 25'b0000000000000000010000101;
    rom[5317] = 25'b0000000000000000010000001;
    rom[5318] = 25'b0000000000000000001111110;
    rom[5319] = 25'b0000000000000000001111010;
    rom[5320] = 25'b0000000000000000001110111;
    rom[5321] = 25'b0000000000000000001110011;
    rom[5322] = 25'b0000000000000000001110000;
    rom[5323] = 25'b0000000000000000001101100;
    rom[5324] = 25'b0000000000000000001101001;
    rom[5325] = 25'b0000000000000000001100101;
    rom[5326] = 25'b0000000000000000001100001;
    rom[5327] = 25'b0000000000000000001011110;
    rom[5328] = 25'b0000000000000000001011010;
    rom[5329] = 25'b0000000000000000001010111;
    rom[5330] = 25'b0000000000000000001010011;
    rom[5331] = 25'b0000000000000000001001111;
    rom[5332] = 25'b0000000000000000001001100;
    rom[5333] = 25'b0000000000000000001001000;
    rom[5334] = 25'b0000000000000000001000101;
    rom[5335] = 25'b0000000000000000001000001;
    rom[5336] = 25'b0000000000000000000111110;
    rom[5337] = 25'b0000000000000000000111010;
    rom[5338] = 25'b0000000000000000000110110;
    rom[5339] = 25'b0000000000000000000110010;
    rom[5340] = 25'b0000000000000000000101111;
    rom[5341] = 25'b0000000000000000000101100;
    rom[5342] = 25'b0000000000000000000101000;
    rom[5343] = 25'b0000000000000000000100100;
    rom[5344] = 25'b0000000000000000000100000;
    rom[5345] = 25'b0000000000000000000011101;
    rom[5346] = 25'b0000000000000000000011001;
    rom[5347] = 25'b0000000000000000000010110;
    rom[5348] = 25'b0000000000000000000010010;
    rom[5349] = 25'b0000000000000000000001110;
    rom[5350] = 25'b0000000000000000000001011;
    rom[5351] = 25'b0000000000000000000000111;
    rom[5352] = 25'b0000000000000000000000011;
    rom[5353] = 25'b0000000000000000000000000;
    rom[5354] = 25'b1111111111111111111111101;
    rom[5355] = 25'b1111111111111111111111001;
    rom[5356] = 25'b1111111111111111111110110;
    rom[5357] = 25'b1111111111111111111110010;
    rom[5358] = 25'b1111111111111111111101110;
    rom[5359] = 25'b1111111111111111111101011;
    rom[5360] = 25'b1111111111111111111100111;
    rom[5361] = 25'b1111111111111111111100011;
    rom[5362] = 25'b1111111111111111111011111;
    rom[5363] = 25'b1111111111111111111011100;
    rom[5364] = 25'b1111111111111111111011000;
    rom[5365] = 25'b1111111111111111111010100;
    rom[5366] = 25'b1111111111111111111010000;
    rom[5367] = 25'b1111111111111111111001101;
    rom[5368] = 25'b1111111111111111111001001;
    rom[5369] = 25'b1111111111111111111000101;
    rom[5370] = 25'b1111111111111111111000001;
    rom[5371] = 25'b1111111111111111110111110;
    rom[5372] = 25'b1111111111111111110111011;
    rom[5373] = 25'b1111111111111111110110111;
    rom[5374] = 25'b1111111111111111110110011;
    rom[5375] = 25'b1111111111111111110110000;
    rom[5376] = 25'b1111111111111111110101100;
    rom[5377] = 25'b1111111111111111110101000;
    rom[5378] = 25'b1111111111111111110100100;
    rom[5379] = 25'b1111111111111111110100001;
    rom[5380] = 25'b1111111111111111110011101;
    rom[5381] = 25'b1111111111111111110011001;
    rom[5382] = 25'b1111111111111111110010101;
    rom[5383] = 25'b1111111111111111110010010;
    rom[5384] = 25'b1111111111111111110001110;
    rom[5385] = 25'b1111111111111111110001010;
    rom[5386] = 25'b1111111111111111110000110;
    rom[5387] = 25'b1111111111111111110000011;
    rom[5388] = 25'b1111111111111111101111111;
    rom[5389] = 25'b1111111111111111101111011;
    rom[5390] = 25'b1111111111111111101110111;
    rom[5391] = 25'b1111111111111111101110011;
    rom[5392] = 25'b1111111111111111101101111;
    rom[5393] = 25'b1111111111111111101101100;
    rom[5394] = 25'b1111111111111111101101000;
    rom[5395] = 25'b1111111111111111101100100;
    rom[5396] = 25'b1111111111111111101100000;
    rom[5397] = 25'b1111111111111111101011101;
    rom[5398] = 25'b1111111111111111101011001;
    rom[5399] = 25'b1111111111111111101010101;
    rom[5400] = 25'b1111111111111111101010001;
    rom[5401] = 25'b1111111111111111101001110;
    rom[5402] = 25'b1111111111111111101001010;
    rom[5403] = 25'b1111111111111111101000110;
    rom[5404] = 25'b1111111111111111101000010;
    rom[5405] = 25'b1111111111111111100111110;
    rom[5406] = 25'b1111111111111111100111010;
    rom[5407] = 25'b1111111111111111100110111;
    rom[5408] = 25'b1111111111111111100110011;
    rom[5409] = 25'b1111111111111111100101111;
    rom[5410] = 25'b1111111111111111100101011;
    rom[5411] = 25'b1111111111111111100101000;
    rom[5412] = 25'b1111111111111111100100100;
    rom[5413] = 25'b1111111111111111100100000;
    rom[5414] = 25'b1111111111111111100011100;
    rom[5415] = 25'b1111111111111111100011000;
    rom[5416] = 25'b1111111111111111100010100;
    rom[5417] = 25'b1111111111111111100010000;
    rom[5418] = 25'b1111111111111111100001101;
    rom[5419] = 25'b1111111111111111100001001;
    rom[5420] = 25'b1111111111111111100000101;
    rom[5421] = 25'b1111111111111111100000001;
    rom[5422] = 25'b1111111111111111011111101;
    rom[5423] = 25'b1111111111111111011111001;
    rom[5424] = 25'b1111111111111111011110110;
    rom[5425] = 25'b1111111111111111011110010;
    rom[5426] = 25'b1111111111111111011101110;
    rom[5427] = 25'b1111111111111111011101010;
    rom[5428] = 25'b1111111111111111011100110;
    rom[5429] = 25'b1111111111111111011100010;
    rom[5430] = 25'b1111111111111111011011110;
    rom[5431] = 25'b1111111111111111011011011;
    rom[5432] = 25'b1111111111111111011010111;
    rom[5433] = 25'b1111111111111111011010010;
    rom[5434] = 25'b1111111111111111011001111;
    rom[5435] = 25'b1111111111111111011001011;
    rom[5436] = 25'b1111111111111111011000111;
    rom[5437] = 25'b1111111111111111011000011;
    rom[5438] = 25'b1111111111111111010111111;
    rom[5439] = 25'b1111111111111111010111011;
    rom[5440] = 25'b1111111111111111010111000;
    rom[5441] = 25'b1111111111111111010110100;
    rom[5442] = 25'b1111111111111111010110000;
    rom[5443] = 25'b1111111111111111010101100;
    rom[5444] = 25'b1111111111111111010101000;
    rom[5445] = 25'b1111111111111111010100100;
    rom[5446] = 25'b1111111111111111010100000;
    rom[5447] = 25'b1111111111111111010011100;
    rom[5448] = 25'b1111111111111111010011000;
    rom[5449] = 25'b1111111111111111010010100;
    rom[5450] = 25'b1111111111111111010010001;
    rom[5451] = 25'b1111111111111111010001100;
    rom[5452] = 25'b1111111111111111010001000;
    rom[5453] = 25'b1111111111111111010000101;
    rom[5454] = 25'b1111111111111111010000001;
    rom[5455] = 25'b1111111111111111001111101;
    rom[5456] = 25'b1111111111111111001111001;
    rom[5457] = 25'b1111111111111111001110101;
    rom[5458] = 25'b1111111111111111001110001;
    rom[5459] = 25'b1111111111111111001101101;
    rom[5460] = 25'b1111111111111111001101001;
    rom[5461] = 25'b1111111111111111001100101;
    rom[5462] = 25'b1111111111111111001100001;
    rom[5463] = 25'b1111111111111111001011101;
    rom[5464] = 25'b1111111111111111001011001;
    rom[5465] = 25'b1111111111111111001010110;
    rom[5466] = 25'b1111111111111111001010001;
    rom[5467] = 25'b1111111111111111001001101;
    rom[5468] = 25'b1111111111111111001001010;
    rom[5469] = 25'b1111111111111111001000101;
    rom[5470] = 25'b1111111111111111001000001;
    rom[5471] = 25'b1111111111111111000111110;
    rom[5472] = 25'b1111111111111111000111001;
    rom[5473] = 25'b1111111111111111000110110;
    rom[5474] = 25'b1111111111111111000110010;
    rom[5475] = 25'b1111111111111111000101101;
    rom[5476] = 25'b1111111111111111000101010;
    rom[5477] = 25'b1111111111111111000100110;
    rom[5478] = 25'b1111111111111111000100001;
    rom[5479] = 25'b1111111111111111000011110;
    rom[5480] = 25'b1111111111111111000011010;
    rom[5481] = 25'b1111111111111111000010101;
    rom[5482] = 25'b1111111111111111000010010;
    rom[5483] = 25'b1111111111111111000001110;
    rom[5484] = 25'b1111111111111111000001001;
    rom[5485] = 25'b1111111111111111000000110;
    rom[5486] = 25'b1111111111111111000000010;
    rom[5487] = 25'b1111111111111110111111101;
    rom[5488] = 25'b1111111111111110111111010;
    rom[5489] = 25'b1111111111111110111110101;
    rom[5490] = 25'b1111111111111110111110010;
    rom[5491] = 25'b1111111111111110111101110;
    rom[5492] = 25'b1111111111111110111101001;
    rom[5493] = 25'b1111111111111110111100110;
    rom[5494] = 25'b1111111111111110111100001;
    rom[5495] = 25'b1111111111111110111011101;
    rom[5496] = 25'b1111111111111110111011010;
    rom[5497] = 25'b1111111111111110111010101;
    rom[5498] = 25'b1111111111111110111010001;
    rom[5499] = 25'b1111111111111110111001101;
    rom[5500] = 25'b1111111111111110111001001;
    rom[5501] = 25'b1111111111111110111000101;
    rom[5502] = 25'b1111111111111110111000001;
    rom[5503] = 25'b1111111111111110110111101;
    rom[5504] = 25'b1111111111111110110111001;
    rom[5505] = 25'b1111111111111110110110101;
    rom[5506] = 25'b1111111111111110110110001;
    rom[5507] = 25'b1111111111111110110101101;
    rom[5508] = 25'b1111111111111110110101001;
    rom[5509] = 25'b1111111111111110110100101;
    rom[5510] = 25'b1111111111111110110100001;
    rom[5511] = 25'b1111111111111110110011100;
    rom[5512] = 25'b1111111111111110110011001;
    rom[5513] = 25'b1111111111111110110010100;
    rom[5514] = 25'b1111111111111110110010000;
    rom[5515] = 25'b1111111111111110110001100;
    rom[5516] = 25'b1111111111111110110001000;
    rom[5517] = 25'b1111111111111110110000100;
    rom[5518] = 25'b1111111111111110110000000;
    rom[5519] = 25'b1111111111111110101111100;
    rom[5520] = 25'b1111111111111110101111000;
    rom[5521] = 25'b1111111111111110101110100;
    rom[5522] = 25'b1111111111111110101110000;
    rom[5523] = 25'b1111111111111110101101100;
    rom[5524] = 25'b1111111111111110101100111;
    rom[5525] = 25'b1111111111111110101100100;
    rom[5526] = 25'b1111111111111110101011111;
    rom[5527] = 25'b1111111111111110101011011;
    rom[5528] = 25'b1111111111111110101010111;
    rom[5529] = 25'b1111111111111110101010011;
    rom[5530] = 25'b1111111111111110101001111;
    rom[5531] = 25'b1111111111111110101001011;
    rom[5532] = 25'b1111111111111110101000110;
    rom[5533] = 25'b1111111111111110101000011;
    rom[5534] = 25'b1111111111111110100111110;
    rom[5535] = 25'b1111111111111110100111011;
    rom[5536] = 25'b1111111111111110100110110;
    rom[5537] = 25'b1111111111111110100110010;
    rom[5538] = 25'b1111111111111110100101110;
    rom[5539] = 25'b1111111111111110100101010;
    rom[5540] = 25'b1111111111111110100100110;
    rom[5541] = 25'b1111111111111110100100001;
    rom[5542] = 25'b1111111111111110100011101;
    rom[5543] = 25'b1111111111111110100011001;
    rom[5544] = 25'b1111111111111110100010101;
    rom[5545] = 25'b1111111111111110100010001;
    rom[5546] = 25'b1111111111111110100001101;
    rom[5547] = 25'b1111111111111110100001000;
    rom[5548] = 25'b1111111111111110100000101;
    rom[5549] = 25'b1111111111111110100000000;
    rom[5550] = 25'b1111111111111110011111100;
    rom[5551] = 25'b1111111111111110011111000;
    rom[5552] = 25'b1111111111111110011110100;
    rom[5553] = 25'b1111111111111110011110000;
    rom[5554] = 25'b1111111111111110011101011;
    rom[5555] = 25'b1111111111111110011101000;
    rom[5556] = 25'b1111111111111110011100011;
    rom[5557] = 25'b1111111111111110011011111;
    rom[5558] = 25'b1111111111111110011011011;
    rom[5559] = 25'b1111111111111110011010110;
    rom[5560] = 25'b1111111111111110011010011;
    rom[5561] = 25'b1111111111111110011001110;
    rom[5562] = 25'b1111111111111110011001010;
    rom[5563] = 25'b1111111111111110011000110;
    rom[5564] = 25'b1111111111111110011000001;
    rom[5565] = 25'b1111111111111110010111110;
    rom[5566] = 25'b1111111111111110010111001;
    rom[5567] = 25'b1111111111111110010110101;
    rom[5568] = 25'b1111111111111110010110001;
    rom[5569] = 25'b1111111111111110010101101;
    rom[5570] = 25'b1111111111111110010101001;
    rom[5571] = 25'b1111111111111110010100100;
    rom[5572] = 25'b1111111111111110010100000;
    rom[5573] = 25'b1111111111111110010011100;
    rom[5574] = 25'b1111111111111110010011000;
    rom[5575] = 25'b1111111111111110010010100;
    rom[5576] = 25'b1111111111111110010001111;
    rom[5577] = 25'b1111111111111110010001011;
    rom[5578] = 25'b1111111111111110010000111;
    rom[5579] = 25'b1111111111111110010000011;
    rom[5580] = 25'b1111111111111110001111110;
    rom[5581] = 25'b1111111111111110001111011;
    rom[5582] = 25'b1111111111111110001110110;
    rom[5583] = 25'b1111111111111110001110010;
    rom[5584] = 25'b1111111111111110001101110;
    rom[5585] = 25'b1111111111111110001101001;
    rom[5586] = 25'b1111111111111110001100101;
    rom[5587] = 25'b1111111111111110001100001;
    rom[5588] = 25'b1111111111111110001011101;
    rom[5589] = 25'b1111111111111110001011000;
    rom[5590] = 25'b1111111111111110001010100;
    rom[5591] = 25'b1111111111111110001010000;
    rom[5592] = 25'b1111111111111110001001011;
    rom[5593] = 25'b1111111111111110001001000;
    rom[5594] = 25'b1111111111111110001000011;
    rom[5595] = 25'b1111111111111110000111111;
    rom[5596] = 25'b1111111111111110000111011;
    rom[5597] = 25'b1111111111111110000110111;
    rom[5598] = 25'b1111111111111110000110010;
    rom[5599] = 25'b1111111111111110000101110;
    rom[5600] = 25'b1111111111111110000101010;
    rom[5601] = 25'b1111111111111110000100101;
    rom[5602] = 25'b1111111111111110000100001;
    rom[5603] = 25'b1111111111111110000011101;
    rom[5604] = 25'b1111111111111110000011001;
    rom[5605] = 25'b1111111111111110000010100;
    rom[5606] = 25'b1111111111111110000010000;
    rom[5607] = 25'b1111111111111110000001100;
    rom[5608] = 25'b1111111111111110000000111;
    rom[5609] = 25'b1111111111111110000000011;
    rom[5610] = 25'b1111111111111101111111111;
    rom[5611] = 25'b1111111111111101111111011;
    rom[5612] = 25'b1111111111111101111110110;
    rom[5613] = 25'b1111111111111101111110011;
    rom[5614] = 25'b1111111111111101111101110;
    rom[5615] = 25'b1111111111111101111101010;
    rom[5616] = 25'b1111111111111101111100101;
    rom[5617] = 25'b1111111111111101111100001;
    rom[5618] = 25'b1111111111111101111011101;
    rom[5619] = 25'b1111111111111101111011000;
    rom[5620] = 25'b1111111111111101111010100;
    rom[5621] = 25'b1111111111111101111010000;
    rom[5622] = 25'b1111111111111101111001100;
    rom[5623] = 25'b1111111111111101111000111;
    rom[5624] = 25'b1111111111111101111000011;
    rom[5625] = 25'b1111111111111101110111111;
    rom[5626] = 25'b1111111111111101110111010;
    rom[5627] = 25'b1111111111111101110110110;
    rom[5628] = 25'b1111111111111101110110010;
    rom[5629] = 25'b1111111111111101110101110;
    rom[5630] = 25'b1111111111111101110101001;
    rom[5631] = 25'b1111111111111101110100101;
    rom[5632] = 25'b1111111111111101110100000;
    rom[5633] = 25'b1111111111111101110011101;
    rom[5634] = 25'b1111111111111101110011000;
    rom[5635] = 25'b1111111111111101110010100;
    rom[5636] = 25'b1111111111111101110001111;
    rom[5637] = 25'b1111111111111101110001011;
    rom[5638] = 25'b1111111111111101110000111;
    rom[5639] = 25'b1111111111111101110000010;
    rom[5640] = 25'b1111111111111101101111110;
    rom[5641] = 25'b1111111111111101101111010;
    rom[5642] = 25'b1111111111111101101110101;
    rom[5643] = 25'b1111111111111101101110001;
    rom[5644] = 25'b1111111111111101101101101;
    rom[5645] = 25'b1111111111111101101101000;
    rom[5646] = 25'b1111111111111101101100100;
    rom[5647] = 25'b1111111111111101101011111;
    rom[5648] = 25'b1111111111111101101011100;
    rom[5649] = 25'b1111111111111101101010111;
    rom[5650] = 25'b1111111111111101101010011;
    rom[5651] = 25'b1111111111111101101001110;
    rom[5652] = 25'b1111111111111101101001010;
    rom[5653] = 25'b1111111111111101101000110;
    rom[5654] = 25'b1111111111111101101000001;
    rom[5655] = 25'b1111111111111101100111101;
    rom[5656] = 25'b1111111111111101100111001;
    rom[5657] = 25'b1111111111111101100110100;
    rom[5658] = 25'b1111111111111101100110000;
    rom[5659] = 25'b1111111111111101100101100;
    rom[5660] = 25'b1111111111111101100100111;
    rom[5661] = 25'b1111111111111101100100011;
    rom[5662] = 25'b1111111111111101100011110;
    rom[5663] = 25'b1111111111111101100011010;
    rom[5664] = 25'b1111111111111101100010101;
    rom[5665] = 25'b1111111111111101100010010;
    rom[5666] = 25'b1111111111111101100001101;
    rom[5667] = 25'b1111111111111101100001001;
    rom[5668] = 25'b1111111111111101100000100;
    rom[5669] = 25'b1111111111111101100000000;
    rom[5670] = 25'b1111111111111101011111011;
    rom[5671] = 25'b1111111111111101011110111;
    rom[5672] = 25'b1111111111111101011110011;
    rom[5673] = 25'b1111111111111101011101111;
    rom[5674] = 25'b1111111111111101011101010;
    rom[5675] = 25'b1111111111111101011100110;
    rom[5676] = 25'b1111111111111101011100001;
    rom[5677] = 25'b1111111111111101011011101;
    rom[5678] = 25'b1111111111111101011011000;
    rom[5679] = 25'b1111111111111101011010100;
    rom[5680] = 25'b1111111111111101011010000;
    rom[5681] = 25'b1111111111111101011001011;
    rom[5682] = 25'b1111111111111101011000111;
    rom[5683] = 25'b1111111111111101011000010;
    rom[5684] = 25'b1111111111111101010111110;
    rom[5685] = 25'b1111111111111101010111001;
    rom[5686] = 25'b1111111111111101010110101;
    rom[5687] = 25'b1111111111111101010110001;
    rom[5688] = 25'b1111111111111101010101100;
    rom[5689] = 25'b1111111111111101010101000;
    rom[5690] = 25'b1111111111111101010100100;
    rom[5691] = 25'b1111111111111101010011111;
    rom[5692] = 25'b1111111111111101010011011;
    rom[5693] = 25'b1111111111111101010010110;
    rom[5694] = 25'b1111111111111101010010010;
    rom[5695] = 25'b1111111111111101010001101;
    rom[5696] = 25'b1111111111111101010001001;
    rom[5697] = 25'b1111111111111101010000100;
    rom[5698] = 25'b1111111111111101010000000;
    rom[5699] = 25'b1111111111111101001111100;
    rom[5700] = 25'b1111111111111101001111000;
    rom[5701] = 25'b1111111111111101001110011;
    rom[5702] = 25'b1111111111111101001101111;
    rom[5703] = 25'b1111111111111101001101010;
    rom[5704] = 25'b1111111111111101001100110;
    rom[5705] = 25'b1111111111111101001100001;
    rom[5706] = 25'b1111111111111101001011101;
    rom[5707] = 25'b1111111111111101001011000;
    rom[5708] = 25'b1111111111111101001010100;
    rom[5709] = 25'b1111111111111101001001111;
    rom[5710] = 25'b1111111111111101001001011;
    rom[5711] = 25'b1111111111111101001000110;
    rom[5712] = 25'b1111111111111101001000011;
    rom[5713] = 25'b1111111111111101000111110;
    rom[5714] = 25'b1111111111111101000111010;
    rom[5715] = 25'b1111111111111101000110101;
    rom[5716] = 25'b1111111111111101000110001;
    rom[5717] = 25'b1111111111111101000101100;
    rom[5718] = 25'b1111111111111101000101000;
    rom[5719] = 25'b1111111111111101000100011;
    rom[5720] = 25'b1111111111111101000011111;
    rom[5721] = 25'b1111111111111101000011010;
    rom[5722] = 25'b1111111111111101000010110;
    rom[5723] = 25'b1111111111111101000010001;
    rom[5724] = 25'b1111111111111101000001101;
    rom[5725] = 25'b1111111111111101000001000;
    rom[5726] = 25'b1111111111111101000000100;
    rom[5727] = 25'b1111111111111100111111111;
    rom[5728] = 25'b1111111111111100111111011;
    rom[5729] = 25'b1111111111111100111110111;
    rom[5730] = 25'b1111111111111100111110010;
    rom[5731] = 25'b1111111111111100111101110;
    rom[5732] = 25'b1111111111111100111101001;
    rom[5733] = 25'b1111111111111100111100101;
    rom[5734] = 25'b1111111111111100111100001;
    rom[5735] = 25'b1111111111111100111011100;
    rom[5736] = 25'b1111111111111100111011000;
    rom[5737] = 25'b1111111111111100111010011;
    rom[5738] = 25'b1111111111111100111001111;
    rom[5739] = 25'b1111111111111100111001010;
    rom[5740] = 25'b1111111111111100111000110;
    rom[5741] = 25'b1111111111111100111000001;
    rom[5742] = 25'b1111111111111100110111101;
    rom[5743] = 25'b1111111111111100110111000;
    rom[5744] = 25'b1111111111111100110110100;
    rom[5745] = 25'b1111111111111100110110000;
    rom[5746] = 25'b1111111111111100110101011;
    rom[5747] = 25'b1111111111111100110100111;
    rom[5748] = 25'b1111111111111100110100010;
    rom[5749] = 25'b1111111111111100110011110;
    rom[5750] = 25'b1111111111111100110011001;
    rom[5751] = 25'b1111111111111100110010101;
    rom[5752] = 25'b1111111111111100110010000;
    rom[5753] = 25'b1111111111111100110001100;
    rom[5754] = 25'b1111111111111100110000111;
    rom[5755] = 25'b1111111111111100110000011;
    rom[5756] = 25'b1111111111111100101111110;
    rom[5757] = 25'b1111111111111100101111010;
    rom[5758] = 25'b1111111111111100101110101;
    rom[5759] = 25'b1111111111111100101110001;
    rom[5760] = 25'b1111111111111100101101100;
    rom[5761] = 25'b1111111111111100101101000;
    rom[5762] = 25'b1111111111111100101100011;
    rom[5763] = 25'b1111111111111100101011111;
    rom[5764] = 25'b1111111111111100101011010;
    rom[5765] = 25'b1111111111111100101010110;
    rom[5766] = 25'b1111111111111100101010001;
    rom[5767] = 25'b1111111111111100101001101;
    rom[5768] = 25'b1111111111111100101001000;
    rom[5769] = 25'b1111111111111100101000100;
    rom[5770] = 25'b1111111111111100100111111;
    rom[5771] = 25'b1111111111111100100111011;
    rom[5772] = 25'b1111111111111100100110111;
    rom[5773] = 25'b1111111111111100100110010;
    rom[5774] = 25'b1111111111111100100101110;
    rom[5775] = 25'b1111111111111100100101000;
    rom[5776] = 25'b1111111111111100100100100;
    rom[5777] = 25'b1111111111111100100011111;
    rom[5778] = 25'b1111111111111100100011011;
    rom[5779] = 25'b1111111111111100100010110;
    rom[5780] = 25'b1111111111111100100010010;
    rom[5781] = 25'b1111111111111100100001101;
    rom[5782] = 25'b1111111111111100100001001;
    rom[5783] = 25'b1111111111111100100000100;
    rom[5784] = 25'b1111111111111100100000000;
    rom[5785] = 25'b1111111111111100011111011;
    rom[5786] = 25'b1111111111111100011110111;
    rom[5787] = 25'b1111111111111100011110011;
    rom[5788] = 25'b1111111111111100011101110;
    rom[5789] = 25'b1111111111111100011101010;
    rom[5790] = 25'b1111111111111100011100101;
    rom[5791] = 25'b1111111111111100011100001;
    rom[5792] = 25'b1111111111111100011011100;
    rom[5793] = 25'b1111111111111100011011000;
    rom[5794] = 25'b1111111111111100011010011;
    rom[5795] = 25'b1111111111111100011001111;
    rom[5796] = 25'b1111111111111100011001010;
    rom[5797] = 25'b1111111111111100011000110;
    rom[5798] = 25'b1111111111111100011000001;
    rom[5799] = 25'b1111111111111100010111100;
    rom[5800] = 25'b1111111111111100010110111;
    rom[5801] = 25'b1111111111111100010110011;
    rom[5802] = 25'b1111111111111100010101111;
    rom[5803] = 25'b1111111111111100010101010;
    rom[5804] = 25'b1111111111111100010100110;
    rom[5805] = 25'b1111111111111100010100001;
    rom[5806] = 25'b1111111111111100010011101;
    rom[5807] = 25'b1111111111111100010011000;
    rom[5808] = 25'b1111111111111100010010100;
    rom[5809] = 25'b1111111111111100010001111;
    rom[5810] = 25'b1111111111111100010001011;
    rom[5811] = 25'b1111111111111100010000110;
    rom[5812] = 25'b1111111111111100010000010;
    rom[5813] = 25'b1111111111111100001111101;
    rom[5814] = 25'b1111111111111100001111001;
    rom[5815] = 25'b1111111111111100001110100;
    rom[5816] = 25'b1111111111111100001101111;
    rom[5817] = 25'b1111111111111100001101011;
    rom[5818] = 25'b1111111111111100001100110;
    rom[5819] = 25'b1111111111111100001100010;
    rom[5820] = 25'b1111111111111100001011101;
    rom[5821] = 25'b1111111111111100001011001;
    rom[5822] = 25'b1111111111111100001010100;
    rom[5823] = 25'b1111111111111100001010000;
    rom[5824] = 25'b1111111111111100001001011;
    rom[5825] = 25'b1111111111111100001000111;
    rom[5826] = 25'b1111111111111100001000010;
    rom[5827] = 25'b1111111111111100000111110;
    rom[5828] = 25'b1111111111111100000111000;
    rom[5829] = 25'b1111111111111100000110100;
    rom[5830] = 25'b1111111111111100000110000;
    rom[5831] = 25'b1111111111111100000101011;
    rom[5832] = 25'b1111111111111100000100111;
    rom[5833] = 25'b1111111111111100000100010;
    rom[5834] = 25'b1111111111111100000011110;
    rom[5835] = 25'b1111111111111100000011001;
    rom[5836] = 25'b1111111111111100000010101;
    rom[5837] = 25'b1111111111111100000010000;
    rom[5838] = 25'b1111111111111100000001100;
    rom[5839] = 25'b1111111111111100000000111;
    rom[5840] = 25'b1111111111111100000000010;
    rom[5841] = 25'b1111111111111011111111101;
    rom[5842] = 25'b1111111111111011111111001;
    rom[5843] = 25'b1111111111111011111110101;
    rom[5844] = 25'b1111111111111011111110000;
    rom[5845] = 25'b1111111111111011111101100;
    rom[5846] = 25'b1111111111111011111100111;
    rom[5847] = 25'b1111111111111011111100011;
    rom[5848] = 25'b1111111111111011111011110;
    rom[5849] = 25'b1111111111111011111011010;
    rom[5850] = 25'b1111111111111011111010100;
    rom[5851] = 25'b1111111111111011111010000;
    rom[5852] = 25'b1111111111111011111001011;
    rom[5853] = 25'b1111111111111011111000111;
    rom[5854] = 25'b1111111111111011111000010;
    rom[5855] = 25'b1111111111111011110111110;
    rom[5856] = 25'b1111111111111011110111001;
    rom[5857] = 25'b1111111111111011110110101;
    rom[5858] = 25'b1111111111111011110110001;
    rom[5859] = 25'b1111111111111011110101100;
    rom[5860] = 25'b1111111111111011110100111;
    rom[5861] = 25'b1111111111111011110100010;
    rom[5862] = 25'b1111111111111011110011110;
    rom[5863] = 25'b1111111111111011110011001;
    rom[5864] = 25'b1111111111111011110010101;
    rom[5865] = 25'b1111111111111011110010000;
    rom[5866] = 25'b1111111111111011110001100;
    rom[5867] = 25'b1111111111111011110000111;
    rom[5868] = 25'b1111111111111011110000011;
    rom[5869] = 25'b1111111111111011101111110;
    rom[5870] = 25'b1111111111111011101111001;
    rom[5871] = 25'b1111111111111011101110101;
    rom[5872] = 25'b1111111111111011101110000;
    rom[5873] = 25'b1111111111111011101101100;
    rom[5874] = 25'b1111111111111011101100111;
    rom[5875] = 25'b1111111111111011101100011;
    rom[5876] = 25'b1111111111111011101011110;
    rom[5877] = 25'b1111111111111011101011010;
    rom[5878] = 25'b1111111111111011101010101;
    rom[5879] = 25'b1111111111111011101010000;
    rom[5880] = 25'b1111111111111011101001100;
    rom[5881] = 25'b1111111111111011101000111;
    rom[5882] = 25'b1111111111111011101000011;
    rom[5883] = 25'b1111111111111011100111110;
    rom[5884] = 25'b1111111111111011100111010;
    rom[5885] = 25'b1111111111111011100110101;
    rom[5886] = 25'b1111111111111011100110001;
    rom[5887] = 25'b1111111111111011100101100;
    rom[5888] = 25'b1111111111111011100100111;
    rom[5889] = 25'b1111111111111011100100011;
    rom[5890] = 25'b1111111111111011100011110;
    rom[5891] = 25'b1111111111111011100011010;
    rom[5892] = 25'b1111111111111011100010101;
    rom[5893] = 25'b1111111111111011100010001;
    rom[5894] = 25'b1111111111111011100001100;
    rom[5895] = 25'b1111111111111011100001000;
    rom[5896] = 25'b1111111111111011100000011;
    rom[5897] = 25'b1111111111111011011111110;
    rom[5898] = 25'b1111111111111011011111001;
    rom[5899] = 25'b1111111111111011011110101;
    rom[5900] = 25'b1111111111111011011110001;
    rom[5901] = 25'b1111111111111011011101100;
    rom[5902] = 25'b1111111111111011011101000;
    rom[5903] = 25'b1111111111111011011100011;
    rom[5904] = 25'b1111111111111011011011111;
    rom[5905] = 25'b1111111111111011011011001;
    rom[5906] = 25'b1111111111111011011010101;
    rom[5907] = 25'b1111111111111011011010000;
    rom[5908] = 25'b1111111111111011011001100;
    rom[5909] = 25'b1111111111111011011000111;
    rom[5910] = 25'b1111111111111011011000011;
    rom[5911] = 25'b1111111111111011010111110;
    rom[5912] = 25'b1111111111111011010111010;
    rom[5913] = 25'b1111111111111011010110101;
    rom[5914] = 25'b1111111111111011010110000;
    rom[5915] = 25'b1111111111111011010101100;
    rom[5916] = 25'b1111111111111011010100111;
    rom[5917] = 25'b1111111111111011010100011;
    rom[5918] = 25'b1111111111111011010011110;
    rom[5919] = 25'b1111111111111011010011010;
    rom[5920] = 25'b1111111111111011010010101;
    rom[5921] = 25'b1111111111111011010010001;
    rom[5922] = 25'b1111111111111011010001100;
    rom[5923] = 25'b1111111111111011010000111;
    rom[5924] = 25'b1111111111111011010000011;
    rom[5925] = 25'b1111111111111011001111110;
    rom[5926] = 25'b1111111111111011001111010;
    rom[5927] = 25'b1111111111111011001110101;
    rom[5928] = 25'b1111111111111011001110001;
    rom[5929] = 25'b1111111111111011001101100;
    rom[5930] = 25'b1111111111111011001101000;
    rom[5931] = 25'b1111111111111011001100011;
    rom[5932] = 25'b1111111111111011001011110;
    rom[5933] = 25'b1111111111111011001011010;
    rom[5934] = 25'b1111111111111011001010101;
    rom[5935] = 25'b1111111111111011001010001;
    rom[5936] = 25'b1111111111111011001001100;
    rom[5937] = 25'b1111111111111011001001000;
    rom[5938] = 25'b1111111111111011001000011;
    rom[5939] = 25'b1111111111111011000111111;
    rom[5940] = 25'b1111111111111011000111001;
    rom[5941] = 25'b1111111111111011000110101;
    rom[5942] = 25'b1111111111111011000110001;
    rom[5943] = 25'b1111111111111011000101100;
    rom[5944] = 25'b1111111111111011000101000;
    rom[5945] = 25'b1111111111111011000100011;
    rom[5946] = 25'b1111111111111011000011111;
    rom[5947] = 25'b1111111111111011000011010;
    rom[5948] = 25'b1111111111111011000010110;
    rom[5949] = 25'b1111111111111011000010000;
    rom[5950] = 25'b1111111111111011000001100;
    rom[5951] = 25'b1111111111111011000000111;
    rom[5952] = 25'b1111111111111011000000011;
    rom[5953] = 25'b1111111111111010111111110;
    rom[5954] = 25'b1111111111111010111111010;
    rom[5955] = 25'b1111111111111010111110101;
    rom[5956] = 25'b1111111111111010111110001;
    rom[5957] = 25'b1111111111111010111101101;
    rom[5958] = 25'b1111111111111010111100111;
    rom[5959] = 25'b1111111111111010111100011;
    rom[5960] = 25'b1111111111111010111011110;
    rom[5961] = 25'b1111111111111010111011010;
    rom[5962] = 25'b1111111111111010111010101;
    rom[5963] = 25'b1111111111111010111010001;
    rom[5964] = 25'b1111111111111010111001100;
    rom[5965] = 25'b1111111111111010111001000;
    rom[5966] = 25'b1111111111111010111000011;
    rom[5967] = 25'b1111111111111010110111110;
    rom[5968] = 25'b1111111111111010110111010;
    rom[5969] = 25'b1111111111111010110110101;
    rom[5970] = 25'b1111111111111010110110001;
    rom[5971] = 25'b1111111111111010110101100;
    rom[5972] = 25'b1111111111111010110101000;
    rom[5973] = 25'b1111111111111010110100011;
    rom[5974] = 25'b1111111111111010110011111;
    rom[5975] = 25'b1111111111111010110011010;
    rom[5976] = 25'b1111111111111010110010110;
    rom[5977] = 25'b1111111111111010110010001;
    rom[5978] = 25'b1111111111111010110001100;
    rom[5979] = 25'b1111111111111010110001000;
    rom[5980] = 25'b1111111111111010110000011;
    rom[5981] = 25'b1111111111111010101111111;
    rom[5982] = 25'b1111111111111010101111010;
    rom[5983] = 25'b1111111111111010101110110;
    rom[5984] = 25'b1111111111111010101110001;
    rom[5985] = 25'b1111111111111010101101101;
    rom[5986] = 25'b1111111111111010101101000;
    rom[5987] = 25'b1111111111111010101100011;
    rom[5988] = 25'b1111111111111010101011111;
    rom[5989] = 25'b1111111111111010101011010;
    rom[5990] = 25'b1111111111111010101010110;
    rom[5991] = 25'b1111111111111010101010001;
    rom[5992] = 25'b1111111111111010101001101;
    rom[5993] = 25'b1111111111111010101001000;
    rom[5994] = 25'b1111111111111010101000100;
    rom[5995] = 25'b1111111111111010100111111;
    rom[5996] = 25'b1111111111111010100111011;
    rom[5997] = 25'b1111111111111010100110110;
    rom[5998] = 25'b1111111111111010100110001;
    rom[5999] = 25'b1111111111111010100101101;
    rom[6000] = 25'b1111111111111010100101000;
    rom[6001] = 25'b1111111111111010100100100;
    rom[6002] = 25'b1111111111111010100011111;
    rom[6003] = 25'b1111111111111010100011011;
    rom[6004] = 25'b1111111111111010100010110;
    rom[6005] = 25'b1111111111111010100010010;
    rom[6006] = 25'b1111111111111010100001101;
    rom[6007] = 25'b1111111111111010100001001;
    rom[6008] = 25'b1111111111111010100000100;
    rom[6009] = 25'b1111111111111010100000000;
    rom[6010] = 25'b1111111111111010011111011;
    rom[6011] = 25'b1111111111111010011110110;
    rom[6012] = 25'b1111111111111010011110001;
    rom[6013] = 25'b1111111111111010011101101;
    rom[6014] = 25'b1111111111111010011101001;
    rom[6015] = 25'b1111111111111010011100100;
    rom[6016] = 25'b1111111111111010011100000;
    rom[6017] = 25'b1111111111111010011011011;
    rom[6018] = 25'b1111111111111010011010111;
    rom[6019] = 25'b1111111111111010011010010;
    rom[6020] = 25'b1111111111111010011001110;
    rom[6021] = 25'b1111111111111010011001001;
    rom[6022] = 25'b1111111111111010011000101;
    rom[6023] = 25'b1111111111111010011000000;
    rom[6024] = 25'b1111111111111010010111100;
    rom[6025] = 25'b1111111111111010010110110;
    rom[6026] = 25'b1111111111111010010110010;
    rom[6027] = 25'b1111111111111010010101110;
    rom[6028] = 25'b1111111111111010010101001;
    rom[6029] = 25'b1111111111111010010100101;
    rom[6030] = 25'b1111111111111010010100000;
    rom[6031] = 25'b1111111111111010010011100;
    rom[6032] = 25'b1111111111111010010010111;
    rom[6033] = 25'b1111111111111010010010011;
    rom[6034] = 25'b1111111111111010010001110;
    rom[6035] = 25'b1111111111111010010001010;
    rom[6036] = 25'b1111111111111010010000101;
    rom[6037] = 25'b1111111111111010010000001;
    rom[6038] = 25'b1111111111111010001111100;
    rom[6039] = 25'b1111111111111010001111000;
    rom[6040] = 25'b1111111111111010001110011;
    rom[6041] = 25'b1111111111111010001101111;
    rom[6042] = 25'b1111111111111010001101010;
    rom[6043] = 25'b1111111111111010001100110;
    rom[6044] = 25'b1111111111111010001100001;
    rom[6045] = 25'b1111111111111010001011100;
    rom[6046] = 25'b1111111111111010001011000;
    rom[6047] = 25'b1111111111111010001010011;
    rom[6048] = 25'b1111111111111010001001111;
    rom[6049] = 25'b1111111111111010001001010;
    rom[6050] = 25'b1111111111111010001000110;
    rom[6051] = 25'b1111111111111010001000001;
    rom[6052] = 25'b1111111111111010000111101;
    rom[6053] = 25'b1111111111111010000111000;
    rom[6054] = 25'b1111111111111010000110100;
    rom[6055] = 25'b1111111111111010000101111;
    rom[6056] = 25'b1111111111111010000101011;
    rom[6057] = 25'b1111111111111010000100110;
    rom[6058] = 25'b1111111111111010000100010;
    rom[6059] = 25'b1111111111111010000011101;
    rom[6060] = 25'b1111111111111010000011001;
    rom[6061] = 25'b1111111111111010000010100;
    rom[6062] = 25'b1111111111111010000010000;
    rom[6063] = 25'b1111111111111010000001011;
    rom[6064] = 25'b1111111111111010000000111;
    rom[6065] = 25'b1111111111111010000000010;
    rom[6066] = 25'b1111111111111001111111110;
    rom[6067] = 25'b1111111111111001111111001;
    rom[6068] = 25'b1111111111111001111110101;
    rom[6069] = 25'b1111111111111001111110000;
    rom[6070] = 25'b1111111111111001111101100;
    rom[6071] = 25'b1111111111111001111101000;
    rom[6072] = 25'b1111111111111001111100011;
    rom[6073] = 25'b1111111111111001111011111;
    rom[6074] = 25'b1111111111111001111011010;
    rom[6075] = 25'b1111111111111001111010110;
    rom[6076] = 25'b1111111111111001111010001;
    rom[6077] = 25'b1111111111111001111001101;
    rom[6078] = 25'b1111111111111001111001000;
    rom[6079] = 25'b1111111111111001111000100;
    rom[6080] = 25'b1111111111111001110111111;
    rom[6081] = 25'b1111111111111001110111011;
    rom[6082] = 25'b1111111111111001110110110;
    rom[6083] = 25'b1111111111111001110110010;
    rom[6084] = 25'b1111111111111001110101101;
    rom[6085] = 25'b1111111111111001110101001;
    rom[6086] = 25'b1111111111111001110100100;
    rom[6087] = 25'b1111111111111001110100000;
    rom[6088] = 25'b1111111111111001110011011;
    rom[6089] = 25'b1111111111111001110010111;
    rom[6090] = 25'b1111111111111001110010010;
    rom[6091] = 25'b1111111111111001110001110;
    rom[6092] = 25'b1111111111111001110001001;
    rom[6093] = 25'b1111111111111001110000101;
    rom[6094] = 25'b1111111111111001110000000;
    rom[6095] = 25'b1111111111111001101111100;
    rom[6096] = 25'b1111111111111001101110111;
    rom[6097] = 25'b1111111111111001101110011;
    rom[6098] = 25'b1111111111111001101101111;
    rom[6099] = 25'b1111111111111001101101010;
    rom[6100] = 25'b1111111111111001101100110;
    rom[6101] = 25'b1111111111111001101100010;
    rom[6102] = 25'b1111111111111001101011101;
    rom[6103] = 25'b1111111111111001101011001;
    rom[6104] = 25'b1111111111111001101010100;
    rom[6105] = 25'b1111111111111001101010000;
    rom[6106] = 25'b1111111111111001101001011;
    rom[6107] = 25'b1111111111111001101000111;
    rom[6108] = 25'b1111111111111001101000010;
    rom[6109] = 25'b1111111111111001100111110;
    rom[6110] = 25'b1111111111111001100111001;
    rom[6111] = 25'b1111111111111001100110101;
    rom[6112] = 25'b1111111111111001100110000;
    rom[6113] = 25'b1111111111111001100101100;
    rom[6114] = 25'b1111111111111001100101000;
    rom[6115] = 25'b1111111111111001100100011;
    rom[6116] = 25'b1111111111111001100011111;
    rom[6117] = 25'b1111111111111001100011011;
    rom[6118] = 25'b1111111111111001100010110;
    rom[6119] = 25'b1111111111111001100010010;
    rom[6120] = 25'b1111111111111001100001101;
    rom[6121] = 25'b1111111111111001100001001;
    rom[6122] = 25'b1111111111111001100000100;
    rom[6123] = 25'b1111111111111001100000000;
    rom[6124] = 25'b1111111111111001011111011;
    rom[6125] = 25'b1111111111111001011110111;
    rom[6126] = 25'b1111111111111001011110010;
    rom[6127] = 25'b1111111111111001011101110;
    rom[6128] = 25'b1111111111111001011101010;
    rom[6129] = 25'b1111111111111001011100110;
    rom[6130] = 25'b1111111111111001011100001;
    rom[6131] = 25'b1111111111111001011011101;
    rom[6132] = 25'b1111111111111001011011000;
    rom[6133] = 25'b1111111111111001011010100;
    rom[6134] = 25'b1111111111111001011001111;
    rom[6135] = 25'b1111111111111001011001011;
    rom[6136] = 25'b1111111111111001011000110;
    rom[6137] = 25'b1111111111111001011000010;
    rom[6138] = 25'b1111111111111001010111110;
    rom[6139] = 25'b1111111111111001010111010;
    rom[6140] = 25'b1111111111111001010110101;
    rom[6141] = 25'b1111111111111001010110001;
    rom[6142] = 25'b1111111111111001010101100;
    rom[6143] = 25'b1111111111111001010101000;
    rom[6144] = 25'b1111111111111001010100011;
    rom[6145] = 25'b1111111111111001010011111;
    rom[6146] = 25'b1111111111111001010011011;
    rom[6147] = 25'b1111111111111001010010111;
    rom[6148] = 25'b1111111111111001010010010;
    rom[6149] = 25'b1111111111111001010001110;
    rom[6150] = 25'b1111111111111001010001001;
    rom[6151] = 25'b1111111111111001010000101;
    rom[6152] = 25'b1111111111111001010000000;
    rom[6153] = 25'b1111111111111001001111100;
    rom[6154] = 25'b1111111111111001001111000;
    rom[6155] = 25'b1111111111111001001110011;
    rom[6156] = 25'b1111111111111001001101111;
    rom[6157] = 25'b1111111111111001001101011;
    rom[6158] = 25'b1111111111111001001100110;
    rom[6159] = 25'b1111111111111001001100010;
    rom[6160] = 25'b1111111111111001001011110;
    rom[6161] = 25'b1111111111111001001011001;
    rom[6162] = 25'b1111111111111001001010101;
    rom[6163] = 25'b1111111111111001001010000;
    rom[6164] = 25'b1111111111111001001001100;
    rom[6165] = 25'b1111111111111001001001000;
    rom[6166] = 25'b1111111111111001001000100;
    rom[6167] = 25'b1111111111111001000111111;
    rom[6168] = 25'b1111111111111001000111011;
    rom[6169] = 25'b1111111111111001000110110;
    rom[6170] = 25'b1111111111111001000110010;
    rom[6171] = 25'b1111111111111001000101110;
    rom[6172] = 25'b1111111111111001000101010;
    rom[6173] = 25'b1111111111111001000100101;
    rom[6174] = 25'b1111111111111001000100001;
    rom[6175] = 25'b1111111111111001000011101;
    rom[6176] = 25'b1111111111111001000011000;
    rom[6177] = 25'b1111111111111001000010100;
    rom[6178] = 25'b1111111111111001000001111;
    rom[6179] = 25'b1111111111111001000001011;
    rom[6180] = 25'b1111111111111001000000111;
    rom[6181] = 25'b1111111111111001000000011;
    rom[6182] = 25'b1111111111111000111111110;
    rom[6183] = 25'b1111111111111000111111010;
    rom[6184] = 25'b1111111111111000111110110;
    rom[6185] = 25'b1111111111111000111110001;
    rom[6186] = 25'b1111111111111000111101101;
    rom[6187] = 25'b1111111111111000111101001;
    rom[6188] = 25'b1111111111111000111100101;
    rom[6189] = 25'b1111111111111000111100000;
    rom[6190] = 25'b1111111111111000111011100;
    rom[6191] = 25'b1111111111111000111010111;
    rom[6192] = 25'b1111111111111000111010100;
    rom[6193] = 25'b1111111111111000111001111;
    rom[6194] = 25'b1111111111111000111001011;
    rom[6195] = 25'b1111111111111000111000110;
    rom[6196] = 25'b1111111111111000111000010;
    rom[6197] = 25'b1111111111111000110111110;
    rom[6198] = 25'b1111111111111000110111001;
    rom[6199] = 25'b1111111111111000110110101;
    rom[6200] = 25'b1111111111111000110110001;
    rom[6201] = 25'b1111111111111000110101101;
    rom[6202] = 25'b1111111111111000110101000;
    rom[6203] = 25'b1111111111111000110100101;
    rom[6204] = 25'b1111111111111000110100000;
    rom[6205] = 25'b1111111111111000110011100;
    rom[6206] = 25'b1111111111111000110010111;
    rom[6207] = 25'b1111111111111000110010011;
    rom[6208] = 25'b1111111111111000110001111;
    rom[6209] = 25'b1111111111111000110001010;
    rom[6210] = 25'b1111111111111000110000111;
    rom[6211] = 25'b1111111111111000110000010;
    rom[6212] = 25'b1111111111111000101111110;
    rom[6213] = 25'b1111111111111000101111001;
    rom[6214] = 25'b1111111111111000101110101;
    rom[6215] = 25'b1111111111111000101110001;
    rom[6216] = 25'b1111111111111000101101101;
    rom[6217] = 25'b1111111111111000101101001;
    rom[6218] = 25'b1111111111111000101100100;
    rom[6219] = 25'b1111111111111000101100000;
    rom[6220] = 25'b1111111111111000101011100;
    rom[6221] = 25'b1111111111111000101011000;
    rom[6222] = 25'b1111111111111000101010011;
    rom[6223] = 25'b1111111111111000101001111;
    rom[6224] = 25'b1111111111111000101001011;
    rom[6225] = 25'b1111111111111000101000110;
    rom[6226] = 25'b1111111111111000101000011;
    rom[6227] = 25'b1111111111111000100111110;
    rom[6228] = 25'b1111111111111000100111010;
    rom[6229] = 25'b1111111111111000100110110;
    rom[6230] = 25'b1111111111111000100110001;
    rom[6231] = 25'b1111111111111000100101110;
    rom[6232] = 25'b1111111111111000100101001;
    rom[6233] = 25'b1111111111111000100100101;
    rom[6234] = 25'b1111111111111000100100001;
    rom[6235] = 25'b1111111111111000100011101;
    rom[6236] = 25'b1111111111111000100011001;
    rom[6237] = 25'b1111111111111000100010100;
    rom[6238] = 25'b1111111111111000100010000;
    rom[6239] = 25'b1111111111111000100001100;
    rom[6240] = 25'b1111111111111000100001000;
    rom[6241] = 25'b1111111111111000100000011;
    rom[6242] = 25'b1111111111111000011111111;
    rom[6243] = 25'b1111111111111000011111011;
    rom[6244] = 25'b1111111111111000011110111;
    rom[6245] = 25'b1111111111111000011110011;
    rom[6246] = 25'b1111111111111000011101111;
    rom[6247] = 25'b1111111111111000011101011;
    rom[6248] = 25'b1111111111111000011100110;
    rom[6249] = 25'b1111111111111000011100010;
    rom[6250] = 25'b1111111111111000011011110;
    rom[6251] = 25'b1111111111111000011011010;
    rom[6252] = 25'b1111111111111000011010110;
    rom[6253] = 25'b1111111111111000011010010;
    rom[6254] = 25'b1111111111111000011001101;
    rom[6255] = 25'b1111111111111000011001001;
    rom[6256] = 25'b1111111111111000011000101;
    rom[6257] = 25'b1111111111111000011000001;
    rom[6258] = 25'b1111111111111000010111101;
    rom[6259] = 25'b1111111111111000010111000;
    rom[6260] = 25'b1111111111111000010110101;
    rom[6261] = 25'b1111111111111000010110000;
    rom[6262] = 25'b1111111111111000010101100;
    rom[6263] = 25'b1111111111111000010101000;
    rom[6264] = 25'b1111111111111000010100100;
    rom[6265] = 25'b1111111111111000010100000;
    rom[6266] = 25'b1111111111111000010011100;
    rom[6267] = 25'b1111111111111000010011000;
    rom[6268] = 25'b1111111111111000010010100;
    rom[6269] = 25'b1111111111111000010001111;
    rom[6270] = 25'b1111111111111000010001100;
    rom[6271] = 25'b1111111111111000010000111;
    rom[6272] = 25'b1111111111111000010000011;
    rom[6273] = 25'b1111111111111000001111111;
    rom[6274] = 25'b1111111111111000001111011;
    rom[6275] = 25'b1111111111111000001110111;
    rom[6276] = 25'b1111111111111000001110011;
    rom[6277] = 25'b1111111111111000001101110;
    rom[6278] = 25'b1111111111111000001101011;
    rom[6279] = 25'b1111111111111000001100110;
    rom[6280] = 25'b1111111111111000001100011;
    rom[6281] = 25'b1111111111111000001011110;
    rom[6282] = 25'b1111111111111000001011010;
    rom[6283] = 25'b1111111111111000001010110;
    rom[6284] = 25'b1111111111111000001010010;
    rom[6285] = 25'b1111111111111000001001110;
    rom[6286] = 25'b1111111111111000001001010;
    rom[6287] = 25'b1111111111111000001000110;
    rom[6288] = 25'b1111111111111000001000010;
    rom[6289] = 25'b1111111111111000000111110;
    rom[6290] = 25'b1111111111111000000111001;
    rom[6291] = 25'b1111111111111000000110110;
    rom[6292] = 25'b1111111111111000000110001;
    rom[6293] = 25'b1111111111111000000101101;
    rom[6294] = 25'b1111111111111000000101010;
    rom[6295] = 25'b1111111111111000000100101;
    rom[6296] = 25'b1111111111111000000100010;
    rom[6297] = 25'b1111111111111000000011101;
    rom[6298] = 25'b1111111111111000000011001;
    rom[6299] = 25'b1111111111111000000010110;
    rom[6300] = 25'b1111111111111000000010001;
    rom[6301] = 25'b1111111111111000000001101;
    rom[6302] = 25'b1111111111111000000001010;
    rom[6303] = 25'b1111111111111000000000101;
    rom[6304] = 25'b1111111111111000000000001;
    rom[6305] = 25'b1111111111110111111111101;
    rom[6306] = 25'b1111111111110111111111001;
    rom[6307] = 25'b1111111111110111111110101;
    rom[6308] = 25'b1111111111110111111110001;
    rom[6309] = 25'b1111111111110111111101101;
    rom[6310] = 25'b1111111111110111111101010;
    rom[6311] = 25'b1111111111110111111100101;
    rom[6312] = 25'b1111111111110111111100001;
    rom[6313] = 25'b1111111111110111111011110;
    rom[6314] = 25'b1111111111110111111011001;
    rom[6315] = 25'b1111111111110111111010101;
    rom[6316] = 25'b1111111111110111111010010;
    rom[6317] = 25'b1111111111110111111001101;
    rom[6318] = 25'b1111111111110111111001001;
    rom[6319] = 25'b1111111111110111111000110;
    rom[6320] = 25'b1111111111110111111000001;
    rom[6321] = 25'b1111111111110111110111101;
    rom[6322] = 25'b1111111111110111110111010;
    rom[6323] = 25'b1111111111110111110110101;
    rom[6324] = 25'b1111111111110111110110001;
    rom[6325] = 25'b1111111111110111110101110;
    rom[6326] = 25'b1111111111110111110101010;
    rom[6327] = 25'b1111111111110111110100110;
    rom[6328] = 25'b1111111111110111110100010;
    rom[6329] = 25'b1111111111110111110011110;
    rom[6330] = 25'b1111111111110111110011010;
    rom[6331] = 25'b1111111111110111110010110;
    rom[6332] = 25'b1111111111110111110010010;
    rom[6333] = 25'b1111111111110111110001110;
    rom[6334] = 25'b1111111111110111110001010;
    rom[6335] = 25'b1111111111110111110000110;
    rom[6336] = 25'b1111111111110111110000010;
    rom[6337] = 25'b1111111111110111101111111;
    rom[6338] = 25'b1111111111110111101111011;
    rom[6339] = 25'b1111111111110111101110110;
    rom[6340] = 25'b1111111111110111101110011;
    rom[6341] = 25'b1111111111110111101101111;
    rom[6342] = 25'b1111111111110111101101011;
    rom[6343] = 25'b1111111111110111101100111;
    rom[6344] = 25'b1111111111110111101100011;
    rom[6345] = 25'b1111111111110111101011111;
    rom[6346] = 25'b1111111111110111101011100;
    rom[6347] = 25'b1111111111110111101011000;
    rom[6348] = 25'b1111111111110111101010011;
    rom[6349] = 25'b1111111111110111101010000;
    rom[6350] = 25'b1111111111110111101001100;
    rom[6351] = 25'b1111111111110111101001000;
    rom[6352] = 25'b1111111111110111101000100;
    rom[6353] = 25'b1111111111110111101000001;
    rom[6354] = 25'b1111111111110111100111100;
    rom[6355] = 25'b1111111111110111100111000;
    rom[6356] = 25'b1111111111110111100110101;
    rom[6357] = 25'b1111111111110111100110001;
    rom[6358] = 25'b1111111111110111100101101;
    rom[6359] = 25'b1111111111110111100101010;
    rom[6360] = 25'b1111111111110111100100110;
    rom[6361] = 25'b1111111111110111100100001;
    rom[6362] = 25'b1111111111110111100011110;
    rom[6363] = 25'b1111111111110111100011010;
    rom[6364] = 25'b1111111111110111100010110;
    rom[6365] = 25'b1111111111110111100010010;
    rom[6366] = 25'b1111111111110111100001111;
    rom[6367] = 25'b1111111111110111100001011;
    rom[6368] = 25'b1111111111110111100000111;
    rom[6369] = 25'b1111111111110111100000011;
    rom[6370] = 25'b1111111111110111100000000;
    rom[6371] = 25'b1111111111110111011111011;
    rom[6372] = 25'b1111111111110111011110111;
    rom[6373] = 25'b1111111111110111011110100;
    rom[6374] = 25'b1111111111110111011110000;
    rom[6375] = 25'b1111111111110111011101100;
    rom[6376] = 25'b1111111111110111011101001;
    rom[6377] = 25'b1111111111110111011100101;
    rom[6378] = 25'b1111111111110111011100001;
    rom[6379] = 25'b1111111111110111011011101;
    rom[6380] = 25'b1111111111110111011011010;
    rom[6381] = 25'b1111111111110111011010110;
    rom[6382] = 25'b1111111111110111011010010;
    rom[6383] = 25'b1111111111110111011001110;
    rom[6384] = 25'b1111111111110111011001011;
    rom[6385] = 25'b1111111111110111011000111;
    rom[6386] = 25'b1111111111110111011000011;
    rom[6387] = 25'b1111111111110111010111111;
    rom[6388] = 25'b1111111111110111010111100;
    rom[6389] = 25'b1111111111110111010111000;
    rom[6390] = 25'b1111111111110111010110100;
    rom[6391] = 25'b1111111111110111010110000;
    rom[6392] = 25'b1111111111110111010101101;
    rom[6393] = 25'b1111111111110111010101001;
    rom[6394] = 25'b1111111111110111010100101;
    rom[6395] = 25'b1111111111110111010100010;
    rom[6396] = 25'b1111111111110111010011110;
    rom[6397] = 25'b1111111111110111010011010;
    rom[6398] = 25'b1111111111110111010010110;
    rom[6399] = 25'b1111111111110111010010011;
    rom[6400] = 25'b1111111111110111010001111;
    rom[6401] = 25'b1111111111110111010001011;
    rom[6402] = 25'b1111111111110111010000111;
    rom[6403] = 25'b1111111111110111010000100;
    rom[6404] = 25'b1111111111110111010000000;
    rom[6405] = 25'b1111111111110111001111101;
    rom[6406] = 25'b1111111111110111001111001;
    rom[6407] = 25'b1111111111110111001110101;
    rom[6408] = 25'b1111111111110111001110010;
    rom[6409] = 25'b1111111111110111001101110;
    rom[6410] = 25'b1111111111110111001101010;
    rom[6411] = 25'b1111111111110111001100111;
    rom[6412] = 25'b1111111111110111001100011;
    rom[6413] = 25'b1111111111110111001011111;
    rom[6414] = 25'b1111111111110111001011100;
    rom[6415] = 25'b1111111111110111001011000;
    rom[6416] = 25'b1111111111110111001010101;
    rom[6417] = 25'b1111111111110111001010001;
    rom[6418] = 25'b1111111111110111001001101;
    rom[6419] = 25'b1111111111110111001001001;
    rom[6420] = 25'b1111111111110111001000110;
    rom[6421] = 25'b1111111111110111001000011;
    rom[6422] = 25'b1111111111110111000111111;
    rom[6423] = 25'b1111111111110111000111011;
    rom[6424] = 25'b1111111111110111000110111;
    rom[6425] = 25'b1111111111110111000110100;
    rom[6426] = 25'b1111111111110111000110001;
    rom[6427] = 25'b1111111111110111000101101;
    rom[6428] = 25'b1111111111110111000101001;
    rom[6429] = 25'b1111111111110111000100110;
    rom[6430] = 25'b1111111111110111000100010;
    rom[6431] = 25'b1111111111110111000011111;
    rom[6432] = 25'b1111111111110111000011011;
    rom[6433] = 25'b1111111111110111000010111;
    rom[6434] = 25'b1111111111110111000010100;
    rom[6435] = 25'b1111111111110111000010001;
    rom[6436] = 25'b1111111111110111000001101;
    rom[6437] = 25'b1111111111110111000001001;
    rom[6438] = 25'b1111111111110111000000101;
    rom[6439] = 25'b1111111111110111000000010;
    rom[6440] = 25'b1111111111110110111111111;
    rom[6441] = 25'b1111111111110110111111011;
    rom[6442] = 25'b1111111111110110111110111;
    rom[6443] = 25'b1111111111110110111110100;
    rom[6444] = 25'b1111111111110110111110000;
    rom[6445] = 25'b1111111111110110111101101;
    rom[6446] = 25'b1111111111110110111101010;
    rom[6447] = 25'b1111111111110110111100110;
    rom[6448] = 25'b1111111111110110111100010;
    rom[6449] = 25'b1111111111110110111011111;
    rom[6450] = 25'b1111111111110110111011100;
    rom[6451] = 25'b1111111111110110111011000;
    rom[6452] = 25'b1111111111110110111010100;
    rom[6453] = 25'b1111111111110110111010001;
    rom[6454] = 25'b1111111111110110111001101;
    rom[6455] = 25'b1111111111110110111001010;
    rom[6456] = 25'b1111111111110110111000111;
    rom[6457] = 25'b1111111111110110111000011;
    rom[6458] = 25'b1111111111110110111000000;
    rom[6459] = 25'b1111111111110110110111100;
    rom[6460] = 25'b1111111111110110110111000;
    rom[6461] = 25'b1111111111110110110110101;
    rom[6462] = 25'b1111111111110110110110010;
    rom[6463] = 25'b1111111111110110110101111;
    rom[6464] = 25'b1111111111110110110101011;
    rom[6465] = 25'b1111111111110110110100111;
    rom[6466] = 25'b1111111111110110110100100;
    rom[6467] = 25'b1111111111110110110100001;
    rom[6468] = 25'b1111111111110110110011110;
    rom[6469] = 25'b1111111111110110110011010;
    rom[6470] = 25'b1111111111110110110010111;
    rom[6471] = 25'b1111111111110110110010011;
    rom[6472] = 25'b1111111111110110110001111;
    rom[6473] = 25'b1111111111110110110001100;
    rom[6474] = 25'b1111111111110110110001001;
    rom[6475] = 25'b1111111111110110110000110;
    rom[6476] = 25'b1111111111110110110000010;
    rom[6477] = 25'b1111111111110110101111111;
    rom[6478] = 25'b1111111111110110101111011;
    rom[6479] = 25'b1111111111110110101111000;
    rom[6480] = 25'b1111111111110110101110100;
    rom[6481] = 25'b1111111111110110101110001;
    rom[6482] = 25'b1111111111110110101101110;
    rom[6483] = 25'b1111111111110110101101011;
    rom[6484] = 25'b1111111111110110101100111;
    rom[6485] = 25'b1111111111110110101100100;
    rom[6486] = 25'b1111111111110110101100000;
    rom[6487] = 25'b1111111111110110101011101;
    rom[6488] = 25'b1111111111110110101011010;
    rom[6489] = 25'b1111111111110110101010111;
    rom[6490] = 25'b1111111111110110101010100;
    rom[6491] = 25'b1111111111110110101010000;
    rom[6492] = 25'b1111111111110110101001101;
    rom[6493] = 25'b1111111111110110101001001;
    rom[6494] = 25'b1111111111110110101000110;
    rom[6495] = 25'b1111111111110110101000010;
    rom[6496] = 25'b1111111111110110100111111;
    rom[6497] = 25'b1111111111110110100111100;
    rom[6498] = 25'b1111111111110110100111001;
    rom[6499] = 25'b1111111111110110100110110;
    rom[6500] = 25'b1111111111110110100110010;
    rom[6501] = 25'b1111111111110110100101111;
    rom[6502] = 25'b1111111111110110100101100;
    rom[6503] = 25'b1111111111110110100101000;
    rom[6504] = 25'b1111111111110110100100101;
    rom[6505] = 25'b1111111111110110100100010;
    rom[6506] = 25'b1111111111110110100011111;
    rom[6507] = 25'b1111111111110110100011100;
    rom[6508] = 25'b1111111111110110100011001;
    rom[6509] = 25'b1111111111110110100010101;
    rom[6510] = 25'b1111111111110110100010010;
    rom[6511] = 25'b1111111111110110100001111;
    rom[6512] = 25'b1111111111110110100001011;
    rom[6513] = 25'b1111111111110110100001000;
    rom[6514] = 25'b1111111111110110100000101;
    rom[6515] = 25'b1111111111110110100000001;
    rom[6516] = 25'b1111111111110110011111110;
    rom[6517] = 25'b1111111111110110011111011;
    rom[6518] = 25'b1111111111110110011111000;
    rom[6519] = 25'b1111111111110110011110101;
    rom[6520] = 25'b1111111111110110011110010;
    rom[6521] = 25'b1111111111110110011101111;
    rom[6522] = 25'b1111111111110110011101100;
    rom[6523] = 25'b1111111111110110011101000;
    rom[6524] = 25'b1111111111110110011100101;
    rom[6525] = 25'b1111111111110110011100010;
    rom[6526] = 25'b1111111111110110011011111;
    rom[6527] = 25'b1111111111110110011011100;
    rom[6528] = 25'b1111111111110110011011000;
    rom[6529] = 25'b1111111111110110011010101;
    rom[6530] = 25'b1111111111110110011010010;
    rom[6531] = 25'b1111111111110110011001111;
    rom[6532] = 25'b1111111111110110011001100;
    rom[6533] = 25'b1111111111110110011001001;
    rom[6534] = 25'b1111111111110110011000110;
    rom[6535] = 25'b1111111111110110011000011;
    rom[6536] = 25'b1111111111110110011000000;
    rom[6537] = 25'b1111111111110110010111101;
    rom[6538] = 25'b1111111111110110010111010;
    rom[6539] = 25'b1111111111110110010110110;
    rom[6540] = 25'b1111111111110110010110011;
    rom[6541] = 25'b1111111111110110010110000;
    rom[6542] = 25'b1111111111110110010101101;
    rom[6543] = 25'b1111111111110110010101010;
    rom[6544] = 25'b1111111111110110010100111;
    rom[6545] = 25'b1111111111110110010100100;
    rom[6546] = 25'b1111111111110110010100001;
    rom[6547] = 25'b1111111111110110010011110;
    rom[6548] = 25'b1111111111110110010011011;
    rom[6549] = 25'b1111111111110110010011000;
    rom[6550] = 25'b1111111111110110010010100;
    rom[6551] = 25'b1111111111110110010010001;
    rom[6552] = 25'b1111111111110110010001110;
    rom[6553] = 25'b1111111111110110010001011;
    rom[6554] = 25'b1111111111110110010001000;
    rom[6555] = 25'b1111111111110110010000101;
    rom[6556] = 25'b1111111111110110010000010;
    rom[6557] = 25'b1111111111110110001111111;
    rom[6558] = 25'b1111111111110110001111100;
    rom[6559] = 25'b1111111111110110001111001;
    rom[6560] = 25'b1111111111110110001110110;
    rom[6561] = 25'b1111111111110110001110011;
    rom[6562] = 25'b1111111111110110001110000;
    rom[6563] = 25'b1111111111110110001101101;
    rom[6564] = 25'b1111111111110110001101010;
    rom[6565] = 25'b1111111111110110001100111;
    rom[6566] = 25'b1111111111110110001100101;
    rom[6567] = 25'b1111111111110110001100010;
    rom[6568] = 25'b1111111111110110001011111;
    rom[6569] = 25'b1111111111110110001011100;
    rom[6570] = 25'b1111111111110110001011001;
    rom[6571] = 25'b1111111111110110001010110;
    rom[6572] = 25'b1111111111110110001010011;
    rom[6573] = 25'b1111111111110110001010000;
    rom[6574] = 25'b1111111111110110001001101;
    rom[6575] = 25'b1111111111110110001001010;
    rom[6576] = 25'b1111111111110110001000111;
    rom[6577] = 25'b1111111111110110001000100;
    rom[6578] = 25'b1111111111110110001000010;
    rom[6579] = 25'b1111111111110110000111111;
    rom[6580] = 25'b1111111111110110000111100;
    rom[6581] = 25'b1111111111110110000111001;
    rom[6582] = 25'b1111111111110110000110110;
    rom[6583] = 25'b1111111111110110000110011;
    rom[6584] = 25'b1111111111110110000110000;
    rom[6585] = 25'b1111111111110110000101110;
    rom[6586] = 25'b1111111111110110000101011;
    rom[6587] = 25'b1111111111110110000101000;
    rom[6588] = 25'b1111111111110110000100101;
    rom[6589] = 25'b1111111111110110000100010;
    rom[6590] = 25'b1111111111110110000100000;
    rom[6591] = 25'b1111111111110110000011101;
    rom[6592] = 25'b1111111111110110000011010;
    rom[6593] = 25'b1111111111110110000010111;
    rom[6594] = 25'b1111111111110110000010101;
    rom[6595] = 25'b1111111111110110000010010;
    rom[6596] = 25'b1111111111110110000001111;
    rom[6597] = 25'b1111111111110110000001100;
    rom[6598] = 25'b1111111111110110000001001;
    rom[6599] = 25'b1111111111110110000000110;
    rom[6600] = 25'b1111111111110110000000011;
    rom[6601] = 25'b1111111111110110000000001;
    rom[6602] = 25'b1111111111110101111111110;
    rom[6603] = 25'b1111111111110101111111011;
    rom[6604] = 25'b1111111111110101111111000;
    rom[6605] = 25'b1111111111110101111110110;
    rom[6606] = 25'b1111111111110101111110011;
    rom[6607] = 25'b1111111111110101111110000;
    rom[6608] = 25'b1111111111110101111101110;
    rom[6609] = 25'b1111111111110101111101011;
    rom[6610] = 25'b1111111111110101111101000;
    rom[6611] = 25'b1111111111110101111100110;
    rom[6612] = 25'b1111111111110101111100011;
    rom[6613] = 25'b1111111111110101111100000;
    rom[6614] = 25'b1111111111110101111011101;
    rom[6615] = 25'b1111111111110101111011010;
    rom[6616] = 25'b1111111111110101111011000;
    rom[6617] = 25'b1111111111110101111010101;
    rom[6618] = 25'b1111111111110101111010011;
    rom[6619] = 25'b1111111111110101111010000;
    rom[6620] = 25'b1111111111110101111001110;
    rom[6621] = 25'b1111111111110101111001011;
    rom[6622] = 25'b1111111111110101111001000;
    rom[6623] = 25'b1111111111110101111000101;
    rom[6624] = 25'b1111111111110101111000010;
    rom[6625] = 25'b1111111111110101111000000;
    rom[6626] = 25'b1111111111110101110111101;
    rom[6627] = 25'b1111111111110101110111011;
    rom[6628] = 25'b1111111111110101110111000;
    rom[6629] = 25'b1111111111110101110110110;
    rom[6630] = 25'b1111111111110101110110011;
    rom[6631] = 25'b1111111111110101110110000;
    rom[6632] = 25'b1111111111110101110101101;
    rom[6633] = 25'b1111111111110101110101011;
    rom[6634] = 25'b1111111111110101110101000;
    rom[6635] = 25'b1111111111110101110100110;
    rom[6636] = 25'b1111111111110101110100100;
    rom[6637] = 25'b1111111111110101110100001;
    rom[6638] = 25'b1111111111110101110011111;
    rom[6639] = 25'b1111111111110101110011100;
    rom[6640] = 25'b1111111111110101110011001;
    rom[6641] = 25'b1111111111110101110010110;
    rom[6642] = 25'b1111111111110101110010100;
    rom[6643] = 25'b1111111111110101110010010;
    rom[6644] = 25'b1111111111110101110001111;
    rom[6645] = 25'b1111111111110101110001101;
    rom[6646] = 25'b1111111111110101110001010;
    rom[6647] = 25'b1111111111110101110000111;
    rom[6648] = 25'b1111111111110101110000101;
    rom[6649] = 25'b1111111111110101110000010;
    rom[6650] = 25'b1111111111110101110000000;
    rom[6651] = 25'b1111111111110101101111110;
    rom[6652] = 25'b1111111111110101101111011;
    rom[6653] = 25'b1111111111110101101111000;
    rom[6654] = 25'b1111111111110101101110110;
    rom[6655] = 25'b1111111111110101101110100;
    rom[6656] = 25'b1111111111110101101110001;
    rom[6657] = 25'b1111111111110101101101111;
    rom[6658] = 25'b1111111111110101101101100;
    rom[6659] = 25'b1111111111110101101101001;
    rom[6660] = 25'b1111111111110101101100111;
    rom[6661] = 25'b1111111111110101101100101;
    rom[6662] = 25'b1111111111110101101100011;
    rom[6663] = 25'b1111111111110101101100000;
    rom[6664] = 25'b1111111111110101101011110;
    rom[6665] = 25'b1111111111110101101011011;
    rom[6666] = 25'b1111111111110101101011001;
    rom[6667] = 25'b1111111111110101101010111;
    rom[6668] = 25'b1111111111110101101010100;
    rom[6669] = 25'b1111111111110101101010010;
    rom[6670] = 25'b1111111111110101101001111;
    rom[6671] = 25'b1111111111110101101001101;
    rom[6672] = 25'b1111111111110101101001011;
    rom[6673] = 25'b1111111111110101101001001;
    rom[6674] = 25'b1111111111110101101000110;
    rom[6675] = 25'b1111111111110101101000011;
    rom[6676] = 25'b1111111111110101101000001;
    rom[6677] = 25'b1111111111110101100111111;
    rom[6678] = 25'b1111111111110101100111101;
    rom[6679] = 25'b1111111111110101100111010;
    rom[6680] = 25'b1111111111110101100111000;
    rom[6681] = 25'b1111111111110101100110110;
    rom[6682] = 25'b1111111111110101100110100;
    rom[6683] = 25'b1111111111110101100110001;
    rom[6684] = 25'b1111111111110101100101110;
    rom[6685] = 25'b1111111111110101100101100;
    rom[6686] = 25'b1111111111110101100101010;
    rom[6687] = 25'b1111111111110101100101000;
    rom[6688] = 25'b1111111111110101100100101;
    rom[6689] = 25'b1111111111110101100100011;
    rom[6690] = 25'b1111111111110101100100001;
    rom[6691] = 25'b1111111111110101100011111;
    rom[6692] = 25'b1111111111110101100011101;
    rom[6693] = 25'b1111111111110101100011010;
    rom[6694] = 25'b1111111111110101100011000;
    rom[6695] = 25'b1111111111110101100010110;
    rom[6696] = 25'b1111111111110101100010100;
    rom[6697] = 25'b1111111111110101100010001;
    rom[6698] = 25'b1111111111110101100001111;
    rom[6699] = 25'b1111111111110101100001101;
    rom[6700] = 25'b1111111111110101100001011;
    rom[6701] = 25'b1111111111110101100001001;
    rom[6702] = 25'b1111111111110101100000111;
    rom[6703] = 25'b1111111111110101100000101;
    rom[6704] = 25'b1111111111110101100000010;
    rom[6705] = 25'b1111111111110101100000000;
    rom[6706] = 25'b1111111111110101011111110;
    rom[6707] = 25'b1111111111110101011111100;
    rom[6708] = 25'b1111111111110101011111001;
    rom[6709] = 25'b1111111111110101011110111;
    rom[6710] = 25'b1111111111110101011110110;
    rom[6711] = 25'b1111111111110101011110011;
    rom[6712] = 25'b1111111111110101011110001;
    rom[6713] = 25'b1111111111110101011101111;
    rom[6714] = 25'b1111111111110101011101101;
    rom[6715] = 25'b1111111111110101011101011;
    rom[6716] = 25'b1111111111110101011101001;
    rom[6717] = 25'b1111111111110101011100111;
    rom[6718] = 25'b1111111111110101011100101;
    rom[6719] = 25'b1111111111110101011100010;
    rom[6720] = 25'b1111111111110101011100001;
    rom[6721] = 25'b1111111111110101011011111;
    rom[6722] = 25'b1111111111110101011011100;
    rom[6723] = 25'b1111111111110101011011010;
    rom[6724] = 25'b1111111111110101011011001;
    rom[6725] = 25'b1111111111110101011010110;
    rom[6726] = 25'b1111111111110101011010100;
    rom[6727] = 25'b1111111111110101011010011;
    rom[6728] = 25'b1111111111110101011010000;
    rom[6729] = 25'b1111111111110101011001110;
    rom[6730] = 25'b1111111111110101011001100;
    rom[6731] = 25'b1111111111110101011001010;
    rom[6732] = 25'b1111111111110101011001000;
    rom[6733] = 25'b1111111111110101011000110;
    rom[6734] = 25'b1111111111110101011000100;
    rom[6735] = 25'b1111111111110101011000010;
    rom[6736] = 25'b1111111111110101011000001;
    rom[6737] = 25'b1111111111110101010111110;
    rom[6738] = 25'b1111111111110101010111100;
    rom[6739] = 25'b1111111111110101010111011;
    rom[6740] = 25'b1111111111110101010111000;
    rom[6741] = 25'b1111111111110101010110111;
    rom[6742] = 25'b1111111111110101010110101;
    rom[6743] = 25'b1111111111110101010110010;
    rom[6744] = 25'b1111111111110101010110001;
    rom[6745] = 25'b1111111111110101010101111;
    rom[6746] = 25'b1111111111110101010101101;
    rom[6747] = 25'b1111111111110101010101011;
    rom[6748] = 25'b1111111111110101010101001;
    rom[6749] = 25'b1111111111110101010100111;
    rom[6750] = 25'b1111111111110101010100110;
    rom[6751] = 25'b1111111111110101010100100;
    rom[6752] = 25'b1111111111110101010100010;
    rom[6753] = 25'b1111111111110101010100000;
    rom[6754] = 25'b1111111111110101010011110;
    rom[6755] = 25'b1111111111110101010011100;
    rom[6756] = 25'b1111111111110101010011011;
    rom[6757] = 25'b1111111111110101010011000;
    rom[6758] = 25'b1111111111110101010010111;
    rom[6759] = 25'b1111111111110101010010101;
    rom[6760] = 25'b1111111111110101010010011;
    rom[6761] = 25'b1111111111110101010010010;
    rom[6762] = 25'b1111111111110101010001111;
    rom[6763] = 25'b1111111111110101010001110;
    rom[6764] = 25'b1111111111110101010001100;
    rom[6765] = 25'b1111111111110101010001010;
    rom[6766] = 25'b1111111111110101010001001;
    rom[6767] = 25'b1111111111110101010000111;
    rom[6768] = 25'b1111111111110101010000101;
    rom[6769] = 25'b1111111111110101010000011;
    rom[6770] = 25'b1111111111110101010000010;
    rom[6771] = 25'b1111111111110101010000000;
    rom[6772] = 25'b1111111111110101001111110;
    rom[6773] = 25'b1111111111110101001111101;
    rom[6774] = 25'b1111111111110101001111010;
    rom[6775] = 25'b1111111111110101001111001;
    rom[6776] = 25'b1111111111110101001110111;
    rom[6777] = 25'b1111111111110101001110110;
    rom[6778] = 25'b1111111111110101001110100;
    rom[6779] = 25'b1111111111110101001110010;
    rom[6780] = 25'b1111111111110101001110001;
    rom[6781] = 25'b1111111111110101001101111;
    rom[6782] = 25'b1111111111110101001101101;
    rom[6783] = 25'b1111111111110101001101011;
    rom[6784] = 25'b1111111111110101001101010;
    rom[6785] = 25'b1111111111110101001101000;
    rom[6786] = 25'b1111111111110101001100111;
    rom[6787] = 25'b1111111111110101001100101;
    rom[6788] = 25'b1111111111110101001100011;
    rom[6789] = 25'b1111111111110101001100010;
    rom[6790] = 25'b1111111111110101001100000;
    rom[6791] = 25'b1111111111110101001011111;
    rom[6792] = 25'b1111111111110101001011101;
    rom[6793] = 25'b1111111111110101001011100;
    rom[6794] = 25'b1111111111110101001011010;
    rom[6795] = 25'b1111111111110101001011000;
    rom[6796] = 25'b1111111111110101001010111;
    rom[6797] = 25'b1111111111110101001010101;
    rom[6798] = 25'b1111111111110101001010100;
    rom[6799] = 25'b1111111111110101001010010;
    rom[6800] = 25'b1111111111110101001010001;
    rom[6801] = 25'b1111111111110101001001111;
    rom[6802] = 25'b1111111111110101001001110;
    rom[6803] = 25'b1111111111110101001001100;
    rom[6804] = 25'b1111111111110101001001011;
    rom[6805] = 25'b1111111111110101001001001;
    rom[6806] = 25'b1111111111110101001001000;
    rom[6807] = 25'b1111111111110101001000110;
    rom[6808] = 25'b1111111111110101001000101;
    rom[6809] = 25'b1111111111110101001000011;
    rom[6810] = 25'b1111111111110101001000010;
    rom[6811] = 25'b1111111111110101001000000;
    rom[6812] = 25'b1111111111110101000111111;
    rom[6813] = 25'b1111111111110101000111101;
    rom[6814] = 25'b1111111111110101000111100;
    rom[6815] = 25'b1111111111110101000111010;
    rom[6816] = 25'b1111111111110101000111001;
    rom[6817] = 25'b1111111111110101000111000;
    rom[6818] = 25'b1111111111110101000110110;
    rom[6819] = 25'b1111111111110101000110101;
    rom[6820] = 25'b1111111111110101000110011;
    rom[6821] = 25'b1111111111110101000110010;
    rom[6822] = 25'b1111111111110101000110000;
    rom[6823] = 25'b1111111111110101000110000;
    rom[6824] = 25'b1111111111110101000101110;
    rom[6825] = 25'b1111111111110101000101101;
    rom[6826] = 25'b1111111111110101000101011;
    rom[6827] = 25'b1111111111110101000101010;
    rom[6828] = 25'b1111111111110101000101001;
    rom[6829] = 25'b1111111111110101000100111;
    rom[6830] = 25'b1111111111110101000100110;
    rom[6831] = 25'b1111111111110101000100100;
    rom[6832] = 25'b1111111111110101000100011;
    rom[6833] = 25'b1111111111110101000100010;
    rom[6834] = 25'b1111111111110101000100001;
    rom[6835] = 25'b1111111111110101000011111;
    rom[6836] = 25'b1111111111110101000011111;
    rom[6837] = 25'b1111111111110101000011101;
    rom[6838] = 25'b1111111111110101000011100;
    rom[6839] = 25'b1111111111110101000011011;
    rom[6840] = 25'b1111111111110101000011001;
    rom[6841] = 25'b1111111111110101000011000;
    rom[6842] = 25'b1111111111110101000010111;
    rom[6843] = 25'b1111111111110101000010110;
    rom[6844] = 25'b1111111111110101000010100;
    rom[6845] = 25'b1111111111110101000010011;
    rom[6846] = 25'b1111111111110101000010010;
    rom[6847] = 25'b1111111111110101000010001;
    rom[6848] = 25'b1111111111110101000010000;
    rom[6849] = 25'b1111111111110101000001110;
    rom[6850] = 25'b1111111111110101000001101;
    rom[6851] = 25'b1111111111110101000001100;
    rom[6852] = 25'b1111111111110101000001011;
    rom[6853] = 25'b1111111111110101000001010;
    rom[6854] = 25'b1111111111110101000001001;
    rom[6855] = 25'b1111111111110101000000111;
    rom[6856] = 25'b1111111111110101000000111;
    rom[6857] = 25'b1111111111110101000000101;
    rom[6858] = 25'b1111111111110101000000100;
    rom[6859] = 25'b1111111111110101000000011;
    rom[6860] = 25'b1111111111110101000000010;
    rom[6861] = 25'b1111111111110101000000001;
    rom[6862] = 25'b1111111111110101000000000;
    rom[6863] = 25'b1111111111110100111111110;
    rom[6864] = 25'b1111111111110100111111110;
    rom[6865] = 25'b1111111111110100111111100;
    rom[6866] = 25'b1111111111110100111111011;
    rom[6867] = 25'b1111111111110100111111011;
    rom[6868] = 25'b1111111111110100111111001;
    rom[6869] = 25'b1111111111110100111111000;
    rom[6870] = 25'b1111111111110100111110111;
    rom[6871] = 25'b1111111111110100111110110;
    rom[6872] = 25'b1111111111110100111110101;
    rom[6873] = 25'b1111111111110100111110100;
    rom[6874] = 25'b1111111111110100111110011;
    rom[6875] = 25'b1111111111110100111110010;
    rom[6876] = 25'b1111111111110100111110001;
    rom[6877] = 25'b1111111111110100111110000;
    rom[6878] = 25'b1111111111110100111101111;
    rom[6879] = 25'b1111111111110100111101111;
    rom[6880] = 25'b1111111111110100111101101;
    rom[6881] = 25'b1111111111110100111101100;
    rom[6882] = 25'b1111111111110100111101100;
    rom[6883] = 25'b1111111111110100111101011;
    rom[6884] = 25'b1111111111110100111101001;
    rom[6885] = 25'b1111111111110100111101001;
    rom[6886] = 25'b1111111111110100111101000;
    rom[6887] = 25'b1111111111110100111100111;
    rom[6888] = 25'b1111111111110100111100110;
    rom[6889] = 25'b1111111111110100111100101;
    rom[6890] = 25'b1111111111110100111100100;
    rom[6891] = 25'b1111111111110100111100011;
    rom[6892] = 25'b1111111111110100111100011;
    rom[6893] = 25'b1111111111110100111100010;
    rom[6894] = 25'b1111111111110100111100001;
    rom[6895] = 25'b1111111111110100111100001;
    rom[6896] = 25'b1111111111110100111011111;
    rom[6897] = 25'b1111111111110100111011110;
    rom[6898] = 25'b1111111111110100111011110;
    rom[6899] = 25'b1111111111110100111011101;
    rom[6900] = 25'b1111111111110100111011100;
    rom[6901] = 25'b1111111111110100111011011;
    rom[6902] = 25'b1111111111110100111011011;
    rom[6903] = 25'b1111111111110100111011010;
    rom[6904] = 25'b1111111111110100111011001;
    rom[6905] = 25'b1111111111110100111011000;
    rom[6906] = 25'b1111111111110100111011000;
    rom[6907] = 25'b1111111111110100111010111;
    rom[6908] = 25'b1111111111110100111010110;
    rom[6909] = 25'b1111111111110100111010101;
    rom[6910] = 25'b1111111111110100111010101;
    rom[6911] = 25'b1111111111110100111010100;
    rom[6912] = 25'b1111111111110100111010011;
    rom[6913] = 25'b1111111111110100111010010;
    rom[6914] = 25'b1111111111110100111010010;
    rom[6915] = 25'b1111111111110100111010001;
    rom[6916] = 25'b1111111111110100111010000;
    rom[6917] = 25'b1111111111110100111010000;
    rom[6918] = 25'b1111111111110100111001111;
    rom[6919] = 25'b1111111111110100111001111;
    rom[6920] = 25'b1111111111110100111001110;
    rom[6921] = 25'b1111111111110100111001101;
    rom[6922] = 25'b1111111111110100111001100;
    rom[6923] = 25'b1111111111110100111001100;
    rom[6924] = 25'b1111111111110100111001100;
    rom[6925] = 25'b1111111111110100111001011;
    rom[6926] = 25'b1111111111110100111001010;
    rom[6927] = 25'b1111111111110100111001001;
    rom[6928] = 25'b1111111111110100111001001;
    rom[6929] = 25'b1111111111110100111001001;
    rom[6930] = 25'b1111111111110100111001000;
    rom[6931] = 25'b1111111111110100111000111;
    rom[6932] = 25'b1111111111110100111000111;
    rom[6933] = 25'b1111111111110100111000110;
    rom[6934] = 25'b1111111111110100111000110;
    rom[6935] = 25'b1111111111110100111000101;
    rom[6936] = 25'b1111111111110100111000101;
    rom[6937] = 25'b1111111111110100111000100;
    rom[6938] = 25'b1111111111110100111000011;
    rom[6939] = 25'b1111111111110100111000011;
    rom[6940] = 25'b1111111111110100111000011;
    rom[6941] = 25'b1111111111110100111000010;
    rom[6942] = 25'b1111111111110100111000010;
    rom[6943] = 25'b1111111111110100111000001;
    rom[6944] = 25'b1111111111110100111000001;
    rom[6945] = 25'b1111111111110100111000000;
    rom[6946] = 25'b1111111111110100111000000;
    rom[6947] = 25'b1111111111110100111000000;
    rom[6948] = 25'b1111111111110100110111111;
    rom[6949] = 25'b1111111111110100110111111;
    rom[6950] = 25'b1111111111110100110111110;
    rom[6951] = 25'b1111111111110100110111110;
    rom[6952] = 25'b1111111111110100110111101;
    rom[6953] = 25'b1111111111110100110111101;
    rom[6954] = 25'b1111111111110100110111101;
    rom[6955] = 25'b1111111111110100110111101;
    rom[6956] = 25'b1111111111110100110111100;
    rom[6957] = 25'b1111111111110100110111100;
    rom[6958] = 25'b1111111111110100110111011;
    rom[6959] = 25'b1111111111110100110111011;
    rom[6960] = 25'b1111111111110100110111010;
    rom[6961] = 25'b1111111111110100110111010;
    rom[6962] = 25'b1111111111110100110111010;
    rom[6963] = 25'b1111111111110100110111010;
    rom[6964] = 25'b1111111111110100110111010;
    rom[6965] = 25'b1111111111110100110111001;
    rom[6966] = 25'b1111111111110100110111001;
    rom[6967] = 25'b1111111111110100110111001;
    rom[6968] = 25'b1111111111110100110111000;
    rom[6969] = 25'b1111111111110100110111000;
    rom[6970] = 25'b1111111111110100110111000;
    rom[6971] = 25'b1111111111110100110110111;
    rom[6972] = 25'b1111111111110100110110111;
    rom[6973] = 25'b1111111111110100110110111;
    rom[6974] = 25'b1111111111110100110110111;
    rom[6975] = 25'b1111111111110100110110111;
    rom[6976] = 25'b1111111111110100110110111;
    rom[6977] = 25'b1111111111110100110110111;
    rom[6978] = 25'b1111111111110100110110111;
    rom[6979] = 25'b1111111111110100110110110;
    rom[6980] = 25'b1111111111110100110110110;
    rom[6981] = 25'b1111111111110100110110110;
    rom[6982] = 25'b1111111111110100110110110;
    rom[6983] = 25'b1111111111110100110110110;
    rom[6984] = 25'b1111111111110100110110101;
    rom[6985] = 25'b1111111111110100110110101;
    rom[6986] = 25'b1111111111110100110110101;
    rom[6987] = 25'b1111111111110100110110101;
    rom[6988] = 25'b1111111111110100110110101;
    rom[6989] = 25'b1111111111110100110110101;
    rom[6990] = 25'b1111111111110100110110101;
    rom[6991] = 25'b1111111111110100110110101;
    rom[6992] = 25'b1111111111110100110110100;
    rom[6993] = 25'b1111111111110100110110100;
    rom[6994] = 25'b1111111111110100110110100;
    rom[6995] = 25'b1111111111110100110110100;
    rom[6996] = 25'b1111111111110100110110100;
    rom[6997] = 25'b1111111111110100110110100;
    rom[6998] = 25'b1111111111110100110110100;
    rom[6999] = 25'b1111111111110100110110100;
    rom[7000] = 25'b1111111111110100110110100;
    rom[7001] = 25'b1111111111110100110110100;
    rom[7002] = 25'b1111111111110100110110100;
    rom[7003] = 25'b1111111111110100110110100;
    rom[7004] = 25'b1111111111110100110110100;
    rom[7005] = 25'b1111111111110100110110100;
    rom[7006] = 25'b1111111111110100110110101;
    rom[7007] = 25'b1111111111110100110110101;
    rom[7008] = 25'b1111111111110100110110101;
    rom[7009] = 25'b1111111111110100110110101;
    rom[7010] = 25'b1111111111110100110110101;
    rom[7011] = 25'b1111111111110100110110101;
    rom[7012] = 25'b1111111111110100110110101;
    rom[7013] = 25'b1111111111110100110110101;
    rom[7014] = 25'b1111111111110100110110110;
    rom[7015] = 25'b1111111111110100110110110;
    rom[7016] = 25'b1111111111110100110110110;
    rom[7017] = 25'b1111111111110100110110110;
    rom[7018] = 25'b1111111111110100110110110;
    rom[7019] = 25'b1111111111110100110110111;
    rom[7020] = 25'b1111111111110100110110111;
    rom[7021] = 25'b1111111111110100110110111;
    rom[7022] = 25'b1111111111110100110110111;
    rom[7023] = 25'b1111111111110100110110111;
    rom[7024] = 25'b1111111111110100110110111;
    rom[7025] = 25'b1111111111110100110110111;
    rom[7026] = 25'b1111111111110100110110111;
    rom[7027] = 25'b1111111111110100110111000;
    rom[7028] = 25'b1111111111110100110111000;
    rom[7029] = 25'b1111111111110100110111000;
    rom[7030] = 25'b1111111111110100110111001;
    rom[7031] = 25'b1111111111110100110111001;
    rom[7032] = 25'b1111111111110100110111010;
    rom[7033] = 25'b1111111111110100110111010;
    rom[7034] = 25'b1111111111110100110111010;
    rom[7035] = 25'b1111111111110100110111010;
    rom[7036] = 25'b1111111111110100110111010;
    rom[7037] = 25'b1111111111110100110111011;
    rom[7038] = 25'b1111111111110100110111011;
    rom[7039] = 25'b1111111111110100110111011;
    rom[7040] = 25'b1111111111110100110111100;
    rom[7041] = 25'b1111111111110100110111100;
    rom[7042] = 25'b1111111111110100110111101;
    rom[7043] = 25'b1111111111110100110111101;
    rom[7044] = 25'b1111111111110100110111101;
    rom[7045] = 25'b1111111111110100110111101;
    rom[7046] = 25'b1111111111110100110111110;
    rom[7047] = 25'b1111111111110100110111110;
    rom[7048] = 25'b1111111111110100110111111;
    rom[7049] = 25'b1111111111110100111000000;
    rom[7050] = 25'b1111111111110100111000000;
    rom[7051] = 25'b1111111111110100111000000;
    rom[7052] = 25'b1111111111110100111000000;
    rom[7053] = 25'b1111111111110100111000001;
    rom[7054] = 25'b1111111111110100111000010;
    rom[7055] = 25'b1111111111110100111000010;
    rom[7056] = 25'b1111111111110100111000011;
    rom[7057] = 25'b1111111111110100111000011;
    rom[7058] = 25'b1111111111110100111000011;
    rom[7059] = 25'b1111111111110100111000100;
    rom[7060] = 25'b1111111111110100111000101;
    rom[7061] = 25'b1111111111110100111000101;
    rom[7062] = 25'b1111111111110100111000110;
    rom[7063] = 25'b1111111111110100111000110;
    rom[7064] = 25'b1111111111110100111000111;
    rom[7065] = 25'b1111111111110100111000111;
    rom[7066] = 25'b1111111111110100111001000;
    rom[7067] = 25'b1111111111110100111001001;
    rom[7068] = 25'b1111111111110100111001001;
    rom[7069] = 25'b1111111111110100111001001;
    rom[7070] = 25'b1111111111110100111001010;
    rom[7071] = 25'b1111111111110100111001011;
    rom[7072] = 25'b1111111111110100111001100;
    rom[7073] = 25'b1111111111110100111001100;
    rom[7074] = 25'b1111111111110100111001101;
    rom[7075] = 25'b1111111111110100111001101;
    rom[7076] = 25'b1111111111110100111001110;
    rom[7077] = 25'b1111111111110100111001111;
    rom[7078] = 25'b1111111111110100111001111;
    rom[7079] = 25'b1111111111110100111010000;
    rom[7080] = 25'b1111111111110100111010001;
    rom[7081] = 25'b1111111111110100111010010;
    rom[7082] = 25'b1111111111110100111010010;
    rom[7083] = 25'b1111111111110100111010011;
    rom[7084] = 25'b1111111111110100111010100;
    rom[7085] = 25'b1111111111110100111010101;
    rom[7086] = 25'b1111111111110100111010101;
    rom[7087] = 25'b1111111111110100111010110;
    rom[7088] = 25'b1111111111110100111010111;
    rom[7089] = 25'b1111111111110100111011000;
    rom[7090] = 25'b1111111111110100111011000;
    rom[7091] = 25'b1111111111110100111011001;
    rom[7092] = 25'b1111111111110100111011010;
    rom[7093] = 25'b1111111111110100111011011;
    rom[7094] = 25'b1111111111110100111011011;
    rom[7095] = 25'b1111111111110100111011100;
    rom[7096] = 25'b1111111111110100111011110;
    rom[7097] = 25'b1111111111110100111011110;
    rom[7098] = 25'b1111111111110100111011111;
    rom[7099] = 25'b1111111111110100111100000;
    rom[7100] = 25'b1111111111110100111100001;
    rom[7101] = 25'b1111111111110100111100001;
    rom[7102] = 25'b1111111111110100111100010;
    rom[7103] = 25'b1111111111110100111100011;
    rom[7104] = 25'b1111111111110100111100100;
    rom[7105] = 25'b1111111111110100111100101;
    rom[7106] = 25'b1111111111110100111100110;
    rom[7107] = 25'b1111111111110100111100111;
    rom[7108] = 25'b1111111111110100111101000;
    rom[7109] = 25'b1111111111110100111101001;
    rom[7110] = 25'b1111111111110100111101001;
    rom[7111] = 25'b1111111111110100111101011;
    rom[7112] = 25'b1111111111110100111101100;
    rom[7113] = 25'b1111111111110100111101100;
    rom[7114] = 25'b1111111111110100111101110;
    rom[7115] = 25'b1111111111110100111101111;
    rom[7116] = 25'b1111111111110100111101111;
    rom[7117] = 25'b1111111111110100111110001;
    rom[7118] = 25'b1111111111110100111110010;
    rom[7119] = 25'b1111111111110100111110011;
    rom[7120] = 25'b1111111111110100111110100;
    rom[7121] = 25'b1111111111110100111110101;
    rom[7122] = 25'b1111111111110100111110110;
    rom[7123] = 25'b1111111111110100111110111;
    rom[7124] = 25'b1111111111110100111111000;
    rom[7125] = 25'b1111111111110100111111001;
    rom[7126] = 25'b1111111111110100111111011;
    rom[7127] = 25'b1111111111110100111111011;
    rom[7128] = 25'b1111111111110100111111101;
    rom[7129] = 25'b1111111111110100111111110;
    rom[7130] = 25'b1111111111110100111111111;
    rom[7131] = 25'b1111111111110101000000000;
    rom[7132] = 25'b1111111111110101000000001;
    rom[7133] = 25'b1111111111110101000000010;
    rom[7134] = 25'b1111111111110101000000100;
    rom[7135] = 25'b1111111111110101000000101;
    rom[7136] = 25'b1111111111110101000000110;
    rom[7137] = 25'b1111111111110101000000111;
    rom[7138] = 25'b1111111111110101000001000;
    rom[7139] = 25'b1111111111110101000001010;
    rom[7140] = 25'b1111111111110101000001011;
    rom[7141] = 25'b1111111111110101000001100;
    rom[7142] = 25'b1111111111110101000001101;
    rom[7143] = 25'b1111111111110101000001111;
    rom[7144] = 25'b1111111111110101000010000;
    rom[7145] = 25'b1111111111110101000010001;
    rom[7146] = 25'b1111111111110101000010011;
    rom[7147] = 25'b1111111111110101000010100;
    rom[7148] = 25'b1111111111110101000010101;
    rom[7149] = 25'b1111111111110101000010110;
    rom[7150] = 25'b1111111111110101000011000;
    rom[7151] = 25'b1111111111110101000011001;
    rom[7152] = 25'b1111111111110101000011010;
    rom[7153] = 25'b1111111111110101000011100;
    rom[7154] = 25'b1111111111110101000011101;
    rom[7155] = 25'b1111111111110101000011111;
    rom[7156] = 25'b1111111111110101000100000;
    rom[7157] = 25'b1111111111110101000100010;
    rom[7158] = 25'b1111111111110101000100011;
    rom[7159] = 25'b1111111111110101000100100;
    rom[7160] = 25'b1111111111110101000100101;
    rom[7161] = 25'b1111111111110101000100111;
    rom[7162] = 25'b1111111111110101000101000;
    rom[7163] = 25'b1111111111110101000101010;
    rom[7164] = 25'b1111111111110101000101011;
    rom[7165] = 25'b1111111111110101000101101;
    rom[7166] = 25'b1111111111110101000101110;
    rom[7167] = 25'b1111111111110101000110000;
    rom[7168] = 25'b1111111111110101000110001;
    rom[7169] = 25'b1111111111110101000110011;
    rom[7170] = 25'b1111111111110101000110100;
    rom[7171] = 25'b1111111111110101000110110;
    rom[7172] = 25'b1111111111110101000110111;
    rom[7173] = 25'b1111111111110101000111001;
    rom[7174] = 25'b1111111111110101000111010;
    rom[7175] = 25'b1111111111110101000111100;
    rom[7176] = 25'b1111111111110101000111101;
    rom[7177] = 25'b1111111111110101000111111;
    rom[7178] = 25'b1111111111110101001000001;
    rom[7179] = 25'b1111111111110101001000010;
    rom[7180] = 25'b1111111111110101001000100;
    rom[7181] = 25'b1111111111110101001000101;
    rom[7182] = 25'b1111111111110101001000111;
    rom[7183] = 25'b1111111111110101001001000;
    rom[7184] = 25'b1111111111110101001001011;
    rom[7185] = 25'b1111111111110101001001100;
    rom[7186] = 25'b1111111111110101001001110;
    rom[7187] = 25'b1111111111110101001001111;
    rom[7188] = 25'b1111111111110101001010001;
    rom[7189] = 25'b1111111111110101001010011;
    rom[7190] = 25'b1111111111110101001010100;
    rom[7191] = 25'b1111111111110101001010110;
    rom[7192] = 25'b1111111111110101001011000;
    rom[7193] = 25'b1111111111110101001011010;
    rom[7194] = 25'b1111111111110101001011011;
    rom[7195] = 25'b1111111111110101001011101;
    rom[7196] = 25'b1111111111110101001011111;
    rom[7197] = 25'b1111111111110101001100000;
    rom[7198] = 25'b1111111111110101001100011;
    rom[7199] = 25'b1111111111110101001100100;
    rom[7200] = 25'b1111111111110101001100101;
    rom[7201] = 25'b1111111111110101001101000;
    rom[7202] = 25'b1111111111110101001101001;
    rom[7203] = 25'b1111111111110101001101011;
    rom[7204] = 25'b1111111111110101001101101;
    rom[7205] = 25'b1111111111110101001101111;
    rom[7206] = 25'b1111111111110101001110001;
    rom[7207] = 25'b1111111111110101001110011;
    rom[7208] = 25'b1111111111110101001110100;
    rom[7209] = 25'b1111111111110101001110111;
    rom[7210] = 25'b1111111111110101001111000;
    rom[7211] = 25'b1111111111110101001111010;
    rom[7212] = 25'b1111111111110101001111100;
    rom[7213] = 25'b1111111111110101001111110;
    rom[7214] = 25'b1111111111110101010000000;
    rom[7215] = 25'b1111111111110101010000010;
    rom[7216] = 25'b1111111111110101010000011;
    rom[7217] = 25'b1111111111110101010000110;
    rom[7218] = 25'b1111111111110101010001000;
    rom[7219] = 25'b1111111111110101010001001;
    rom[7220] = 25'b1111111111110101010001100;
    rom[7221] = 25'b1111111111110101010001110;
    rom[7222] = 25'b1111111111110101010001111;
    rom[7223] = 25'b1111111111110101010010010;
    rom[7224] = 25'b1111111111110101010010100;
    rom[7225] = 25'b1111111111110101010010101;
    rom[7226] = 25'b1111111111110101010011000;
    rom[7227] = 25'b1111111111110101010011010;
    rom[7228] = 25'b1111111111110101010011100;
    rom[7229] = 25'b1111111111110101010011110;
    rom[7230] = 25'b1111111111110101010100000;
    rom[7231] = 25'b1111111111110101010100010;
    rom[7232] = 25'b1111111111110101010100100;
    rom[7233] = 25'b1111111111110101010100110;
    rom[7234] = 25'b1111111111110101010101000;
    rom[7235] = 25'b1111111111110101010101010;
    rom[7236] = 25'b1111111111110101010101100;
    rom[7237] = 25'b1111111111110101010101111;
    rom[7238] = 25'b1111111111110101010110001;
    rom[7239] = 25'b1111111111110101010110011;
    rom[7240] = 25'b1111111111110101010110101;
    rom[7241] = 25'b1111111111110101010111000;
    rom[7242] = 25'b1111111111110101010111001;
    rom[7243] = 25'b1111111111110101010111011;
    rom[7244] = 25'b1111111111110101010111110;
    rom[7245] = 25'b1111111111110101011000000;
    rom[7246] = 25'b1111111111110101011000010;
    rom[7247] = 25'b1111111111110101011000100;
    rom[7248] = 25'b1111111111110101011000111;
    rom[7249] = 25'b1111111111110101011001001;
    rom[7250] = 25'b1111111111110101011001011;
    rom[7251] = 25'b1111111111110101011001101;
    rom[7252] = 25'b1111111111110101011010000;
    rom[7253] = 25'b1111111111110101011010010;
    rom[7254] = 25'b1111111111110101011010101;
    rom[7255] = 25'b1111111111110101011010111;
    rom[7256] = 25'b1111111111110101011011001;
    rom[7257] = 25'b1111111111110101011011100;
    rom[7258] = 25'b1111111111110101011011110;
    rom[7259] = 25'b1111111111110101011100000;
    rom[7260] = 25'b1111111111110101011100010;
    rom[7261] = 25'b1111111111110101011100101;
    rom[7262] = 25'b1111111111110101011100111;
    rom[7263] = 25'b1111111111110101011101010;
    rom[7264] = 25'b1111111111110101011101100;
    rom[7265] = 25'b1111111111110101011101110;
    rom[7266] = 25'b1111111111110101011110001;
    rom[7267] = 25'b1111111111110101011110011;
    rom[7268] = 25'b1111111111110101011110110;
    rom[7269] = 25'b1111111111110101011111000;
    rom[7270] = 25'b1111111111110101011111011;
    rom[7271] = 25'b1111111111110101011111101;
    rom[7272] = 25'b1111111111110101011111111;
    rom[7273] = 25'b1111111111110101100000010;
    rom[7274] = 25'b1111111111110101100000101;
    rom[7275] = 25'b1111111111110101100000111;
    rom[7276] = 25'b1111111111110101100001010;
    rom[7277] = 25'b1111111111110101100001100;
    rom[7278] = 25'b1111111111110101100001110;
    rom[7279] = 25'b1111111111110101100010001;
    rom[7280] = 25'b1111111111110101100010100;
    rom[7281] = 25'b1111111111110101100010111;
    rom[7282] = 25'b1111111111110101100011001;
    rom[7283] = 25'b1111111111110101100011100;
    rom[7284] = 25'b1111111111110101100011110;
    rom[7285] = 25'b1111111111110101100100001;
    rom[7286] = 25'b1111111111110101100100011;
    rom[7287] = 25'b1111111111110101100100110;
    rom[7288] = 25'b1111111111110101100101000;
    rom[7289] = 25'b1111111111110101100101011;
    rom[7290] = 25'b1111111111110101100101110;
    rom[7291] = 25'b1111111111110101100110001;
    rom[7292] = 25'b1111111111110101100110011;
    rom[7293] = 25'b1111111111110101100110110;
    rom[7294] = 25'b1111111111110101100111000;
    rom[7295] = 25'b1111111111110101100111011;
    rom[7296] = 25'b1111111111110101100111110;
    rom[7297] = 25'b1111111111110101101000000;
    rom[7298] = 25'b1111111111110101101000011;
    rom[7299] = 25'b1111111111110101101000110;
    rom[7300] = 25'b1111111111110101101001001;
    rom[7301] = 25'b1111111111110101101001100;
    rom[7302] = 25'b1111111111110101101001111;
    rom[7303] = 25'b1111111111110101101010001;
    rom[7304] = 25'b1111111111110101101010100;
    rom[7305] = 25'b1111111111110101101010111;
    rom[7306] = 25'b1111111111110101101011010;
    rom[7307] = 25'b1111111111110101101011100;
    rom[7308] = 25'b1111111111110101101011111;
    rom[7309] = 25'b1111111111110101101100010;
    rom[7310] = 25'b1111111111110101101100101;
    rom[7311] = 25'b1111111111110101101101000;
    rom[7312] = 25'b1111111111110101101101011;
    rom[7313] = 25'b1111111111110101101101101;
    rom[7314] = 25'b1111111111110101101110000;
    rom[7315] = 25'b1111111111110101101110011;
    rom[7316] = 25'b1111111111110101101110110;
    rom[7317] = 25'b1111111111110101101111001;
    rom[7318] = 25'b1111111111110101101111100;
    rom[7319] = 25'b1111111111110101101111111;
    rom[7320] = 25'b1111111111110101110000010;
    rom[7321] = 25'b1111111111110101110000101;
    rom[7322] = 25'b1111111111110101110001000;
    rom[7323] = 25'b1111111111110101110001011;
    rom[7324] = 25'b1111111111110101110001110;
    rom[7325] = 25'b1111111111110101110010001;
    rom[7326] = 25'b1111111111110101110010100;
    rom[7327] = 25'b1111111111110101110010111;
    rom[7328] = 25'b1111111111110101110011010;
    rom[7329] = 25'b1111111111110101110011101;
    rom[7330] = 25'b1111111111110101110100000;
    rom[7331] = 25'b1111111111110101110100011;
    rom[7332] = 25'b1111111111110101110100110;
    rom[7333] = 25'b1111111111110101110101001;
    rom[7334] = 25'b1111111111110101110101100;
    rom[7335] = 25'b1111111111110101110101111;
    rom[7336] = 25'b1111111111110101110110011;
    rom[7337] = 25'b1111111111110101110110110;
    rom[7338] = 25'b1111111111110101110111001;
    rom[7339] = 25'b1111111111110101110111100;
    rom[7340] = 25'b1111111111110101110111111;
    rom[7341] = 25'b1111111111110101111000010;
    rom[7342] = 25'b1111111111110101111000101;
    rom[7343] = 25'b1111111111110101111001000;
    rom[7344] = 25'b1111111111110101111001011;
    rom[7345] = 25'b1111111111110101111001110;
    rom[7346] = 25'b1111111111110101111010010;
    rom[7347] = 25'b1111111111110101111010101;
    rom[7348] = 25'b1111111111110101111011000;
    rom[7349] = 25'b1111111111110101111011100;
    rom[7350] = 25'b1111111111110101111011111;
    rom[7351] = 25'b1111111111110101111100010;
    rom[7352] = 25'b1111111111110101111100110;
    rom[7353] = 25'b1111111111110101111101000;
    rom[7354] = 25'b1111111111110101111101100;
    rom[7355] = 25'b1111111111110101111101111;
    rom[7356] = 25'b1111111111110101111110010;
    rom[7357] = 25'b1111111111110101111110110;
    rom[7358] = 25'b1111111111110101111111001;
    rom[7359] = 25'b1111111111110101111111101;
    rom[7360] = 25'b1111111111110110000000000;
    rom[7361] = 25'b1111111111110110000000011;
    rom[7362] = 25'b1111111111110110000000110;
    rom[7363] = 25'b1111111111110110000001010;
    rom[7364] = 25'b1111111111110110000001101;
    rom[7365] = 25'b1111111111110110000010001;
    rom[7366] = 25'b1111111111110110000010100;
    rom[7367] = 25'b1111111111110110000011000;
    rom[7368] = 25'b1111111111110110000011011;
    rom[7369] = 25'b1111111111110110000011110;
    rom[7370] = 25'b1111111111110110000100010;
    rom[7371] = 25'b1111111111110110000100101;
    rom[7372] = 25'b1111111111110110000101001;
    rom[7373] = 25'b1111111111110110000101100;
    rom[7374] = 25'b1111111111110110000101111;
    rom[7375] = 25'b1111111111110110000110011;
    rom[7376] = 25'b1111111111110110000110110;
    rom[7377] = 25'b1111111111110110000111010;
    rom[7378] = 25'b1111111111110110000111110;
    rom[7379] = 25'b1111111111110110001000001;
    rom[7380] = 25'b1111111111110110001000100;
    rom[7381] = 25'b1111111111110110001001000;
    rom[7382] = 25'b1111111111110110001001100;
    rom[7383] = 25'b1111111111110110001010000;
    rom[7384] = 25'b1111111111110110001010011;
    rom[7385] = 25'b1111111111110110001010110;
    rom[7386] = 25'b1111111111110110001011010;
    rom[7387] = 25'b1111111111110110001011110;
    rom[7388] = 25'b1111111111110110001100010;
    rom[7389] = 25'b1111111111110110001100101;
    rom[7390] = 25'b1111111111110110001101000;
    rom[7391] = 25'b1111111111110110001101100;
    rom[7392] = 25'b1111111111110110001110000;
    rom[7393] = 25'b1111111111110110001110011;
    rom[7394] = 25'b1111111111110110001110111;
    rom[7395] = 25'b1111111111110110001111011;
    rom[7396] = 25'b1111111111110110001111111;
    rom[7397] = 25'b1111111111110110010000010;
    rom[7398] = 25'b1111111111110110010000110;
    rom[7399] = 25'b1111111111110110010001010;
    rom[7400] = 25'b1111111111110110010001110;
    rom[7401] = 25'b1111111111110110010010001;
    rom[7402] = 25'b1111111111110110010010101;
    rom[7403] = 25'b1111111111110110010011001;
    rom[7404] = 25'b1111111111110110010011101;
    rom[7405] = 25'b1111111111110110010100000;
    rom[7406] = 25'b1111111111110110010100100;
    rom[7407] = 25'b1111111111110110010101000;
    rom[7408] = 25'b1111111111110110010101011;
    rom[7409] = 25'b1111111111110110010101111;
    rom[7410] = 25'b1111111111110110010110100;
    rom[7411] = 25'b1111111111110110010110111;
    rom[7412] = 25'b1111111111110110010111011;
    rom[7413] = 25'b1111111111110110010111111;
    rom[7414] = 25'b1111111111110110011000011;
    rom[7415] = 25'b1111111111110110011000111;
    rom[7416] = 25'b1111111111110110011001011;
    rom[7417] = 25'b1111111111110110011001111;
    rom[7418] = 25'b1111111111110110011010010;
    rom[7419] = 25'b1111111111110110011010110;
    rom[7420] = 25'b1111111111110110011011011;
    rom[7421] = 25'b1111111111110110011011110;
    rom[7422] = 25'b1111111111110110011100010;
    rom[7423] = 25'b1111111111110110011100111;
    rom[7424] = 25'b1111111111110110011101010;
    rom[7425] = 25'b1111111111110110011101110;
    rom[7426] = 25'b1111111111110110011110010;
    rom[7427] = 25'b1111111111110110011110110;
    rom[7428] = 25'b1111111111110110011111010;
    rom[7429] = 25'b1111111111110110011111110;
    rom[7430] = 25'b1111111111110110100000010;
    rom[7431] = 25'b1111111111110110100000111;
    rom[7432] = 25'b1111111111110110100001010;
    rom[7433] = 25'b1111111111110110100001110;
    rom[7434] = 25'b1111111111110110100010011;
    rom[7435] = 25'b1111111111110110100010110;
    rom[7436] = 25'b1111111111110110100011011;
    rom[7437] = 25'b1111111111110110100011111;
    rom[7438] = 25'b1111111111110110100100011;
    rom[7439] = 25'b1111111111110110100100111;
    rom[7440] = 25'b1111111111110110100101011;
    rom[7441] = 25'b1111111111110110100110000;
    rom[7442] = 25'b1111111111110110100110011;
    rom[7443] = 25'b1111111111110110100111000;
    rom[7444] = 25'b1111111111110110100111100;
    rom[7445] = 25'b1111111111110110101000000;
    rom[7446] = 25'b1111111111110110101000101;
    rom[7447] = 25'b1111111111110110101001000;
    rom[7448] = 25'b1111111111110110101001101;
    rom[7449] = 25'b1111111111110110101010001;
    rom[7450] = 25'b1111111111110110101010101;
    rom[7451] = 25'b1111111111110110101011010;
    rom[7452] = 25'b1111111111110110101011110;
    rom[7453] = 25'b1111111111110110101100010;
    rom[7454] = 25'b1111111111110110101100110;
    rom[7455] = 25'b1111111111110110101101011;
    rom[7456] = 25'b1111111111110110101101110;
    rom[7457] = 25'b1111111111110110101110011;
    rom[7458] = 25'b1111111111110110101110111;
    rom[7459] = 25'b1111111111110110101111100;
    rom[7460] = 25'b1111111111110110110000000;
    rom[7461] = 25'b1111111111110110110000100;
    rom[7462] = 25'b1111111111110110110001001;
    rom[7463] = 25'b1111111111110110110001101;
    rom[7464] = 25'b1111111111110110110010010;
    rom[7465] = 25'b1111111111110110110010110;
    rom[7466] = 25'b1111111111110110110011011;
    rom[7467] = 25'b1111111111110110110011111;
    rom[7468] = 25'b1111111111110110110100100;
    rom[7469] = 25'b1111111111110110110101000;
    rom[7470] = 25'b1111111111110110110101100;
    rom[7471] = 25'b1111111111110110110110000;
    rom[7472] = 25'b1111111111110110110110101;
    rom[7473] = 25'b1111111111110110110111001;
    rom[7474] = 25'b1111111111110110110111110;
    rom[7475] = 25'b1111111111110110111000010;
    rom[7476] = 25'b1111111111110110111000111;
    rom[7477] = 25'b1111111111110110111001011;
    rom[7478] = 25'b1111111111110110111010000;
    rom[7479] = 25'b1111111111110110111010101;
    rom[7480] = 25'b1111111111110110111011001;
    rom[7481] = 25'b1111111111110110111011110;
    rom[7482] = 25'b1111111111110110111100010;
    rom[7483] = 25'b1111111111110110111100111;
    rom[7484] = 25'b1111111111110110111101011;
    rom[7485] = 25'b1111111111110110111110000;
    rom[7486] = 25'b1111111111110110111110100;
    rom[7487] = 25'b1111111111110110111111001;
    rom[7488] = 25'b1111111111110110111111110;
    rom[7489] = 25'b1111111111110111000000010;
    rom[7490] = 25'b1111111111110111000000111;
    rom[7491] = 25'b1111111111110111000001011;
    rom[7492] = 25'b1111111111110111000010001;
    rom[7493] = 25'b1111111111110111000010101;
    rom[7494] = 25'b1111111111110111000011010;
    rom[7495] = 25'b1111111111110111000011110;
    rom[7496] = 25'b1111111111110111000100011;
    rom[7497] = 25'b1111111111110111000101000;
    rom[7498] = 25'b1111111111110111000101100;
    rom[7499] = 25'b1111111111110111000110001;
    rom[7500] = 25'b1111111111110111000110110;
    rom[7501] = 25'b1111111111110111000111010;
    rom[7502] = 25'b1111111111110111001000000;
    rom[7503] = 25'b1111111111110111001000100;
    rom[7504] = 25'b1111111111110111001001001;
    rom[7505] = 25'b1111111111110111001001110;
    rom[7506] = 25'b1111111111110111001010010;
    rom[7507] = 25'b1111111111110111001011000;
    rom[7508] = 25'b1111111111110111001011100;
    rom[7509] = 25'b1111111111110111001100001;
    rom[7510] = 25'b1111111111110111001100110;
    rom[7511] = 25'b1111111111110111001101011;
    rom[7512] = 25'b1111111111110111001101111;
    rom[7513] = 25'b1111111111110111001110101;
    rom[7514] = 25'b1111111111110111001111001;
    rom[7515] = 25'b1111111111110111001111110;
    rom[7516] = 25'b1111111111110111010000100;
    rom[7517] = 25'b1111111111110111010001000;
    rom[7518] = 25'b1111111111110111010001101;
    rom[7519] = 25'b1111111111110111010010010;
    rom[7520] = 25'b1111111111110111010010111;
    rom[7521] = 25'b1111111111110111010011100;
    rom[7522] = 25'b1111111111110111010100001;
    rom[7523] = 25'b1111111111110111010100110;
    rom[7524] = 25'b1111111111110111010101011;
    rom[7525] = 25'b1111111111110111010110000;
    rom[7526] = 25'b1111111111110111010110101;
    rom[7527] = 25'b1111111111110111010111010;
    rom[7528] = 25'b1111111111110111010111111;
    rom[7529] = 25'b1111111111110111011000100;
    rom[7530] = 25'b1111111111110111011001001;
    rom[7531] = 25'b1111111111110111011001110;
    rom[7532] = 25'b1111111111110111011010011;
    rom[7533] = 25'b1111111111110111011011000;
    rom[7534] = 25'b1111111111110111011011101;
    rom[7535] = 25'b1111111111110111011100011;
    rom[7536] = 25'b1111111111110111011101000;
    rom[7537] = 25'b1111111111110111011101101;
    rom[7538] = 25'b1111111111110111011110001;
    rom[7539] = 25'b1111111111110111011110111;
    rom[7540] = 25'b1111111111110111011111100;
    rom[7541] = 25'b1111111111110111100000001;
    rom[7542] = 25'b1111111111110111100000110;
    rom[7543] = 25'b1111111111110111100001100;
    rom[7544] = 25'b1111111111110111100010001;
    rom[7545] = 25'b1111111111110111100010110;
    rom[7546] = 25'b1111111111110111100011011;
    rom[7547] = 25'b1111111111110111100100001;
    rom[7548] = 25'b1111111111110111100100110;
    rom[7549] = 25'b1111111111110111100101011;
    rom[7550] = 25'b1111111111110111100110000;
    rom[7551] = 25'b1111111111110111100110101;
    rom[7552] = 25'b1111111111110111100111011;
    rom[7553] = 25'b1111111111110111101000000;
    rom[7554] = 25'b1111111111110111101000101;
    rom[7555] = 25'b1111111111110111101001010;
    rom[7556] = 25'b1111111111110111101010000;
    rom[7557] = 25'b1111111111110111101010101;
    rom[7558] = 25'b1111111111110111101011011;
    rom[7559] = 25'b1111111111110111101100000;
    rom[7560] = 25'b1111111111110111101100101;
    rom[7561] = 25'b1111111111110111101101010;
    rom[7562] = 25'b1111111111110111101110000;
    rom[7563] = 25'b1111111111110111101110101;
    rom[7564] = 25'b1111111111110111101111011;
    rom[7565] = 25'b1111111111110111110000000;
    rom[7566] = 25'b1111111111110111110000101;
    rom[7567] = 25'b1111111111110111110001011;
    rom[7568] = 25'b1111111111110111110010001;
    rom[7569] = 25'b1111111111110111110010110;
    rom[7570] = 25'b1111111111110111110011011;
    rom[7571] = 25'b1111111111110111110100000;
    rom[7572] = 25'b1111111111110111110100110;
    rom[7573] = 25'b1111111111110111110101011;
    rom[7574] = 25'b1111111111110111110110001;
    rom[7575] = 25'b1111111111110111110110111;
    rom[7576] = 25'b1111111111110111110111100;
    rom[7577] = 25'b1111111111110111111000010;
    rom[7578] = 25'b1111111111110111111000111;
    rom[7579] = 25'b1111111111110111111001100;
    rom[7580] = 25'b1111111111110111111010010;
    rom[7581] = 25'b1111111111110111111011000;
    rom[7582] = 25'b1111111111110111111011110;
    rom[7583] = 25'b1111111111110111111100011;
    rom[7584] = 25'b1111111111110111111101001;
    rom[7585] = 25'b1111111111110111111101110;
    rom[7586] = 25'b1111111111110111111110100;
    rom[7587] = 25'b1111111111110111111111001;
    rom[7588] = 25'b1111111111110111111111111;
    rom[7589] = 25'b1111111111111000000000100;
    rom[7590] = 25'b1111111111111000000001010;
    rom[7591] = 25'b1111111111111000000010000;
    rom[7592] = 25'b1111111111111000000010110;
    rom[7593] = 25'b1111111111111000000011100;
    rom[7594] = 25'b1111111111111000000100001;
    rom[7595] = 25'b1111111111111000000100111;
    rom[7596] = 25'b1111111111111000000101101;
    rom[7597] = 25'b1111111111111000000110010;
    rom[7598] = 25'b1111111111111000000111000;
    rom[7599] = 25'b1111111111111000000111110;
    rom[7600] = 25'b1111111111111000001000011;
    rom[7601] = 25'b1111111111111000001001001;
    rom[7602] = 25'b1111111111111000001001111;
    rom[7603] = 25'b1111111111111000001010101;
    rom[7604] = 25'b1111111111111000001011010;
    rom[7605] = 25'b1111111111111000001100000;
    rom[7606] = 25'b1111111111111000001100110;
    rom[7607] = 25'b1111111111111000001101100;
    rom[7608] = 25'b1111111111111000001110001;
    rom[7609] = 25'b1111111111111000001110111;
    rom[7610] = 25'b1111111111111000001111101;
    rom[7611] = 25'b1111111111111000010000011;
    rom[7612] = 25'b1111111111111000010001001;
    rom[7613] = 25'b1111111111111000010001111;
    rom[7614] = 25'b1111111111111000010010101;
    rom[7615] = 25'b1111111111111000010011011;
    rom[7616] = 25'b1111111111111000010100001;
    rom[7617] = 25'b1111111111111000010100111;
    rom[7618] = 25'b1111111111111000010101100;
    rom[7619] = 25'b1111111111111000010110010;
    rom[7620] = 25'b1111111111111000010111000;
    rom[7621] = 25'b1111111111111000010111110;
    rom[7622] = 25'b1111111111111000011000100;
    rom[7623] = 25'b1111111111111000011001010;
    rom[7624] = 25'b1111111111111000011010000;
    rom[7625] = 25'b1111111111111000011010110;
    rom[7626] = 25'b1111111111111000011011100;
    rom[7627] = 25'b1111111111111000011100010;
    rom[7628] = 25'b1111111111111000011101000;
    rom[7629] = 25'b1111111111111000011101111;
    rom[7630] = 25'b1111111111111000011110101;
    rom[7631] = 25'b1111111111111000011111011;
    rom[7632] = 25'b1111111111111000100000001;
    rom[7633] = 25'b1111111111111000100000111;
    rom[7634] = 25'b1111111111111000100001101;
    rom[7635] = 25'b1111111111111000100010011;
    rom[7636] = 25'b1111111111111000100011010;
    rom[7637] = 25'b1111111111111000100100000;
    rom[7638] = 25'b1111111111111000100100110;
    rom[7639] = 25'b1111111111111000100101100;
    rom[7640] = 25'b1111111111111000100110001;
    rom[7641] = 25'b1111111111111000100111000;
    rom[7642] = 25'b1111111111111000100111110;
    rom[7643] = 25'b1111111111111000101000100;
    rom[7644] = 25'b1111111111111000101001010;
    rom[7645] = 25'b1111111111111000101010001;
    rom[7646] = 25'b1111111111111000101010111;
    rom[7647] = 25'b1111111111111000101011101;
    rom[7648] = 25'b1111111111111000101100100;
    rom[7649] = 25'b1111111111111000101101010;
    rom[7650] = 25'b1111111111111000101110000;
    rom[7651] = 25'b1111111111111000101110110;
    rom[7652] = 25'b1111111111111000101111100;
    rom[7653] = 25'b1111111111111000110000011;
    rom[7654] = 25'b1111111111111000110001001;
    rom[7655] = 25'b1111111111111000110010000;
    rom[7656] = 25'b1111111111111000110010110;
    rom[7657] = 25'b1111111111111000110011100;
    rom[7658] = 25'b1111111111111000110100010;
    rom[7659] = 25'b1111111111111000110101000;
    rom[7660] = 25'b1111111111111000110101111;
    rom[7661] = 25'b1111111111111000110110101;
    rom[7662] = 25'b1111111111111000110111100;
    rom[7663] = 25'b1111111111111000111000010;
    rom[7664] = 25'b1111111111111000111001000;
    rom[7665] = 25'b1111111111111000111001111;
    rom[7666] = 25'b1111111111111000111010101;
    rom[7667] = 25'b1111111111111000111011100;
    rom[7668] = 25'b1111111111111000111100010;
    rom[7669] = 25'b1111111111111000111101001;
    rom[7670] = 25'b1111111111111000111101111;
    rom[7671] = 25'b1111111111111000111110101;
    rom[7672] = 25'b1111111111111000111111100;
    rom[7673] = 25'b1111111111111001000000011;
    rom[7674] = 25'b1111111111111001000001001;
    rom[7675] = 25'b1111111111111001000001111;
    rom[7676] = 25'b1111111111111001000010110;
    rom[7677] = 25'b1111111111111001000011101;
    rom[7678] = 25'b1111111111111001000100011;
    rom[7679] = 25'b1111111111111001000101010;
    rom[7680] = 25'b1111111111111001000110000;
    rom[7681] = 25'b1111111111111001000110111;
    rom[7682] = 25'b1111111111111001000111101;
    rom[7683] = 25'b1111111111111001001000100;
    rom[7684] = 25'b1111111111111001001001010;
    rom[7685] = 25'b1111111111111001001010001;
    rom[7686] = 25'b1111111111111001001011000;
    rom[7687] = 25'b1111111111111001001011111;
    rom[7688] = 25'b1111111111111001001100101;
    rom[7689] = 25'b1111111111111001001101011;
    rom[7690] = 25'b1111111111111001001110010;
    rom[7691] = 25'b1111111111111001001111001;
    rom[7692] = 25'b1111111111111001001111111;
    rom[7693] = 25'b1111111111111001010000110;
    rom[7694] = 25'b1111111111111001010001101;
    rom[7695] = 25'b1111111111111001010010100;
    rom[7696] = 25'b1111111111111001010011010;
    rom[7697] = 25'b1111111111111001010100001;
    rom[7698] = 25'b1111111111111001010101000;
    rom[7699] = 25'b1111111111111001010101111;
    rom[7700] = 25'b1111111111111001010110101;
    rom[7701] = 25'b1111111111111001010111100;
    rom[7702] = 25'b1111111111111001011000011;
    rom[7703] = 25'b1111111111111001011001001;
    rom[7704] = 25'b1111111111111001011010000;
    rom[7705] = 25'b1111111111111001011010111;
    rom[7706] = 25'b1111111111111001011011110;
    rom[7707] = 25'b1111111111111001011100101;
    rom[7708] = 25'b1111111111111001011101100;
    rom[7709] = 25'b1111111111111001011110010;
    rom[7710] = 25'b1111111111111001011111001;
    rom[7711] = 25'b1111111111111001100000000;
    rom[7712] = 25'b1111111111111001100000111;
    rom[7713] = 25'b1111111111111001100001110;
    rom[7714] = 25'b1111111111111001100010101;
    rom[7715] = 25'b1111111111111001100011100;
    rom[7716] = 25'b1111111111111001100100010;
    rom[7717] = 25'b1111111111111001100101010;
    rom[7718] = 25'b1111111111111001100110000;
    rom[7719] = 25'b1111111111111001100110111;
    rom[7720] = 25'b1111111111111001100111110;
    rom[7721] = 25'b1111111111111001101000101;
    rom[7722] = 25'b1111111111111001101001100;
    rom[7723] = 25'b1111111111111001101010011;
    rom[7724] = 25'b1111111111111001101011010;
    rom[7725] = 25'b1111111111111001101100001;
    rom[7726] = 25'b1111111111111001101101001;
    rom[7727] = 25'b1111111111111001101101111;
    rom[7728] = 25'b1111111111111001101110110;
    rom[7729] = 25'b1111111111111001101111101;
    rom[7730] = 25'b1111111111111001110000100;
    rom[7731] = 25'b1111111111111001110001100;
    rom[7732] = 25'b1111111111111001110010010;
    rom[7733] = 25'b1111111111111001110011010;
    rom[7734] = 25'b1111111111111001110100001;
    rom[7735] = 25'b1111111111111001110101000;
    rom[7736] = 25'b1111111111111001110101111;
    rom[7737] = 25'b1111111111111001110110110;
    rom[7738] = 25'b1111111111111001110111101;
    rom[7739] = 25'b1111111111111001111000100;
    rom[7740] = 25'b1111111111111001111001011;
    rom[7741] = 25'b1111111111111001111010011;
    rom[7742] = 25'b1111111111111001111011001;
    rom[7743] = 25'b1111111111111001111100001;
    rom[7744] = 25'b1111111111111001111101000;
    rom[7745] = 25'b1111111111111001111101111;
    rom[7746] = 25'b1111111111111001111110110;
    rom[7747] = 25'b1111111111111001111111101;
    rom[7748] = 25'b1111111111111010000000101;
    rom[7749] = 25'b1111111111111010000001100;
    rom[7750] = 25'b1111111111111010000010100;
    rom[7751] = 25'b1111111111111010000011010;
    rom[7752] = 25'b1111111111111010000100010;
    rom[7753] = 25'b1111111111111010000101001;
    rom[7754] = 25'b1111111111111010000110000;
    rom[7755] = 25'b1111111111111010000110111;
    rom[7756] = 25'b1111111111111010000111111;
    rom[7757] = 25'b1111111111111010001000110;
    rom[7758] = 25'b1111111111111010001001101;
    rom[7759] = 25'b1111111111111010001010101;
    rom[7760] = 25'b1111111111111010001011100;
    rom[7761] = 25'b1111111111111010001100100;
    rom[7762] = 25'b1111111111111010001101011;
    rom[7763] = 25'b1111111111111010001110010;
    rom[7764] = 25'b1111111111111010001111010;
    rom[7765] = 25'b1111111111111010010000001;
    rom[7766] = 25'b1111111111111010010001000;
    rom[7767] = 25'b1111111111111010010010000;
    rom[7768] = 25'b1111111111111010010010111;
    rom[7769] = 25'b1111111111111010010011111;
    rom[7770] = 25'b1111111111111010010100110;
    rom[7771] = 25'b1111111111111010010101110;
    rom[7772] = 25'b1111111111111010010110101;
    rom[7773] = 25'b1111111111111010010111100;
    rom[7774] = 25'b1111111111111010011000100;
    rom[7775] = 25'b1111111111111010011001011;
    rom[7776] = 25'b1111111111111010011010011;
    rom[7777] = 25'b1111111111111010011011010;
    rom[7778] = 25'b1111111111111010011100010;
    rom[7779] = 25'b1111111111111010011101001;
    rom[7780] = 25'b1111111111111010011110001;
    rom[7781] = 25'b1111111111111010011111000;
    rom[7782] = 25'b1111111111111010100000000;
    rom[7783] = 25'b1111111111111010100000111;
    rom[7784] = 25'b1111111111111010100001111;
    rom[7785] = 25'b1111111111111010100010111;
    rom[7786] = 25'b1111111111111010100011110;
    rom[7787] = 25'b1111111111111010100100110;
    rom[7788] = 25'b1111111111111010100101101;
    rom[7789] = 25'b1111111111111010100110101;
    rom[7790] = 25'b1111111111111010100111101;
    rom[7791] = 25'b1111111111111010101000100;
    rom[7792] = 25'b1111111111111010101001100;
    rom[7793] = 25'b1111111111111010101010011;
    rom[7794] = 25'b1111111111111010101011100;
    rom[7795] = 25'b1111111111111010101100011;
    rom[7796] = 25'b1111111111111010101101011;
    rom[7797] = 25'b1111111111111010101110010;
    rom[7798] = 25'b1111111111111010101111010;
    rom[7799] = 25'b1111111111111010110000010;
    rom[7800] = 25'b1111111111111010110001001;
    rom[7801] = 25'b1111111111111010110010001;
    rom[7802] = 25'b1111111111111010110011001;
    rom[7803] = 25'b1111111111111010110100000;
    rom[7804] = 25'b1111111111111010110101001;
    rom[7805] = 25'b1111111111111010110110000;
    rom[7806] = 25'b1111111111111010110111000;
    rom[7807] = 25'b1111111111111010111000000;
    rom[7808] = 25'b1111111111111010111000111;
    rom[7809] = 25'b1111111111111010111001111;
    rom[7810] = 25'b1111111111111010111010111;
    rom[7811] = 25'b1111111111111010111011111;
    rom[7812] = 25'b1111111111111010111100111;
    rom[7813] = 25'b1111111111111010111101111;
    rom[7814] = 25'b1111111111111010111110110;
    rom[7815] = 25'b1111111111111010111111110;
    rom[7816] = 25'b1111111111111011000000110;
    rom[7817] = 25'b1111111111111011000001110;
    rom[7818] = 25'b1111111111111011000010110;
    rom[7819] = 25'b1111111111111011000011110;
    rom[7820] = 25'b1111111111111011000100110;
    rom[7821] = 25'b1111111111111011000101110;
    rom[7822] = 25'b1111111111111011000110110;
    rom[7823] = 25'b1111111111111011000111101;
    rom[7824] = 25'b1111111111111011001000101;
    rom[7825] = 25'b1111111111111011001001110;
    rom[7826] = 25'b1111111111111011001010101;
    rom[7827] = 25'b1111111111111011001011101;
    rom[7828] = 25'b1111111111111011001100110;
    rom[7829] = 25'b1111111111111011001101101;
    rom[7830] = 25'b1111111111111011001110101;
    rom[7831] = 25'b1111111111111011001111101;
    rom[7832] = 25'b1111111111111011010000110;
    rom[7833] = 25'b1111111111111011010001101;
    rom[7834] = 25'b1111111111111011010010101;
    rom[7835] = 25'b1111111111111011010011110;
    rom[7836] = 25'b1111111111111011010100110;
    rom[7837] = 25'b1111111111111011010101101;
    rom[7838] = 25'b1111111111111011010110101;
    rom[7839] = 25'b1111111111111011010111110;
    rom[7840] = 25'b1111111111111011011000110;
    rom[7841] = 25'b1111111111111011011001110;
    rom[7842] = 25'b1111111111111011011010110;
    rom[7843] = 25'b1111111111111011011011110;
    rom[7844] = 25'b1111111111111011011100110;
    rom[7845] = 25'b1111111111111011011101110;
    rom[7846] = 25'b1111111111111011011110110;
    rom[7847] = 25'b1111111111111011011111111;
    rom[7848] = 25'b1111111111111011100000111;
    rom[7849] = 25'b1111111111111011100001111;
    rom[7850] = 25'b1111111111111011100010111;
    rom[7851] = 25'b1111111111111011100100000;
    rom[7852] = 25'b1111111111111011100101000;
    rom[7853] = 25'b1111111111111011100110000;
    rom[7854] = 25'b1111111111111011100111000;
    rom[7855] = 25'b1111111111111011101000000;
    rom[7856] = 25'b1111111111111011101001001;
    rom[7857] = 25'b1111111111111011101010001;
    rom[7858] = 25'b1111111111111011101011001;
    rom[7859] = 25'b1111111111111011101100001;
    rom[7860] = 25'b1111111111111011101101010;
    rom[7861] = 25'b1111111111111011101110010;
    rom[7862] = 25'b1111111111111011101111010;
    rom[7863] = 25'b1111111111111011110000010;
    rom[7864] = 25'b1111111111111011110001011;
    rom[7865] = 25'b1111111111111011110010011;
    rom[7866] = 25'b1111111111111011110011100;
    rom[7867] = 25'b1111111111111011110100100;
    rom[7868] = 25'b1111111111111011110101100;
    rom[7869] = 25'b1111111111111011110110100;
    rom[7870] = 25'b1111111111111011110111101;
    rom[7871] = 25'b1111111111111011111000101;
    rom[7872] = 25'b1111111111111011111001110;
    rom[7873] = 25'b1111111111111011111010110;
    rom[7874] = 25'b1111111111111011111011111;
    rom[7875] = 25'b1111111111111011111100111;
    rom[7876] = 25'b1111111111111011111101111;
    rom[7877] = 25'b1111111111111011111110111;
    rom[7878] = 25'b1111111111111100000000000;
    rom[7879] = 25'b1111111111111100000001001;
    rom[7880] = 25'b1111111111111100000010001;
    rom[7881] = 25'b1111111111111100000011010;
    rom[7882] = 25'b1111111111111100000100010;
    rom[7883] = 25'b1111111111111100000101010;
    rom[7884] = 25'b1111111111111100000110011;
    rom[7885] = 25'b1111111111111100000111011;
    rom[7886] = 25'b1111111111111100001000100;
    rom[7887] = 25'b1111111111111100001001101;
    rom[7888] = 25'b1111111111111100001010101;
    rom[7889] = 25'b1111111111111100001011110;
    rom[7890] = 25'b1111111111111100001100110;
    rom[7891] = 25'b1111111111111100001101111;
    rom[7892] = 25'b1111111111111100001110111;
    rom[7893] = 25'b1111111111111100010000000;
    rom[7894] = 25'b1111111111111100010001000;
    rom[7895] = 25'b1111111111111100010010001;
    rom[7896] = 25'b1111111111111100010011010;
    rom[7897] = 25'b1111111111111100010100011;
    rom[7898] = 25'b1111111111111100010101011;
    rom[7899] = 25'b1111111111111100010110100;
    rom[7900] = 25'b1111111111111100010111100;
    rom[7901] = 25'b1111111111111100011000101;
    rom[7902] = 25'b1111111111111100011001101;
    rom[7903] = 25'b1111111111111100011010110;
    rom[7904] = 25'b1111111111111100011011111;
    rom[7905] = 25'b1111111111111100011100111;
    rom[7906] = 25'b1111111111111100011110000;
    rom[7907] = 25'b1111111111111100011111001;
    rom[7908] = 25'b1111111111111100100000001;
    rom[7909] = 25'b1111111111111100100001010;
    rom[7910] = 25'b1111111111111100100010011;
    rom[7911] = 25'b1111111111111100100011100;
    rom[7912] = 25'b1111111111111100100100101;
    rom[7913] = 25'b1111111111111100100101110;
    rom[7914] = 25'b1111111111111100100110110;
    rom[7915] = 25'b1111111111111100100111111;
    rom[7916] = 25'b1111111111111100101001000;
    rom[7917] = 25'b1111111111111100101010001;
    rom[7918] = 25'b1111111111111100101011001;
    rom[7919] = 25'b1111111111111100101100010;
    rom[7920] = 25'b1111111111111100101101011;
    rom[7921] = 25'b1111111111111100101110100;
    rom[7922] = 25'b1111111111111100101111101;
    rom[7923] = 25'b1111111111111100110000110;
    rom[7924] = 25'b1111111111111100110001110;
    rom[7925] = 25'b1111111111111100110010111;
    rom[7926] = 25'b1111111111111100110100000;
    rom[7927] = 25'b1111111111111100110101001;
    rom[7928] = 25'b1111111111111100110110010;
    rom[7929] = 25'b1111111111111100110111011;
    rom[7930] = 25'b1111111111111100111000100;
    rom[7931] = 25'b1111111111111100111001101;
    rom[7932] = 25'b1111111111111100111010110;
    rom[7933] = 25'b1111111111111100111011111;
    rom[7934] = 25'b1111111111111100111101000;
    rom[7935] = 25'b1111111111111100111110000;
    rom[7936] = 25'b1111111111111100111111001;
    rom[7937] = 25'b1111111111111101000000010;
    rom[7938] = 25'b1111111111111101000001011;
    rom[7939] = 25'b1111111111111101000010100;
    rom[7940] = 25'b1111111111111101000011101;
    rom[7941] = 25'b1111111111111101000100110;
    rom[7942] = 25'b1111111111111101000101111;
    rom[7943] = 25'b1111111111111101000111000;
    rom[7944] = 25'b1111111111111101001000001;
    rom[7945] = 25'b1111111111111101001001010;
    rom[7946] = 25'b1111111111111101001010011;
    rom[7947] = 25'b1111111111111101001011100;
    rom[7948] = 25'b1111111111111101001100101;
    rom[7949] = 25'b1111111111111101001101110;
    rom[7950] = 25'b1111111111111101001111000;
    rom[7951] = 25'b1111111111111101010000001;
    rom[7952] = 25'b1111111111111101010001010;
    rom[7953] = 25'b1111111111111101010010011;
    rom[7954] = 25'b1111111111111101010011100;
    rom[7955] = 25'b1111111111111101010100101;
    rom[7956] = 25'b1111111111111101010101110;
    rom[7957] = 25'b1111111111111101010110111;
    rom[7958] = 25'b1111111111111101011000000;
    rom[7959] = 25'b1111111111111101011001001;
    rom[7960] = 25'b1111111111111101011010011;
    rom[7961] = 25'b1111111111111101011011100;
    rom[7962] = 25'b1111111111111101011100101;
    rom[7963] = 25'b1111111111111101011101111;
    rom[7964] = 25'b1111111111111101011111000;
    rom[7965] = 25'b1111111111111101100000000;
    rom[7966] = 25'b1111111111111101100001001;
    rom[7967] = 25'b1111111111111101100010011;
    rom[7968] = 25'b1111111111111101100011100;
    rom[7969] = 25'b1111111111111101100100110;
    rom[7970] = 25'b1111111111111101100101111;
    rom[7971] = 25'b1111111111111101100111000;
    rom[7972] = 25'b1111111111111101101000001;
    rom[7973] = 25'b1111111111111101101001010;
    rom[7974] = 25'b1111111111111101101010100;
    rom[7975] = 25'b1111111111111101101011101;
    rom[7976] = 25'b1111111111111101101100110;
    rom[7977] = 25'b1111111111111101101110000;
    rom[7978] = 25'b1111111111111101101111001;
    rom[7979] = 25'b1111111111111101110000010;
    rom[7980] = 25'b1111111111111101110001011;
    rom[7981] = 25'b1111111111111101110010101;
    rom[7982] = 25'b1111111111111101110011110;
    rom[7983] = 25'b1111111111111101110101000;
    rom[7984] = 25'b1111111111111101110110001;
    rom[7985] = 25'b1111111111111101110111010;
    rom[7986] = 25'b1111111111111101111000100;
    rom[7987] = 25'b1111111111111101111001101;
    rom[7988] = 25'b1111111111111101111010111;
    rom[7989] = 25'b1111111111111101111100000;
    rom[7990] = 25'b1111111111111101111101010;
    rom[7991] = 25'b1111111111111101111110011;
    rom[7992] = 25'b1111111111111101111111100;
    rom[7993] = 25'b1111111111111110000000110;
    rom[7994] = 25'b1111111111111110000001111;
    rom[7995] = 25'b1111111111111110000011001;
    rom[7996] = 25'b1111111111111110000100010;
    rom[7997] = 25'b1111111111111110000101011;
    rom[7998] = 25'b1111111111111110000110101;
    rom[7999] = 25'b1111111111111110000111111;
    rom[8000] = 25'b1111111111111110001001000;
    rom[8001] = 25'b1111111111111110001010001;
    rom[8002] = 25'b1111111111111110001011011;
    rom[8003] = 25'b1111111111111110001100101;
    rom[8004] = 25'b1111111111111110001101110;
    rom[8005] = 25'b1111111111111110001111000;
    rom[8006] = 25'b1111111111111110010000001;
    rom[8007] = 25'b1111111111111110010001011;
    rom[8008] = 25'b1111111111111110010010101;
    rom[8009] = 25'b1111111111111110010011110;
    rom[8010] = 25'b1111111111111110010100111;
    rom[8011] = 25'b1111111111111110010110001;
    rom[8012] = 25'b1111111111111110010111011;
    rom[8013] = 25'b1111111111111110011000100;
    rom[8014] = 25'b1111111111111110011001110;
    rom[8015] = 25'b1111111111111110011010111;
    rom[8016] = 25'b1111111111111110011100001;
    rom[8017] = 25'b1111111111111110011101011;
    rom[8018] = 25'b1111111111111110011110100;
    rom[8019] = 25'b1111111111111110011111110;
    rom[8020] = 25'b1111111111111110100001000;
    rom[8021] = 25'b1111111111111110100010001;
    rom[8022] = 25'b1111111111111110100011011;
    rom[8023] = 25'b1111111111111110100100101;
    rom[8024] = 25'b1111111111111110100101111;
    rom[8025] = 25'b1111111111111110100111000;
    rom[8026] = 25'b1111111111111110101000010;
    rom[8027] = 25'b1111111111111110101001100;
    rom[8028] = 25'b1111111111111110101010101;
    rom[8029] = 25'b1111111111111110101011111;
    rom[8030] = 25'b1111111111111110101101001;
    rom[8031] = 25'b1111111111111110101110011;
    rom[8032] = 25'b1111111111111110101111100;
    rom[8033] = 25'b1111111111111110110000110;
    rom[8034] = 25'b1111111111111110110010000;
    rom[8035] = 25'b1111111111111110110011001;
    rom[8036] = 25'b1111111111111110110100011;
    rom[8037] = 25'b1111111111111110110101101;
    rom[8038] = 25'b1111111111111110110110111;
    rom[8039] = 25'b1111111111111110111000001;
    rom[8040] = 25'b1111111111111110111001011;
    rom[8041] = 25'b1111111111111110111010100;
    rom[8042] = 25'b1111111111111110111011110;
    rom[8043] = 25'b1111111111111110111101000;
    rom[8044] = 25'b1111111111111110111110010;
    rom[8045] = 25'b1111111111111110111111100;
    rom[8046] = 25'b1111111111111111000000110;
    rom[8047] = 25'b1111111111111111000001111;
    rom[8048] = 25'b1111111111111111000011001;
    rom[8049] = 25'b1111111111111111000100100;
    rom[8050] = 25'b1111111111111111000101101;
    rom[8051] = 25'b1111111111111111000110111;
    rom[8052] = 25'b1111111111111111001000001;
    rom[8053] = 25'b1111111111111111001001011;
    rom[8054] = 25'b1111111111111111001010101;
    rom[8055] = 25'b1111111111111111001011111;
    rom[8056] = 25'b1111111111111111001101001;
    rom[8057] = 25'b1111111111111111001110011;
    rom[8058] = 25'b1111111111111111001111101;
    rom[8059] = 25'b1111111111111111010000111;
    rom[8060] = 25'b1111111111111111010010001;
    rom[8061] = 25'b1111111111111111010011010;
    rom[8062] = 25'b1111111111111111010100101;
    rom[8063] = 25'b1111111111111111010101111;
    rom[8064] = 25'b1111111111111111010111000;
    rom[8065] = 25'b1111111111111111011000011;
    rom[8066] = 25'b1111111111111111011001100;
    rom[8067] = 25'b1111111111111111011010111;
    rom[8068] = 25'b1111111111111111011100001;
    rom[8069] = 25'b1111111111111111011101011;
    rom[8070] = 25'b1111111111111111011110101;
    rom[8071] = 25'b1111111111111111011111110;
    rom[8072] = 25'b1111111111111111100001001;
    rom[8073] = 25'b1111111111111111100010011;
    rom[8074] = 25'b1111111111111111100011101;
    rom[8075] = 25'b1111111111111111100100111;
    rom[8076] = 25'b1111111111111111100110001;
    rom[8077] = 25'b1111111111111111100111011;
    rom[8078] = 25'b1111111111111111101000101;
    rom[8079] = 25'b1111111111111111101010000;
    rom[8080] = 25'b1111111111111111101011010;
    rom[8081] = 25'b1111111111111111101100100;
    rom[8082] = 25'b1111111111111111101101110;
    rom[8083] = 25'b1111111111111111101111000;
    rom[8084] = 25'b1111111111111111110000010;
    rom[8085] = 25'b1111111111111111110001100;
    rom[8086] = 25'b1111111111111111110010111;
    rom[8087] = 25'b1111111111111111110100001;
    rom[8088] = 25'b1111111111111111110101011;
    rom[8089] = 25'b1111111111111111110110110;
    rom[8090] = 25'b1111111111111111110111111;
    rom[8091] = 25'b1111111111111111111001010;
    rom[8092] = 25'b1111111111111111111010011;
    rom[8093] = 25'b1111111111111111111011110;
    rom[8094] = 25'b1111111111111111111101000;
    rom[8095] = 25'b1111111111111111111110011;
    rom[8096] = 25'b1111111111111111111111101;
    rom[8097] = 25'b0000000000000000000000110;
    rom[8098] = 25'b0000000000000000000010001;
    rom[8099] = 25'b0000000000000000000011010;
    rom[8100] = 25'b0000000000000000000100101;
    rom[8101] = 25'b0000000000000000000101111;
    rom[8102] = 25'b0000000000000000000111010;
    rom[8103] = 25'b0000000000000000001000100;
    rom[8104] = 25'b0000000000000000001001110;
    rom[8105] = 25'b0000000000000000001011000;
    rom[8106] = 25'b0000000000000000001100011;
    rom[8107] = 25'b0000000000000000001101101;
    rom[8108] = 25'b0000000000000000001111000;
    rom[8109] = 25'b0000000000000000010000001;
    rom[8110] = 25'b0000000000000000010001100;
    rom[8111] = 25'b0000000000000000010010110;
    rom[8112] = 25'b0000000000000000010100001;
    rom[8113] = 25'b0000000000000000010101011;
    rom[8114] = 25'b0000000000000000010110110;
    rom[8115] = 25'b0000000000000000011000000;
    rom[8116] = 25'b0000000000000000011001011;
    rom[8117] = 25'b0000000000000000011010101;
    rom[8118] = 25'b0000000000000000011011111;
    rom[8119] = 25'b0000000000000000011101001;
    rom[8120] = 25'b0000000000000000011110100;
    rom[8121] = 25'b0000000000000000011111110;
    rom[8122] = 25'b0000000000000000100001001;
    rom[8123] = 25'b0000000000000000100010011;
    rom[8124] = 25'b0000000000000000100011110;
    rom[8125] = 25'b0000000000000000100101000;
    rom[8126] = 25'b0000000000000000100110011;
    rom[8127] = 25'b0000000000000000100111101;
    rom[8128] = 25'b0000000000000000101000111;
    rom[8129] = 25'b0000000000000000101010010;
    rom[8130] = 25'b0000000000000000101011100;
    rom[8131] = 25'b0000000000000000101100111;
    rom[8132] = 25'b0000000000000000101110001;
    rom[8133] = 25'b0000000000000000101111100;
    rom[8134] = 25'b0000000000000000110000111;
    rom[8135] = 25'b0000000000000000110010001;
    rom[8136] = 25'b0000000000000000110011100;
    rom[8137] = 25'b0000000000000000110100110;
    rom[8138] = 25'b0000000000000000110110001;
    rom[8139] = 25'b0000000000000000110111011;
    rom[8140] = 25'b0000000000000000111000110;
    rom[8141] = 25'b0000000000000000111010000;
    rom[8142] = 25'b0000000000000000111011011;
    rom[8143] = 25'b0000000000000000111100110;
    rom[8144] = 25'b0000000000000000111110000;
    rom[8145] = 25'b0000000000000000111111011;
    rom[8146] = 25'b0000000000000001000000101;
    rom[8147] = 25'b0000000000000001000010000;
    rom[8148] = 25'b0000000000000001000011011;
    rom[8149] = 25'b0000000000000001000100101;
    rom[8150] = 25'b0000000000000001000110000;
    rom[8151] = 25'b0000000000000001000111010;
    rom[8152] = 25'b0000000000000001001000101;
    rom[8153] = 25'b0000000000000001001010000;
    rom[8154] = 25'b0000000000000001001011010;
    rom[8155] = 25'b0000000000000001001100101;
    rom[8156] = 25'b0000000000000001001110000;
    rom[8157] = 25'b0000000000000001001111011;
    rom[8158] = 25'b0000000000000001010000101;
    rom[8159] = 25'b0000000000000001010001111;
    rom[8160] = 25'b0000000000000001010011011;
    rom[8161] = 25'b0000000000000001010100101;
    rom[8162] = 25'b0000000000000001010110000;
    rom[8163] = 25'b0000000000000001010111011;
    rom[8164] = 25'b0000000000000001011000101;
    rom[8165] = 25'b0000000000000001011010000;
    rom[8166] = 25'b0000000000000001011011011;
    rom[8167] = 25'b0000000000000001011100101;
    rom[8168] = 25'b0000000000000001011110001;
    rom[8169] = 25'b0000000000000001011111011;
    rom[8170] = 25'b0000000000000001100000101;
    rom[8171] = 25'b0000000000000001100010001;
    rom[8172] = 25'b0000000000000001100011011;
    rom[8173] = 25'b0000000000000001100100110;
    rom[8174] = 25'b0000000000000001100110001;
    rom[8175] = 25'b0000000000000001100111011;
    rom[8176] = 25'b0000000000000001101000110;
    rom[8177] = 25'b0000000000000001101010001;
    rom[8178] = 25'b0000000000000001101011100;
    rom[8179] = 25'b0000000000000001101100111;
    rom[8180] = 25'b0000000000000001101110010;
    rom[8181] = 25'b0000000000000001101111100;
    rom[8182] = 25'b0000000000000001110000111;
    rom[8183] = 25'b0000000000000001110010010;
    rom[8184] = 25'b0000000000000001110011101;
    rom[8185] = 25'b0000000000000001110101000;
    rom[8186] = 25'b0000000000000001110110011;
    rom[8187] = 25'b0000000000000001110111110;
    rom[8188] = 25'b0000000000000001111001000;
    rom[8189] = 25'b0000000000000001111010100;
    rom[8190] = 25'b0000000000000001111011110;
    rom[8191] = 25'b0000000000000001111101001;
    rom[8192] = 25'b0000000000000001111110100;
    rom[8193] = 25'b0000000000000001111111111;
    rom[8194] = 25'b0000000000000010000001010;
    rom[8195] = 25'b0000000000000010000010101;
    rom[8196] = 25'b0000000000000010000100000;
    rom[8197] = 25'b0000000000000010000101010;
    rom[8198] = 25'b0000000000000010000110110;
    rom[8199] = 25'b0000000000000010001000001;
    rom[8200] = 25'b0000000000000010001001011;
    rom[8201] = 25'b0000000000000010001010110;
    rom[8202] = 25'b0000000000000010001100010;
    rom[8203] = 25'b0000000000000010001101100;
    rom[8204] = 25'b0000000000000010001110111;
    rom[8205] = 25'b0000000000000010010000011;
    rom[8206] = 25'b0000000000000010010001110;
    rom[8207] = 25'b0000000000000010010011000;
    rom[8208] = 25'b0000000000000010010100011;
    rom[8209] = 25'b0000000000000010010101111;
    rom[8210] = 25'b0000000000000010010111001;
    rom[8211] = 25'b0000000000000010011000100;
    rom[8212] = 25'b0000000000000010011001111;
    rom[8213] = 25'b0000000000000010011011011;
    rom[8214] = 25'b0000000000000010011100101;
    rom[8215] = 25'b0000000000000010011110000;
    rom[8216] = 25'b0000000000000010011111100;
    rom[8217] = 25'b0000000000000010100000111;
    rom[8218] = 25'b0000000000000010100010010;
    rom[8219] = 25'b0000000000000010100011100;
    rom[8220] = 25'b0000000000000010100101000;
    rom[8221] = 25'b0000000000000010100110011;
    rom[8222] = 25'b0000000000000010100111110;
    rom[8223] = 25'b0000000000000010101001001;
    rom[8224] = 25'b0000000000000010101010100;
    rom[8225] = 25'b0000000000000010101100000;
    rom[8226] = 25'b0000000000000010101101010;
    rom[8227] = 25'b0000000000000010101110101;
    rom[8228] = 25'b0000000000000010110000001;
    rom[8229] = 25'b0000000000000010110001100;
    rom[8230] = 25'b0000000000000010110010111;
    rom[8231] = 25'b0000000000000010110100010;
    rom[8232] = 25'b0000000000000010110101101;
    rom[8233] = 25'b0000000000000010110111001;
    rom[8234] = 25'b0000000000000010111000100;
    rom[8235] = 25'b0000000000000010111001111;
    rom[8236] = 25'b0000000000000010111011010;
    rom[8237] = 25'b0000000000000010111100101;
    rom[8238] = 25'b0000000000000010111110000;
    rom[8239] = 25'b0000000000000010111111011;
    rom[8240] = 25'b0000000000000011000000110;
    rom[8241] = 25'b0000000000000011000010001;
    rom[8242] = 25'b0000000000000011000011101;
    rom[8243] = 25'b0000000000000011000101000;
    rom[8244] = 25'b0000000000000011000110011;
    rom[8245] = 25'b0000000000000011000111110;
    rom[8246] = 25'b0000000000000011001001001;
    rom[8247] = 25'b0000000000000011001010101;
    rom[8248] = 25'b0000000000000011001100000;
    rom[8249] = 25'b0000000000000011001101100;
    rom[8250] = 25'b0000000000000011001110111;
    rom[8251] = 25'b0000000000000011010000010;
    rom[8252] = 25'b0000000000000011010001101;
    rom[8253] = 25'b0000000000000011010011001;
    rom[8254] = 25'b0000000000000011010100100;
    rom[8255] = 25'b0000000000000011010101111;
    rom[8256] = 25'b0000000000000011010111010;
    rom[8257] = 25'b0000000000000011011000110;
    rom[8258] = 25'b0000000000000011011010001;
    rom[8259] = 25'b0000000000000011011011100;
    rom[8260] = 25'b0000000000000011011101000;
    rom[8261] = 25'b0000000000000011011110011;
    rom[8262] = 25'b0000000000000011011111110;
    rom[8263] = 25'b0000000000000011100001001;
    rom[8264] = 25'b0000000000000011100010101;
    rom[8265] = 25'b0000000000000011100100000;
    rom[8266] = 25'b0000000000000011100101011;
    rom[8267] = 25'b0000000000000011100110111;
    rom[8268] = 25'b0000000000000011101000010;
    rom[8269] = 25'b0000000000000011101001101;
    rom[8270] = 25'b0000000000000011101011001;
    rom[8271] = 25'b0000000000000011101100100;
    rom[8272] = 25'b0000000000000011101110000;
    rom[8273] = 25'b0000000000000011101111011;
    rom[8274] = 25'b0000000000000011110000110;
    rom[8275] = 25'b0000000000000011110010001;
    rom[8276] = 25'b0000000000000011110011101;
    rom[8277] = 25'b0000000000000011110101001;
    rom[8278] = 25'b0000000000000011110110100;
    rom[8279] = 25'b0000000000000011110111111;
    rom[8280] = 25'b0000000000000011111001011;
    rom[8281] = 25'b0000000000000011111010110;
    rom[8282] = 25'b0000000000000011111100001;
    rom[8283] = 25'b0000000000000011111101101;
    rom[8284] = 25'b0000000000000011111111001;
    rom[8285] = 25'b0000000000000100000000100;
    rom[8286] = 25'b0000000000000100000001111;
    rom[8287] = 25'b0000000000000100000011011;
    rom[8288] = 25'b0000000000000100000100110;
    rom[8289] = 25'b0000000000000100000110001;
    rom[8290] = 25'b0000000000000100000111101;
    rom[8291] = 25'b0000000000000100001001001;
    rom[8292] = 25'b0000000000000100001010100;
    rom[8293] = 25'b0000000000000100001100000;
    rom[8294] = 25'b0000000000000100001101011;
    rom[8295] = 25'b0000000000000100001110111;
    rom[8296] = 25'b0000000000000100010000010;
    rom[8297] = 25'b0000000000000100010001101;
    rom[8298] = 25'b0000000000000100010011001;
    rom[8299] = 25'b0000000000000100010100100;
    rom[8300] = 25'b0000000000000100010110000;
    rom[8301] = 25'b0000000000000100010111100;
    rom[8302] = 25'b0000000000000100011000111;
    rom[8303] = 25'b0000000000000100011010011;
    rom[8304] = 25'b0000000000000100011011110;
    rom[8305] = 25'b0000000000000100011101010;
    rom[8306] = 25'b0000000000000100011110101;
    rom[8307] = 25'b0000000000000100100000001;
    rom[8308] = 25'b0000000000000100100001100;
    rom[8309] = 25'b0000000000000100100010111;
    rom[8310] = 25'b0000000000000100100100011;
    rom[8311] = 25'b0000000000000100100101111;
    rom[8312] = 25'b0000000000000100100111011;
    rom[8313] = 25'b0000000000000100101000110;
    rom[8314] = 25'b0000000000000100101010010;
    rom[8315] = 25'b0000000000000100101011101;
    rom[8316] = 25'b0000000000000100101101001;
    rom[8317] = 25'b0000000000000100101110100;
    rom[8318] = 25'b0000000000000100110000000;
    rom[8319] = 25'b0000000000000100110001011;
    rom[8320] = 25'b0000000000000100110010111;
    rom[8321] = 25'b0000000000000100110100011;
    rom[8322] = 25'b0000000000000100110101110;
    rom[8323] = 25'b0000000000000100110111010;
    rom[8324] = 25'b0000000000000100111000110;
    rom[8325] = 25'b0000000000000100111010001;
    rom[8326] = 25'b0000000000000100111011101;
    rom[8327] = 25'b0000000000000100111101001;
    rom[8328] = 25'b0000000000000100111110101;
    rom[8329] = 25'b0000000000000101000000000;
    rom[8330] = 25'b0000000000000101000001100;
    rom[8331] = 25'b0000000000000101000010111;
    rom[8332] = 25'b0000000000000101000100011;
    rom[8333] = 25'b0000000000000101000101111;
    rom[8334] = 25'b0000000000000101000111010;
    rom[8335] = 25'b0000000000000101001000110;
    rom[8336] = 25'b0000000000000101001010001;
    rom[8337] = 25'b0000000000000101001011101;
    rom[8338] = 25'b0000000000000101001101001;
    rom[8339] = 25'b0000000000000101001110100;
    rom[8340] = 25'b0000000000000101010000000;
    rom[8341] = 25'b0000000000000101010001100;
    rom[8342] = 25'b0000000000000101010010111;
    rom[8343] = 25'b0000000000000101010100011;
    rom[8344] = 25'b0000000000000101010101111;
    rom[8345] = 25'b0000000000000101010111011;
    rom[8346] = 25'b0000000000000101011000111;
    rom[8347] = 25'b0000000000000101011010010;
    rom[8348] = 25'b0000000000000101011011110;
    rom[8349] = 25'b0000000000000101011101010;
    rom[8350] = 25'b0000000000000101011110110;
    rom[8351] = 25'b0000000000000101100000010;
    rom[8352] = 25'b0000000000000101100001101;
    rom[8353] = 25'b0000000000000101100011001;
    rom[8354] = 25'b0000000000000101100100101;
    rom[8355] = 25'b0000000000000101100110001;
    rom[8356] = 25'b0000000000000101100111100;
    rom[8357] = 25'b0000000000000101101001000;
    rom[8358] = 25'b0000000000000101101010100;
    rom[8359] = 25'b0000000000000101101100000;
    rom[8360] = 25'b0000000000000101101101011;
    rom[8361] = 25'b0000000000000101101110111;
    rom[8362] = 25'b0000000000000101110000011;
    rom[8363] = 25'b0000000000000101110001111;
    rom[8364] = 25'b0000000000000101110011011;
    rom[8365] = 25'b0000000000000101110100110;
    rom[8366] = 25'b0000000000000101110110010;
    rom[8367] = 25'b0000000000000101110111110;
    rom[8368] = 25'b0000000000000101111001010;
    rom[8369] = 25'b0000000000000101111010110;
    rom[8370] = 25'b0000000000000101111100001;
    rom[8371] = 25'b0000000000000101111101101;
    rom[8372] = 25'b0000000000000101111111001;
    rom[8373] = 25'b0000000000000110000000101;
    rom[8374] = 25'b0000000000000110000010001;
    rom[8375] = 25'b0000000000000110000011101;
    rom[8376] = 25'b0000000000000110000101001;
    rom[8377] = 25'b0000000000000110000110100;
    rom[8378] = 25'b0000000000000110001000000;
    rom[8379] = 25'b0000000000000110001001100;
    rom[8380] = 25'b0000000000000110001011000;
    rom[8381] = 25'b0000000000000110001100100;
    rom[8382] = 25'b0000000000000110001110000;
    rom[8383] = 25'b0000000000000110001111100;
    rom[8384] = 25'b0000000000000110010001000;
    rom[8385] = 25'b0000000000000110010010011;
    rom[8386] = 25'b0000000000000110010011111;
    rom[8387] = 25'b0000000000000110010101011;
    rom[8388] = 25'b0000000000000110010110111;
    rom[8389] = 25'b0000000000000110011000011;
    rom[8390] = 25'b0000000000000110011001111;
    rom[8391] = 25'b0000000000000110011011010;
    rom[8392] = 25'b0000000000000110011100110;
    rom[8393] = 25'b0000000000000110011110010;
    rom[8394] = 25'b0000000000000110011111110;
    rom[8395] = 25'b0000000000000110100001010;
    rom[8396] = 25'b0000000000000110100010110;
    rom[8397] = 25'b0000000000000110100100010;
    rom[8398] = 25'b0000000000000110100101110;
    rom[8399] = 25'b0000000000000110100111010;
    rom[8400] = 25'b0000000000000110101000110;
    rom[8401] = 25'b0000000000000110101010010;
    rom[8402] = 25'b0000000000000110101011110;
    rom[8403] = 25'b0000000000000110101101010;
    rom[8404] = 25'b0000000000000110101110110;
    rom[8405] = 25'b0000000000000110110000010;
    rom[8406] = 25'b0000000000000110110001110;
    rom[8407] = 25'b0000000000000110110011010;
    rom[8408] = 25'b0000000000000110110100110;
    rom[8409] = 25'b0000000000000110110110010;
    rom[8410] = 25'b0000000000000110110111110;
    rom[8411] = 25'b0000000000000110111001010;
    rom[8412] = 25'b0000000000000110111010101;
    rom[8413] = 25'b0000000000000110111100001;
    rom[8414] = 25'b0000000000000110111101101;
    rom[8415] = 25'b0000000000000110111111001;
    rom[8416] = 25'b0000000000000111000000101;
    rom[8417] = 25'b0000000000000111000010001;
    rom[8418] = 25'b0000000000000111000011101;
    rom[8419] = 25'b0000000000000111000101001;
    rom[8420] = 25'b0000000000000111000110101;
    rom[8421] = 25'b0000000000000111001000001;
    rom[8422] = 25'b0000000000000111001001101;
    rom[8423] = 25'b0000000000000111001011001;
    rom[8424] = 25'b0000000000000111001100101;
    rom[8425] = 25'b0000000000000111001110010;
    rom[8426] = 25'b0000000000000111001111110;
    rom[8427] = 25'b0000000000000111010001010;
    rom[8428] = 25'b0000000000000111010010101;
    rom[8429] = 25'b0000000000000111010100001;
    rom[8430] = 25'b0000000000000111010101101;
    rom[8431] = 25'b0000000000000111010111001;
    rom[8432] = 25'b0000000000000111011000101;
    rom[8433] = 25'b0000000000000111011010001;
    rom[8434] = 25'b0000000000000111011011110;
    rom[8435] = 25'b0000000000000111011101010;
    rom[8436] = 25'b0000000000000111011110110;
    rom[8437] = 25'b0000000000000111100000010;
    rom[8438] = 25'b0000000000000111100001110;
    rom[8439] = 25'b0000000000000111100011010;
    rom[8440] = 25'b0000000000000111100100110;
    rom[8441] = 25'b0000000000000111100110010;
    rom[8442] = 25'b0000000000000111100111110;
    rom[8443] = 25'b0000000000000111101001010;
    rom[8444] = 25'b0000000000000111101010110;
    rom[8445] = 25'b0000000000000111101100010;
    rom[8446] = 25'b0000000000000111101101110;
    rom[8447] = 25'b0000000000000111101111011;
    rom[8448] = 25'b0000000000000111110000111;
    rom[8449] = 25'b0000000000000111110010011;
    rom[8450] = 25'b0000000000000111110011111;
    rom[8451] = 25'b0000000000000111110101011;
    rom[8452] = 25'b0000000000000111110110111;
    rom[8453] = 25'b0000000000000111111000011;
    rom[8454] = 25'b0000000000000111111001111;
    rom[8455] = 25'b0000000000000111111011011;
    rom[8456] = 25'b0000000000000111111100111;
    rom[8457] = 25'b0000000000000111111110100;
    rom[8458] = 25'b0000000000001000000000000;
    rom[8459] = 25'b0000000000001000000001100;
    rom[8460] = 25'b0000000000001000000011000;
    rom[8461] = 25'b0000000000001000000100100;
    rom[8462] = 25'b0000000000001000000110000;
    rom[8463] = 25'b0000000000001000000111100;
    rom[8464] = 25'b0000000000001000001001000;
    rom[8465] = 25'b0000000000001000001010100;
    rom[8466] = 25'b0000000000001000001100001;
    rom[8467] = 25'b0000000000001000001101101;
    rom[8468] = 25'b0000000000001000001111001;
    rom[8469] = 25'b0000000000001000010000101;
    rom[8470] = 25'b0000000000001000010010010;
    rom[8471] = 25'b0000000000001000010011101;
    rom[8472] = 25'b0000000000001000010101001;
    rom[8473] = 25'b0000000000001000010110101;
    rom[8474] = 25'b0000000000001000011000010;
    rom[8475] = 25'b0000000000001000011001110;
    rom[8476] = 25'b0000000000001000011011010;
    rom[8477] = 25'b0000000000001000011100111;
    rom[8478] = 25'b0000000000001000011110011;
    rom[8479] = 25'b0000000000001000011111111;
    rom[8480] = 25'b0000000000001000100001011;
    rom[8481] = 25'b0000000000001000100010111;
    rom[8482] = 25'b0000000000001000100100011;
    rom[8483] = 25'b0000000000001000100101111;
    rom[8484] = 25'b0000000000001000100111100;
    rom[8485] = 25'b0000000000001000101001000;
    rom[8486] = 25'b0000000000001000101010100;
    rom[8487] = 25'b0000000000001000101100000;
    rom[8488] = 25'b0000000000001000101101100;
    rom[8489] = 25'b0000000000001000101111000;
    rom[8490] = 25'b0000000000001000110000100;
    rom[8491] = 25'b0000000000001000110010001;
    rom[8492] = 25'b0000000000001000110011101;
    rom[8493] = 25'b0000000000001000110101001;
    rom[8494] = 25'b0000000000001000110110110;
    rom[8495] = 25'b0000000000001000111000010;
    rom[8496] = 25'b0000000000001000111001110;
    rom[8497] = 25'b0000000000001000111011010;
    rom[8498] = 25'b0000000000001000111100110;
    rom[8499] = 25'b0000000000001000111110010;
    rom[8500] = 25'b0000000000001000111111111;
    rom[8501] = 25'b0000000000001001000001011;
    rom[8502] = 25'b0000000000001001000010111;
    rom[8503] = 25'b0000000000001001000100011;
    rom[8504] = 25'b0000000000001001000101111;
    rom[8505] = 25'b0000000000001001000111100;
    rom[8506] = 25'b0000000000001001001001000;
    rom[8507] = 25'b0000000000001001001010100;
    rom[8508] = 25'b0000000000001001001100001;
    rom[8509] = 25'b0000000000001001001101101;
    rom[8510] = 25'b0000000000001001001111001;
    rom[8511] = 25'b0000000000001001010000101;
    rom[8512] = 25'b0000000000001001010010001;
    rom[8513] = 25'b0000000000001001010011110;
    rom[8514] = 25'b0000000000001001010101010;
    rom[8515] = 25'b0000000000001001010110110;
    rom[8516] = 25'b0000000000001001011000011;
    rom[8517] = 25'b0000000000001001011001111;
    rom[8518] = 25'b0000000000001001011011010;
    rom[8519] = 25'b0000000000001001011100111;
    rom[8520] = 25'b0000000000001001011110011;
    rom[8521] = 25'b0000000000001001100000000;
    rom[8522] = 25'b0000000000001001100001100;
    rom[8523] = 25'b0000000000001001100011000;
    rom[8524] = 25'b0000000000001001100100100;
    rom[8525] = 25'b0000000000001001100110000;
    rom[8526] = 25'b0000000000001001100111101;
    rom[8527] = 25'b0000000000001001101001001;
    rom[8528] = 25'b0000000000001001101010101;
    rom[8529] = 25'b0000000000001001101100010;
    rom[8530] = 25'b0000000000001001101101110;
    rom[8531] = 25'b0000000000001001101111010;
    rom[8532] = 25'b0000000000001001110000110;
    rom[8533] = 25'b0000000000001001110010011;
    rom[8534] = 25'b0000000000001001110011111;
    rom[8535] = 25'b0000000000001001110101011;
    rom[8536] = 25'b0000000000001001110111000;
    rom[8537] = 25'b0000000000001001111000100;
    rom[8538] = 25'b0000000000001001111010000;
    rom[8539] = 25'b0000000000001001111011100;
    rom[8540] = 25'b0000000000001001111101001;
    rom[8541] = 25'b0000000000001001111110101;
    rom[8542] = 25'b0000000000001010000000001;
    rom[8543] = 25'b0000000000001010000001110;
    rom[8544] = 25'b0000000000001010000011001;
    rom[8545] = 25'b0000000000001010000100110;
    rom[8546] = 25'b0000000000001010000110010;
    rom[8547] = 25'b0000000000001010000111111;
    rom[8548] = 25'b0000000000001010001001011;
    rom[8549] = 25'b0000000000001010001011000;
    rom[8550] = 25'b0000000000001010001100011;
    rom[8551] = 25'b0000000000001010001101111;
    rom[8552] = 25'b0000000000001010001111100;
    rom[8553] = 25'b0000000000001010010001000;
    rom[8554] = 25'b0000000000001010010010101;
    rom[8555] = 25'b0000000000001010010100001;
    rom[8556] = 25'b0000000000001010010101101;
    rom[8557] = 25'b0000000000001010010111001;
    rom[8558] = 25'b0000000000001010011000110;
    rom[8559] = 25'b0000000000001010011010010;
    rom[8560] = 25'b0000000000001010011011111;
    rom[8561] = 25'b0000000000001010011101011;
    rom[8562] = 25'b0000000000001010011110111;
    rom[8563] = 25'b0000000000001010100000011;
    rom[8564] = 25'b0000000000001010100001111;
    rom[8565] = 25'b0000000000001010100011100;
    rom[8566] = 25'b0000000000001010100101000;
    rom[8567] = 25'b0000000000001010100110101;
    rom[8568] = 25'b0000000000001010101000001;
    rom[8569] = 25'b0000000000001010101001101;
    rom[8570] = 25'b0000000000001010101011001;
    rom[8571] = 25'b0000000000001010101100110;
    rom[8572] = 25'b0000000000001010101110010;
    rom[8573] = 25'b0000000000001010101111111;
    rom[8574] = 25'b0000000000001010110001011;
    rom[8575] = 25'b0000000000001010110010111;
    rom[8576] = 25'b0000000000001010110100011;
    rom[8577] = 25'b0000000000001010110110000;
    rom[8578] = 25'b0000000000001010110111100;
    rom[8579] = 25'b0000000000001010111001001;
    rom[8580] = 25'b0000000000001010111010101;
    rom[8581] = 25'b0000000000001010111100000;
    rom[8582] = 25'b0000000000001010111101101;
    rom[8583] = 25'b0000000000001010111111001;
    rom[8584] = 25'b0000000000001011000000110;
    rom[8585] = 25'b0000000000001011000010010;
    rom[8586] = 25'b0000000000001011000011110;
    rom[8587] = 25'b0000000000001011000101010;
    rom[8588] = 25'b0000000000001011000110111;
    rom[8589] = 25'b0000000000001011001000011;
    rom[8590] = 25'b0000000000001011001010000;
    rom[8591] = 25'b0000000000001011001011100;
    rom[8592] = 25'b0000000000001011001101000;
    rom[8593] = 25'b0000000000001011001110100;
    rom[8594] = 25'b0000000000001011010000001;
    rom[8595] = 25'b0000000000001011010001101;
    rom[8596] = 25'b0000000000001011010011010;
    rom[8597] = 25'b0000000000001011010100110;
    rom[8598] = 25'b0000000000001011010110010;
    rom[8599] = 25'b0000000000001011010111110;
    rom[8600] = 25'b0000000000001011011001011;
    rom[8601] = 25'b0000000000001011011010111;
    rom[8602] = 25'b0000000000001011011100100;
    rom[8603] = 25'b0000000000001011011110000;
    rom[8604] = 25'b0000000000001011011111100;
    rom[8605] = 25'b0000000000001011100001000;
    rom[8606] = 25'b0000000000001011100010101;
    rom[8607] = 25'b0000000000001011100100001;
    rom[8608] = 25'b0000000000001011100101110;
    rom[8609] = 25'b0000000000001011100111010;
    rom[8610] = 25'b0000000000001011101000110;
    rom[8611] = 25'b0000000000001011101010010;
    rom[8612] = 25'b0000000000001011101011111;
    rom[8613] = 25'b0000000000001011101101011;
    rom[8614] = 25'b0000000000001011101111000;
    rom[8615] = 25'b0000000000001011110000100;
    rom[8616] = 25'b0000000000001011110010000;
    rom[8617] = 25'b0000000000001011110011100;
    rom[8618] = 25'b0000000000001011110101001;
    rom[8619] = 25'b0000000000001011110110101;
    rom[8620] = 25'b0000000000001011111000010;
    rom[8621] = 25'b0000000000001011111001110;
    rom[8622] = 25'b0000000000001011111011010;
    rom[8623] = 25'b0000000000001011111100110;
    rom[8624] = 25'b0000000000001011111110011;
    rom[8625] = 25'b0000000000001011111111111;
    rom[8626] = 25'b0000000000001100000001100;
    rom[8627] = 25'b0000000000001100000011000;
    rom[8628] = 25'b0000000000001100000100100;
    rom[8629] = 25'b0000000000001100000110000;
    rom[8630] = 25'b0000000000001100000111101;
    rom[8631] = 25'b0000000000001100001001001;
    rom[8632] = 25'b0000000000001100001010110;
    rom[8633] = 25'b0000000000001100001100001;
    rom[8634] = 25'b0000000000001100001101110;
    rom[8635] = 25'b0000000000001100001111010;
    rom[8636] = 25'b0000000000001100010000111;
    rom[8637] = 25'b0000000000001100010010011;
    rom[8638] = 25'b0000000000001100010011111;
    rom[8639] = 25'b0000000000001100010101011;
    rom[8640] = 25'b0000000000001100010110111;
    rom[8641] = 25'b0000000000001100011000100;
    rom[8642] = 25'b0000000000001100011010000;
    rom[8643] = 25'b0000000000001100011011101;
    rom[8644] = 25'b0000000000001100011101001;
    rom[8645] = 25'b0000000000001100011110101;
    rom[8646] = 25'b0000000000001100100000001;
    rom[8647] = 25'b0000000000001100100001110;
    rom[8648] = 25'b0000000000001100100011010;
    rom[8649] = 25'b0000000000001100100100111;
    rom[8650] = 25'b0000000000001100100110011;
    rom[8651] = 25'b0000000000001100100111111;
    rom[8652] = 25'b0000000000001100101001011;
    rom[8653] = 25'b0000000000001100101011000;
    rom[8654] = 25'b0000000000001100101100100;
    rom[8655] = 25'b0000000000001100101110001;
    rom[8656] = 25'b0000000000001100101111101;
    rom[8657] = 25'b0000000000001100110001001;
    rom[8658] = 25'b0000000000001100110010101;
    rom[8659] = 25'b0000000000001100110100010;
    rom[8660] = 25'b0000000000001100110101110;
    rom[8661] = 25'b0000000000001100110111011;
    rom[8662] = 25'b0000000000001100111000111;
    rom[8663] = 25'b0000000000001100111010011;
    rom[8664] = 25'b0000000000001100111011111;
    rom[8665] = 25'b0000000000001100111101011;
    rom[8666] = 25'b0000000000001100111111000;
    rom[8667] = 25'b0000000000001101000000100;
    rom[8668] = 25'b0000000000001101000010001;
    rom[8669] = 25'b0000000000001101000011101;
    rom[8670] = 25'b0000000000001101000101001;
    rom[8671] = 25'b0000000000001101000110101;
    rom[8672] = 25'b0000000000001101001000010;
    rom[8673] = 25'b0000000000001101001001110;
    rom[8674] = 25'b0000000000001101001011010;
    rom[8675] = 25'b0000000000001101001100110;
    rom[8676] = 25'b0000000000001101001110010;
    rom[8677] = 25'b0000000000001101001111111;
    rom[8678] = 25'b0000000000001101010001011;
    rom[8679] = 25'b0000000000001101010011000;
    rom[8680] = 25'b0000000000001101010100100;
    rom[8681] = 25'b0000000000001101010110000;
    rom[8682] = 25'b0000000000001101010111100;
    rom[8683] = 25'b0000000000001101011001000;
    rom[8684] = 25'b0000000000001101011010101;
    rom[8685] = 25'b0000000000001101011100001;
    rom[8686] = 25'b0000000000001101011101110;
    rom[8687] = 25'b0000000000001101011111010;
    rom[8688] = 25'b0000000000001101100000110;
    rom[8689] = 25'b0000000000001101100010010;
    rom[8690] = 25'b0000000000001101100011110;
    rom[8691] = 25'b0000000000001101100101011;
    rom[8692] = 25'b0000000000001101100110111;
    rom[8693] = 25'b0000000000001101101000100;
    rom[8694] = 25'b0000000000001101101010000;
    rom[8695] = 25'b0000000000001101101011100;
    rom[8696] = 25'b0000000000001101101101000;
    rom[8697] = 25'b0000000000001101101110100;
    rom[8698] = 25'b0000000000001101110000001;
    rom[8699] = 25'b0000000000001101110001101;
    rom[8700] = 25'b0000000000001101110011010;
    rom[8701] = 25'b0000000000001101110100101;
    rom[8702] = 25'b0000000000001101110110001;
    rom[8703] = 25'b0000000000001101110111110;
    rom[8704] = 25'b0000000000001101111001010;
    rom[8705] = 25'b0000000000001101111010110;
    rom[8706] = 25'b0000000000001101111100011;
    rom[8707] = 25'b0000000000001101111101111;
    rom[8708] = 25'b0000000000001101111111011;
    rom[8709] = 25'b0000000000001110000000111;
    rom[8710] = 25'b0000000000001110000010011;
    rom[8711] = 25'b0000000000001110000100000;
    rom[8712] = 25'b0000000000001110000101100;
    rom[8713] = 25'b0000000000001110000111001;
    rom[8714] = 25'b0000000000001110001000101;
    rom[8715] = 25'b0000000000001110001010001;
    rom[8716] = 25'b0000000000001110001011101;
    rom[8717] = 25'b0000000000001110001101001;
    rom[8718] = 25'b0000000000001110001110101;
    rom[8719] = 25'b0000000000001110010000010;
    rom[8720] = 25'b0000000000001110010001110;
    rom[8721] = 25'b0000000000001110010011010;
    rom[8722] = 25'b0000000000001110010100110;
    rom[8723] = 25'b0000000000001110010110010;
    rom[8724] = 25'b0000000000001110010111110;
    rom[8725] = 25'b0000000000001110011001011;
    rom[8726] = 25'b0000000000001110011010111;
    rom[8727] = 25'b0000000000001110011100011;
    rom[8728] = 25'b0000000000001110011110000;
    rom[8729] = 25'b0000000000001110011111100;
    rom[8730] = 25'b0000000000001110100001000;
    rom[8731] = 25'b0000000000001110100010100;
    rom[8732] = 25'b0000000000001110100100000;
    rom[8733] = 25'b0000000000001110100101100;
    rom[8734] = 25'b0000000000001110100111001;
    rom[8735] = 25'b0000000000001110101000101;
    rom[8736] = 25'b0000000000001110101010001;
    rom[8737] = 25'b0000000000001110101011110;
    rom[8738] = 25'b0000000000001110101101001;
    rom[8739] = 25'b0000000000001110101110101;
    rom[8740] = 25'b0000000000001110110000001;
    rom[8741] = 25'b0000000000001110110001110;
    rom[8742] = 25'b0000000000001110110011010;
    rom[8743] = 25'b0000000000001110110100110;
    rom[8744] = 25'b0000000000001110110110011;
    rom[8745] = 25'b0000000000001110110111111;
    rom[8746] = 25'b0000000000001110111001011;
    rom[8747] = 25'b0000000000001110111010111;
    rom[8748] = 25'b0000000000001110111100011;
    rom[8749] = 25'b0000000000001110111101111;
    rom[8750] = 25'b0000000000001110111111011;
    rom[8751] = 25'b0000000000001111000000111;
    rom[8752] = 25'b0000000000001111000010100;
    rom[8753] = 25'b0000000000001111000100000;
    rom[8754] = 25'b0000000000001111000101100;
    rom[8755] = 25'b0000000000001111000111000;
    rom[8756] = 25'b0000000000001111001000100;
    rom[8757] = 25'b0000000000001111001010000;
    rom[8758] = 25'b0000000000001111001011100;
    rom[8759] = 25'b0000000000001111001101000;
    rom[8760] = 25'b0000000000001111001110101;
    rom[8761] = 25'b0000000000001111010000001;
    rom[8762] = 25'b0000000000001111010001101;
    rom[8763] = 25'b0000000000001111010011001;
    rom[8764] = 25'b0000000000001111010100101;
    rom[8765] = 25'b0000000000001111010110001;
    rom[8766] = 25'b0000000000001111010111101;
    rom[8767] = 25'b0000000000001111011001001;
    rom[8768] = 25'b0000000000001111011010101;
    rom[8769] = 25'b0000000000001111011100001;
    rom[8770] = 25'b0000000000001111011101110;
    rom[8771] = 25'b0000000000001111011111010;
    rom[8772] = 25'b0000000000001111100000110;
    rom[8773] = 25'b0000000000001111100010010;
    rom[8774] = 25'b0000000000001111100011110;
    rom[8775] = 25'b0000000000001111100101010;
    rom[8776] = 25'b0000000000001111100110110;
    rom[8777] = 25'b0000000000001111101000010;
    rom[8778] = 25'b0000000000001111101001110;
    rom[8779] = 25'b0000000000001111101011010;
    rom[8780] = 25'b0000000000001111101100110;
    rom[8781] = 25'b0000000000001111101110010;
    rom[8782] = 25'b0000000000001111101111111;
    rom[8783] = 25'b0000000000001111110001011;
    rom[8784] = 25'b0000000000001111110010111;
    rom[8785] = 25'b0000000000001111110100011;
    rom[8786] = 25'b0000000000001111110101111;
    rom[8787] = 25'b0000000000001111110111011;
    rom[8788] = 25'b0000000000001111111000111;
    rom[8789] = 25'b0000000000001111111010011;
    rom[8790] = 25'b0000000000001111111011111;
    rom[8791] = 25'b0000000000001111111101011;
    rom[8792] = 25'b0000000000001111111110111;
    rom[8793] = 25'b0000000000010000000000011;
    rom[8794] = 25'b0000000000010000000001111;
    rom[8795] = 25'b0000000000010000000011011;
    rom[8796] = 25'b0000000000010000000100111;
    rom[8797] = 25'b0000000000010000000110011;
    rom[8798] = 25'b0000000000010000000111111;
    rom[8799] = 25'b0000000000010000001001011;
    rom[8800] = 25'b0000000000010000001010111;
    rom[8801] = 25'b0000000000010000001100011;
    rom[8802] = 25'b0000000000010000001101111;
    rom[8803] = 25'b0000000000010000001111011;
    rom[8804] = 25'b0000000000010000010000111;
    rom[8805] = 25'b0000000000010000010010011;
    rom[8806] = 25'b0000000000010000010011111;
    rom[8807] = 25'b0000000000010000010101010;
    rom[8808] = 25'b0000000000010000010110110;
    rom[8809] = 25'b0000000000010000011000010;
    rom[8810] = 25'b0000000000010000011001110;
    rom[8811] = 25'b0000000000010000011011010;
    rom[8812] = 25'b0000000000010000011100110;
    rom[8813] = 25'b0000000000010000011110010;
    rom[8814] = 25'b0000000000010000011111110;
    rom[8815] = 25'b0000000000010000100001010;
    rom[8816] = 25'b0000000000010000100010110;
    rom[8817] = 25'b0000000000010000100100010;
    rom[8818] = 25'b0000000000010000100101110;
    rom[8819] = 25'b0000000000010000100111010;
    rom[8820] = 25'b0000000000010000101000110;
    rom[8821] = 25'b0000000000010000101010010;
    rom[8822] = 25'b0000000000010000101011110;
    rom[8823] = 25'b0000000000010000101101010;
    rom[8824] = 25'b0000000000010000101110110;
    rom[8825] = 25'b0000000000010000110000010;
    rom[8826] = 25'b0000000000010000110001110;
    rom[8827] = 25'b0000000000010000110011010;
    rom[8828] = 25'b0000000000010000110100110;
    rom[8829] = 25'b0000000000010000110110001;
    rom[8830] = 25'b0000000000010000110111101;
    rom[8831] = 25'b0000000000010000111001001;
    rom[8832] = 25'b0000000000010000111010101;
    rom[8833] = 25'b0000000000010000111100001;
    rom[8834] = 25'b0000000000010000111101100;
    rom[8835] = 25'b0000000000010000111111000;
    rom[8836] = 25'b0000000000010001000000100;
    rom[8837] = 25'b0000000000010001000010000;
    rom[8838] = 25'b0000000000010001000011100;
    rom[8839] = 25'b0000000000010001000101000;
    rom[8840] = 25'b0000000000010001000110011;
    rom[8841] = 25'b0000000000010001000111111;
    rom[8842] = 25'b0000000000010001001001011;
    rom[8843] = 25'b0000000000010001001010111;
    rom[8844] = 25'b0000000000010001001100011;
    rom[8845] = 25'b0000000000010001001101110;
    rom[8846] = 25'b0000000000010001001111010;
    rom[8847] = 25'b0000000000010001010000110;
    rom[8848] = 25'b0000000000010001010010010;
    rom[8849] = 25'b0000000000010001010011110;
    rom[8850] = 25'b0000000000010001010101010;
    rom[8851] = 25'b0000000000010001010110101;
    rom[8852] = 25'b0000000000010001011000001;
    rom[8853] = 25'b0000000000010001011001101;
    rom[8854] = 25'b0000000000010001011011001;
    rom[8855] = 25'b0000000000010001011100101;
    rom[8856] = 25'b0000000000010001011110000;
    rom[8857] = 25'b0000000000010001011111100;
    rom[8858] = 25'b0000000000010001100001000;
    rom[8859] = 25'b0000000000010001100010100;
    rom[8860] = 25'b0000000000010001100100000;
    rom[8861] = 25'b0000000000010001100101011;
    rom[8862] = 25'b0000000000010001100110111;
    rom[8863] = 25'b0000000000010001101000011;
    rom[8864] = 25'b0000000000010001101001110;
    rom[8865] = 25'b0000000000010001101011010;
    rom[8866] = 25'b0000000000010001101100110;
    rom[8867] = 25'b0000000000010001101110001;
    rom[8868] = 25'b0000000000010001101111101;
    rom[8869] = 25'b0000000000010001110001001;
    rom[8870] = 25'b0000000000010001110010100;
    rom[8871] = 25'b0000000000010001110100000;
    rom[8872] = 25'b0000000000010001110101100;
    rom[8873] = 25'b0000000000010001110110111;
    rom[8874] = 25'b0000000000010001111000011;
    rom[8875] = 25'b0000000000010001111001110;
    rom[8876] = 25'b0000000000010001111011010;
    rom[8877] = 25'b0000000000010001111100110;
    rom[8878] = 25'b0000000000010001111110001;
    rom[8879] = 25'b0000000000010001111111101;
    rom[8880] = 25'b0000000000010010000001001;
    rom[8881] = 25'b0000000000010010000010101;
    rom[8882] = 25'b0000000000010010000100001;
    rom[8883] = 25'b0000000000010010000101100;
    rom[8884] = 25'b0000000000010010000111000;
    rom[8885] = 25'b0000000000010010001000011;
    rom[8886] = 25'b0000000000010010001001111;
    rom[8887] = 25'b0000000000010010001011010;
    rom[8888] = 25'b0000000000010010001100110;
    rom[8889] = 25'b0000000000010010001110001;
    rom[8890] = 25'b0000000000010010001111101;
    rom[8891] = 25'b0000000000010010010001000;
    rom[8892] = 25'b0000000000010010010010100;
    rom[8893] = 25'b0000000000010010010100000;
    rom[8894] = 25'b0000000000010010010101100;
    rom[8895] = 25'b0000000000010010010110111;
    rom[8896] = 25'b0000000000010010011000011;
    rom[8897] = 25'b0000000000010010011001110;
    rom[8898] = 25'b0000000000010010011011010;
    rom[8899] = 25'b0000000000010010011100101;
    rom[8900] = 25'b0000000000010010011110001;
    rom[8901] = 25'b0000000000010010011111100;
    rom[8902] = 25'b0000000000010010100000111;
    rom[8903] = 25'b0000000000010010100010011;
    rom[8904] = 25'b0000000000010010100011111;
    rom[8905] = 25'b0000000000010010100101011;
    rom[8906] = 25'b0000000000010010100110110;
    rom[8907] = 25'b0000000000010010101000001;
    rom[8908] = 25'b0000000000010010101001101;
    rom[8909] = 25'b0000000000010010101011000;
    rom[8910] = 25'b0000000000010010101100100;
    rom[8911] = 25'b0000000000010010101101111;
    rom[8912] = 25'b0000000000010010101111010;
    rom[8913] = 25'b0000000000010010110000110;
    rom[8914] = 25'b0000000000010010110010010;
    rom[8915] = 25'b0000000000010010110011101;
    rom[8916] = 25'b0000000000010010110101001;
    rom[8917] = 25'b0000000000010010110110100;
    rom[8918] = 25'b0000000000010010110111111;
    rom[8919] = 25'b0000000000010010111001010;
    rom[8920] = 25'b0000000000010010111010110;
    rom[8921] = 25'b0000000000010010111100010;
    rom[8922] = 25'b0000000000010010111101101;
    rom[8923] = 25'b0000000000010010111111000;
    rom[8924] = 25'b0000000000010011000000100;
    rom[8925] = 25'b0000000000010011000001111;
    rom[8926] = 25'b0000000000010011000011010;
    rom[8927] = 25'b0000000000010011000100110;
    rom[8928] = 25'b0000000000010011000110001;
    rom[8929] = 25'b0000000000010011000111101;
    rom[8930] = 25'b0000000000010011001001000;
    rom[8931] = 25'b0000000000010011001010011;
    rom[8932] = 25'b0000000000010011001011110;
    rom[8933] = 25'b0000000000010011001101010;
    rom[8934] = 25'b0000000000010011001110101;
    rom[8935] = 25'b0000000000010011010000001;
    rom[8936] = 25'b0000000000010011010001100;
    rom[8937] = 25'b0000000000010011010010111;
    rom[8938] = 25'b0000000000010011010100010;
    rom[8939] = 25'b0000000000010011010101110;
    rom[8940] = 25'b0000000000010011010111001;
    rom[8941] = 25'b0000000000010011011000101;
    rom[8942] = 25'b0000000000010011011010000;
    rom[8943] = 25'b0000000000010011011011011;
    rom[8944] = 25'b0000000000010011011100110;
    rom[8945] = 25'b0000000000010011011110001;
    rom[8946] = 25'b0000000000010011011111101;
    rom[8947] = 25'b0000000000010011100001000;
    rom[8948] = 25'b0000000000010011100010011;
    rom[8949] = 25'b0000000000010011100011110;
    rom[8950] = 25'b0000000000010011100101010;
    rom[8951] = 25'b0000000000010011100110101;
    rom[8952] = 25'b0000000000010011101000000;
    rom[8953] = 25'b0000000000010011101001011;
    rom[8954] = 25'b0000000000010011101010110;
    rom[8955] = 25'b0000000000010011101100010;
    rom[8956] = 25'b0000000000010011101101101;
    rom[8957] = 25'b0000000000010011101111000;
    rom[8958] = 25'b0000000000010011110000011;
    rom[8959] = 25'b0000000000010011110001110;
    rom[8960] = 25'b0000000000010011110011010;
    rom[8961] = 25'b0000000000010011110100101;
    rom[8962] = 25'b0000000000010011110110000;
    rom[8963] = 25'b0000000000010011110111011;
    rom[8964] = 25'b0000000000010011111000110;
    rom[8965] = 25'b0000000000010011111010001;
    rom[8966] = 25'b0000000000010011111011100;
    rom[8967] = 25'b0000000000010011111100111;
    rom[8968] = 25'b0000000000010011111110010;
    rom[8969] = 25'b0000000000010011111111110;
    rom[8970] = 25'b0000000000010100000001001;
    rom[8971] = 25'b0000000000010100000010100;
    rom[8972] = 25'b0000000000010100000011111;
    rom[8973] = 25'b0000000000010100000101010;
    rom[8974] = 25'b0000000000010100000110101;
    rom[8975] = 25'b0000000000010100001000000;
    rom[8976] = 25'b0000000000010100001001011;
    rom[8977] = 25'b0000000000010100001010110;
    rom[8978] = 25'b0000000000010100001100001;
    rom[8979] = 25'b0000000000010100001101100;
    rom[8980] = 25'b0000000000010100001110111;
    rom[8981] = 25'b0000000000010100010000010;
    rom[8982] = 25'b0000000000010100010001101;
    rom[8983] = 25'b0000000000010100010011000;
    rom[8984] = 25'b0000000000010100010100100;
    rom[8985] = 25'b0000000000010100010101110;
    rom[8986] = 25'b0000000000010100010111001;
    rom[8987] = 25'b0000000000010100011000100;
    rom[8988] = 25'b0000000000010100011001111;
    rom[8989] = 25'b0000000000010100011011010;
    rom[8990] = 25'b0000000000010100011100101;
    rom[8991] = 25'b0000000000010100011110000;
    rom[8992] = 25'b0000000000010100011111011;
    rom[8993] = 25'b0000000000010100100000101;
    rom[8994] = 25'b0000000000010100100010001;
    rom[8995] = 25'b0000000000010100100011100;
    rom[8996] = 25'b0000000000010100100100110;
    rom[8997] = 25'b0000000000010100100110010;
    rom[8998] = 25'b0000000000010100100111100;
    rom[8999] = 25'b0000000000010100101000111;
    rom[9000] = 25'b0000000000010100101010010;
    rom[9001] = 25'b0000000000010100101011101;
    rom[9002] = 25'b0000000000010100101100111;
    rom[9003] = 25'b0000000000010100101110011;
    rom[9004] = 25'b0000000000010100101111101;
    rom[9005] = 25'b0000000000010100110001000;
    rom[9006] = 25'b0000000000010100110010011;
    rom[9007] = 25'b0000000000010100110011110;
    rom[9008] = 25'b0000000000010100110101000;
    rom[9009] = 25'b0000000000010100110110100;
    rom[9010] = 25'b0000000000010100110111110;
    rom[9011] = 25'b0000000000010100111001001;
    rom[9012] = 25'b0000000000010100111010100;
    rom[9013] = 25'b0000000000010100111011111;
    rom[9014] = 25'b0000000000010100111101001;
    rom[9015] = 25'b0000000000010100111110100;
    rom[9016] = 25'b0000000000010100111111111;
    rom[9017] = 25'b0000000000010101000001001;
    rom[9018] = 25'b0000000000010101000010100;
    rom[9019] = 25'b0000000000010101000011111;
    rom[9020] = 25'b0000000000010101000101010;
    rom[9021] = 25'b0000000000010101000110100;
    rom[9022] = 25'b0000000000010101000111111;
    rom[9023] = 25'b0000000000010101001001010;
    rom[9024] = 25'b0000000000010101001010100;
    rom[9025] = 25'b0000000000010101001011111;
    rom[9026] = 25'b0000000000010101001101010;
    rom[9027] = 25'b0000000000010101001110100;
    rom[9028] = 25'b0000000000010101001111111;
    rom[9029] = 25'b0000000000010101010001010;
    rom[9030] = 25'b0000000000010101010010100;
    rom[9031] = 25'b0000000000010101010011111;
    rom[9032] = 25'b0000000000010101010101001;
    rom[9033] = 25'b0000000000010101010110100;
    rom[9034] = 25'b0000000000010101010111110;
    rom[9035] = 25'b0000000000010101011001001;
    rom[9036] = 25'b0000000000010101011010100;
    rom[9037] = 25'b0000000000010101011011110;
    rom[9038] = 25'b0000000000010101011101001;
    rom[9039] = 25'b0000000000010101011110011;
    rom[9040] = 25'b0000000000010101011111110;
    rom[9041] = 25'b0000000000010101100001000;
    rom[9042] = 25'b0000000000010101100010011;
    rom[9043] = 25'b0000000000010101100011110;
    rom[9044] = 25'b0000000000010101100101000;
    rom[9045] = 25'b0000000000010101100110011;
    rom[9046] = 25'b0000000000010101100111101;
    rom[9047] = 25'b0000000000010101101001000;
    rom[9048] = 25'b0000000000010101101010010;
    rom[9049] = 25'b0000000000010101101011101;
    rom[9050] = 25'b0000000000010101101100111;
    rom[9051] = 25'b0000000000010101101110010;
    rom[9052] = 25'b0000000000010101101111100;
    rom[9053] = 25'b0000000000010101110000110;
    rom[9054] = 25'b0000000000010101110010001;
    rom[9055] = 25'b0000000000010101110011011;
    rom[9056] = 25'b0000000000010101110100101;
    rom[9057] = 25'b0000000000010101110110000;
    rom[9058] = 25'b0000000000010101110111010;
    rom[9059] = 25'b0000000000010101111000100;
    rom[9060] = 25'b0000000000010101111001111;
    rom[9061] = 25'b0000000000010101111011001;
    rom[9062] = 25'b0000000000010101111100100;
    rom[9063] = 25'b0000000000010101111101110;
    rom[9064] = 25'b0000000000010101111111000;
    rom[9065] = 25'b0000000000010110000000010;
    rom[9066] = 25'b0000000000010110000001101;
    rom[9067] = 25'b0000000000010110000010111;
    rom[9068] = 25'b0000000000010110000100001;
    rom[9069] = 25'b0000000000010110000101100;
    rom[9070] = 25'b0000000000010110000110110;
    rom[9071] = 25'b0000000000010110001000000;
    rom[9072] = 25'b0000000000010110001001010;
    rom[9073] = 25'b0000000000010110001010101;
    rom[9074] = 25'b0000000000010110001011111;
    rom[9075] = 25'b0000000000010110001101010;
    rom[9076] = 25'b0000000000010110001110011;
    rom[9077] = 25'b0000000000010110001111110;
    rom[9078] = 25'b0000000000010110010000111;
    rom[9079] = 25'b0000000000010110010010010;
    rom[9080] = 25'b0000000000010110010011100;
    rom[9081] = 25'b0000000000010110010100110;
    rom[9082] = 25'b0000000000010110010110001;
    rom[9083] = 25'b0000000000010110010111011;
    rom[9084] = 25'b0000000000010110011000101;
    rom[9085] = 25'b0000000000010110011001111;
    rom[9086] = 25'b0000000000010110011011001;
    rom[9087] = 25'b0000000000010110011100011;
    rom[9088] = 25'b0000000000010110011101101;
    rom[9089] = 25'b0000000000010110011111000;
    rom[9090] = 25'b0000000000010110100000001;
    rom[9091] = 25'b0000000000010110100001100;
    rom[9092] = 25'b0000000000010110100010101;
    rom[9093] = 25'b0000000000010110100100000;
    rom[9094] = 25'b0000000000010110100101010;
    rom[9095] = 25'b0000000000010110100110100;
    rom[9096] = 25'b0000000000010110100111110;
    rom[9097] = 25'b0000000000010110101000111;
    rom[9098] = 25'b0000000000010110101010010;
    rom[9099] = 25'b0000000000010110101011100;
    rom[9100] = 25'b0000000000010110101100110;
    rom[9101] = 25'b0000000000010110101110000;
    rom[9102] = 25'b0000000000010110101111001;
    rom[9103] = 25'b0000000000010110110000100;
    rom[9104] = 25'b0000000000010110110001110;
    rom[9105] = 25'b0000000000010110110010111;
    rom[9106] = 25'b0000000000010110110100001;
    rom[9107] = 25'b0000000000010110110101100;
    rom[9108] = 25'b0000000000010110110110101;
    rom[9109] = 25'b0000000000010110110111111;
    rom[9110] = 25'b0000000000010110111001001;
    rom[9111] = 25'b0000000000010110111010011;
    rom[9112] = 25'b0000000000010110111011101;
    rom[9113] = 25'b0000000000010110111100111;
    rom[9114] = 25'b0000000000010110111110000;
    rom[9115] = 25'b0000000000010110111111010;
    rom[9116] = 25'b0000000000010111000000100;
    rom[9117] = 25'b0000000000010111000001110;
    rom[9118] = 25'b0000000000010111000011000;
    rom[9119] = 25'b0000000000010111000100010;
    rom[9120] = 25'b0000000000010111000101011;
    rom[9121] = 25'b0000000000010111000110101;
    rom[9122] = 25'b0000000000010111000111111;
    rom[9123] = 25'b0000000000010111001001000;
    rom[9124] = 25'b0000000000010111001010010;
    rom[9125] = 25'b0000000000010111001011100;
    rom[9126] = 25'b0000000000010111001100110;
    rom[9127] = 25'b0000000000010111001101111;
    rom[9128] = 25'b0000000000010111001111001;
    rom[9129] = 25'b0000000000010111010000011;
    rom[9130] = 25'b0000000000010111010001100;
    rom[9131] = 25'b0000000000010111010010110;
    rom[9132] = 25'b0000000000010111010100000;
    rom[9133] = 25'b0000000000010111010101010;
    rom[9134] = 25'b0000000000010111010110011;
    rom[9135] = 25'b0000000000010111010111101;
    rom[9136] = 25'b0000000000010111011000111;
    rom[9137] = 25'b0000000000010111011010000;
    rom[9138] = 25'b0000000000010111011011001;
    rom[9139] = 25'b0000000000010111011100011;
    rom[9140] = 25'b0000000000010111011101101;
    rom[9141] = 25'b0000000000010111011110111;
    rom[9142] = 25'b0000000000010111100000000;
    rom[9143] = 25'b0000000000010111100001001;
    rom[9144] = 25'b0000000000010111100010011;
    rom[9145] = 25'b0000000000010111100011101;
    rom[9146] = 25'b0000000000010111100100110;
    rom[9147] = 25'b0000000000010111100101111;
    rom[9148] = 25'b0000000000010111100111001;
    rom[9149] = 25'b0000000000010111101000011;
    rom[9150] = 25'b0000000000010111101001100;
    rom[9151] = 25'b0000000000010111101010101;
    rom[9152] = 25'b0000000000010111101011111;
    rom[9153] = 25'b0000000000010111101101000;
    rom[9154] = 25'b0000000000010111101110010;
    rom[9155] = 25'b0000000000010111101111011;
    rom[9156] = 25'b0000000000010111110000100;
    rom[9157] = 25'b0000000000010111110001110;
    rom[9158] = 25'b0000000000010111110010111;
    rom[9159] = 25'b0000000000010111110100001;
    rom[9160] = 25'b0000000000010111110101010;
    rom[9161] = 25'b0000000000010111110110100;
    rom[9162] = 25'b0000000000010111110111100;
    rom[9163] = 25'b0000000000010111111000110;
    rom[9164] = 25'b0000000000010111111001111;
    rom[9165] = 25'b0000000000010111111011000;
    rom[9166] = 25'b0000000000010111111100010;
    rom[9167] = 25'b0000000000010111111101011;
    rom[9168] = 25'b0000000000010111111110101;
    rom[9169] = 25'b0000000000010111111111101;
    rom[9170] = 25'b0000000000011000000000110;
    rom[9171] = 25'b0000000000011000000010000;
    rom[9172] = 25'b0000000000011000000011001;
    rom[9173] = 25'b0000000000011000000100011;
    rom[9174] = 25'b0000000000011000000101100;
    rom[9175] = 25'b0000000000011000000110101;
    rom[9176] = 25'b0000000000011000000111110;
    rom[9177] = 25'b0000000000011000001000111;
    rom[9178] = 25'b0000000000011000001010000;
    rom[9179] = 25'b0000000000011000001011001;
    rom[9180] = 25'b0000000000011000001100010;
    rom[9181] = 25'b0000000000011000001101100;
    rom[9182] = 25'b0000000000011000001110101;
    rom[9183] = 25'b0000000000011000001111110;
    rom[9184] = 25'b0000000000011000010000111;
    rom[9185] = 25'b0000000000011000010010000;
    rom[9186] = 25'b0000000000011000010011001;
    rom[9187] = 25'b0000000000011000010100010;
    rom[9188] = 25'b0000000000011000010101100;
    rom[9189] = 25'b0000000000011000010110101;
    rom[9190] = 25'b0000000000011000010111101;
    rom[9191] = 25'b0000000000011000011000110;
    rom[9192] = 25'b0000000000011000011001111;
    rom[9193] = 25'b0000000000011000011011000;
    rom[9194] = 25'b0000000000011000011100001;
    rom[9195] = 25'b0000000000011000011101010;
    rom[9196] = 25'b0000000000011000011110011;
    rom[9197] = 25'b0000000000011000011111100;
    rom[9198] = 25'b0000000000011000100000101;
    rom[9199] = 25'b0000000000011000100001101;
    rom[9200] = 25'b0000000000011000100010110;
    rom[9201] = 25'b0000000000011000100011111;
    rom[9202] = 25'b0000000000011000100101000;
    rom[9203] = 25'b0000000000011000100110001;
    rom[9204] = 25'b0000000000011000100111010;
    rom[9205] = 25'b0000000000011000101000011;
    rom[9206] = 25'b0000000000011000101001011;
    rom[9207] = 25'b0000000000011000101010100;
    rom[9208] = 25'b0000000000011000101011101;
    rom[9209] = 25'b0000000000011000101100110;
    rom[9210] = 25'b0000000000011000101101111;
    rom[9211] = 25'b0000000000011000101111000;
    rom[9212] = 25'b0000000000011000110000000;
    rom[9213] = 25'b0000000000011000110001001;
    rom[9214] = 25'b0000000000011000110010010;
    rom[9215] = 25'b0000000000011000110011011;
    rom[9216] = 25'b0000000000011000110100100;
    rom[9217] = 25'b0000000000011000110101100;
    rom[9218] = 25'b0000000000011000110110101;
    rom[9219] = 25'b0000000000011000110111101;
    rom[9220] = 25'b0000000000011000111000110;
    rom[9221] = 25'b0000000000011000111001111;
    rom[9222] = 25'b0000000000011000111010111;
    rom[9223] = 25'b0000000000011000111100000;
    rom[9224] = 25'b0000000000011000111101000;
    rom[9225] = 25'b0000000000011000111110001;
    rom[9226] = 25'b0000000000011000111111010;
    rom[9227] = 25'b0000000000011001000000010;
    rom[9228] = 25'b0000000000011001000001011;
    rom[9229] = 25'b0000000000011001000010011;
    rom[9230] = 25'b0000000000011001000011100;
    rom[9231] = 25'b0000000000011001000100100;
    rom[9232] = 25'b0000000000011001000101101;
    rom[9233] = 25'b0000000000011001000110101;
    rom[9234] = 25'b0000000000011001000111110;
    rom[9235] = 25'b0000000000011001001000110;
    rom[9236] = 25'b0000000000011001001001111;
    rom[9237] = 25'b0000000000011001001010111;
    rom[9238] = 25'b0000000000011001001011111;
    rom[9239] = 25'b0000000000011001001101000;
    rom[9240] = 25'b0000000000011001001110000;
    rom[9241] = 25'b0000000000011001001111001;
    rom[9242] = 25'b0000000000011001010000001;
    rom[9243] = 25'b0000000000011001010001001;
    rom[9244] = 25'b0000000000011001010010010;
    rom[9245] = 25'b0000000000011001010011010;
    rom[9246] = 25'b0000000000011001010100010;
    rom[9247] = 25'b0000000000011001010101011;
    rom[9248] = 25'b0000000000011001010110011;
    rom[9249] = 25'b0000000000011001010111011;
    rom[9250] = 25'b0000000000011001011000011;
    rom[9251] = 25'b0000000000011001011001011;
    rom[9252] = 25'b0000000000011001011010100;
    rom[9253] = 25'b0000000000011001011011100;
    rom[9254] = 25'b0000000000011001011100100;
    rom[9255] = 25'b0000000000011001011101100;
    rom[9256] = 25'b0000000000011001011110101;
    rom[9257] = 25'b0000000000011001011111101;
    rom[9258] = 25'b0000000000011001100000101;
    rom[9259] = 25'b0000000000011001100001101;
    rom[9260] = 25'b0000000000011001100010101;
    rom[9261] = 25'b0000000000011001100011110;
    rom[9262] = 25'b0000000000011001100100110;
    rom[9263] = 25'b0000000000011001100101101;
    rom[9264] = 25'b0000000000011001100110110;
    rom[9265] = 25'b0000000000011001100111110;
    rom[9266] = 25'b0000000000011001101000110;
    rom[9267] = 25'b0000000000011001101001110;
    rom[9268] = 25'b0000000000011001101010110;
    rom[9269] = 25'b0000000000011001101011110;
    rom[9270] = 25'b0000000000011001101100110;
    rom[9271] = 25'b0000000000011001101101110;
    rom[9272] = 25'b0000000000011001101110110;
    rom[9273] = 25'b0000000000011001101111110;
    rom[9274] = 25'b0000000000011001110000101;
    rom[9275] = 25'b0000000000011001110001110;
    rom[9276] = 25'b0000000000011001110010110;
    rom[9277] = 25'b0000000000011001110011101;
    rom[9278] = 25'b0000000000011001110100110;
    rom[9279] = 25'b0000000000011001110101101;
    rom[9280] = 25'b0000000000011001110110101;
    rom[9281] = 25'b0000000000011001110111101;
    rom[9282] = 25'b0000000000011001111000101;
    rom[9283] = 25'b0000000000011001111001100;
    rom[9284] = 25'b0000000000011001111010101;
    rom[9285] = 25'b0000000000011001111011100;
    rom[9286] = 25'b0000000000011001111100100;
    rom[9287] = 25'b0000000000011001111101100;
    rom[9288] = 25'b0000000000011001111110011;
    rom[9289] = 25'b0000000000011001111111100;
    rom[9290] = 25'b0000000000011010000000011;
    rom[9291] = 25'b0000000000011010000001010;
    rom[9292] = 25'b0000000000011010000010011;
    rom[9293] = 25'b0000000000011010000011010;
    rom[9294] = 25'b0000000000011010000100010;
    rom[9295] = 25'b0000000000011010000101010;
    rom[9296] = 25'b0000000000011010000110001;
    rom[9297] = 25'b0000000000011010000111001;
    rom[9298] = 25'b0000000000011010001000000;
    rom[9299] = 25'b0000000000011010001001000;
    rom[9300] = 25'b0000000000011010001001111;
    rom[9301] = 25'b0000000000011010001010111;
    rom[9302] = 25'b0000000000011010001011111;
    rom[9303] = 25'b0000000000011010001100110;
    rom[9304] = 25'b0000000000011010001101110;
    rom[9305] = 25'b0000000000011010001110101;
    rom[9306] = 25'b0000000000011010001111101;
    rom[9307] = 25'b0000000000011010010000100;
    rom[9308] = 25'b0000000000011010010001100;
    rom[9309] = 25'b0000000000011010010010011;
    rom[9310] = 25'b0000000000011010010011011;
    rom[9311] = 25'b0000000000011010010100010;
    rom[9312] = 25'b0000000000011010010101010;
    rom[9313] = 25'b0000000000011010010110001;
    rom[9314] = 25'b0000000000011010010111001;
    rom[9315] = 25'b0000000000011010010111111;
    rom[9316] = 25'b0000000000011010011000111;
    rom[9317] = 25'b0000000000011010011001110;
    rom[9318] = 25'b0000000000011010011010110;
    rom[9319] = 25'b0000000000011010011011101;
    rom[9320] = 25'b0000000000011010011100101;
    rom[9321] = 25'b0000000000011010011101011;
    rom[9322] = 25'b0000000000011010011110011;
    rom[9323] = 25'b0000000000011010011111010;
    rom[9324] = 25'b0000000000011010100000001;
    rom[9325] = 25'b0000000000011010100001000;
    rom[9326] = 25'b0000000000011010100010000;
    rom[9327] = 25'b0000000000011010100010111;
    rom[9328] = 25'b0000000000011010100011110;
    rom[9329] = 25'b0000000000011010100100110;
    rom[9330] = 25'b0000000000011010100101100;
    rom[9331] = 25'b0000000000011010100110100;
    rom[9332] = 25'b0000000000011010100111011;
    rom[9333] = 25'b0000000000011010101000010;
    rom[9334] = 25'b0000000000011010101001001;
    rom[9335] = 25'b0000000000011010101010000;
    rom[9336] = 25'b0000000000011010101010111;
    rom[9337] = 25'b0000000000011010101011110;
    rom[9338] = 25'b0000000000011010101100101;
    rom[9339] = 25'b0000000000011010101101100;
    rom[9340] = 25'b0000000000011010101110011;
    rom[9341] = 25'b0000000000011010101111010;
    rom[9342] = 25'b0000000000011010110000010;
    rom[9343] = 25'b0000000000011010110001000;
    rom[9344] = 25'b0000000000011010110001111;
    rom[9345] = 25'b0000000000011010110010110;
    rom[9346] = 25'b0000000000011010110011101;
    rom[9347] = 25'b0000000000011010110100100;
    rom[9348] = 25'b0000000000011010110101011;
    rom[9349] = 25'b0000000000011010110110001;
    rom[9350] = 25'b0000000000011010110111000;
    rom[9351] = 25'b0000000000011010111000000;
    rom[9352] = 25'b0000000000011010111000110;
    rom[9353] = 25'b0000000000011010111001101;
    rom[9354] = 25'b0000000000011010111010100;
    rom[9355] = 25'b0000000000011010111011010;
    rom[9356] = 25'b0000000000011010111100001;
    rom[9357] = 25'b0000000000011010111101000;
    rom[9358] = 25'b0000000000011010111101111;
    rom[9359] = 25'b0000000000011010111110101;
    rom[9360] = 25'b0000000000011010111111100;
    rom[9361] = 25'b0000000000011011000000011;
    rom[9362] = 25'b0000000000011011000001001;
    rom[9363] = 25'b0000000000011011000010000;
    rom[9364] = 25'b0000000000011011000010111;
    rom[9365] = 25'b0000000000011011000011110;
    rom[9366] = 25'b0000000000011011000100100;
    rom[9367] = 25'b0000000000011011000101010;
    rom[9368] = 25'b0000000000011011000110001;
    rom[9369] = 25'b0000000000011011000111000;
    rom[9370] = 25'b0000000000011011000111111;
    rom[9371] = 25'b0000000000011011001000101;
    rom[9372] = 25'b0000000000011011001001011;
    rom[9373] = 25'b0000000000011011001010010;
    rom[9374] = 25'b0000000000011011001011001;
    rom[9375] = 25'b0000000000011011001011111;
    rom[9376] = 25'b0000000000011011001100101;
    rom[9377] = 25'b0000000000011011001101011;
    rom[9378] = 25'b0000000000011011001110010;
    rom[9379] = 25'b0000000000011011001111001;
    rom[9380] = 25'b0000000000011011001111111;
    rom[9381] = 25'b0000000000011011010000101;
    rom[9382] = 25'b0000000000011011010001011;
    rom[9383] = 25'b0000000000011011010010010;
    rom[9384] = 25'b0000000000011011010011000;
    rom[9385] = 25'b0000000000011011010011111;
    rom[9386] = 25'b0000000000011011010100101;
    rom[9387] = 25'b0000000000011011010101011;
    rom[9388] = 25'b0000000000011011010110010;
    rom[9389] = 25'b0000000000011011010111000;
    rom[9390] = 25'b0000000000011011010111110;
    rom[9391] = 25'b0000000000011011011000100;
    rom[9392] = 25'b0000000000011011011001010;
    rom[9393] = 25'b0000000000011011011010000;
    rom[9394] = 25'b0000000000011011011010111;
    rom[9395] = 25'b0000000000011011011011101;
    rom[9396] = 25'b0000000000011011011100011;
    rom[9397] = 25'b0000000000011011011101001;
    rom[9398] = 25'b0000000000011011011110000;
    rom[9399] = 25'b0000000000011011011110110;
    rom[9400] = 25'b0000000000011011011111100;
    rom[9401] = 25'b0000000000011011100000010;
    rom[9402] = 25'b0000000000011011100000111;
    rom[9403] = 25'b0000000000011011100001101;
    rom[9404] = 25'b0000000000011011100010011;
    rom[9405] = 25'b0000000000011011100011001;
    rom[9406] = 25'b0000000000011011100011111;
    rom[9407] = 25'b0000000000011011100100101;
    rom[9408] = 25'b0000000000011011100101011;
    rom[9409] = 25'b0000000000011011100110001;
    rom[9410] = 25'b0000000000011011100110111;
    rom[9411] = 25'b0000000000011011100111101;
    rom[9412] = 25'b0000000000011011101000011;
    rom[9413] = 25'b0000000000011011101001001;
    rom[9414] = 25'b0000000000011011101001110;
    rom[9415] = 25'b0000000000011011101010100;
    rom[9416] = 25'b0000000000011011101011010;
    rom[9417] = 25'b0000000000011011101100000;
    rom[9418] = 25'b0000000000011011101100110;
    rom[9419] = 25'b0000000000011011101101100;
    rom[9420] = 25'b0000000000011011101110010;
    rom[9421] = 25'b0000000000011011101110111;
    rom[9422] = 25'b0000000000011011101111101;
    rom[9423] = 25'b0000000000011011110000011;
    rom[9424] = 25'b0000000000011011110001000;
    rom[9425] = 25'b0000000000011011110001110;
    rom[9426] = 25'b0000000000011011110010011;
    rom[9427] = 25'b0000000000011011110011001;
    rom[9428] = 25'b0000000000011011110011111;
    rom[9429] = 25'b0000000000011011110100100;
    rom[9430] = 25'b0000000000011011110101010;
    rom[9431] = 25'b0000000000011011110110000;
    rom[9432] = 25'b0000000000011011110110101;
    rom[9433] = 25'b0000000000011011110111011;
    rom[9434] = 25'b0000000000011011111000000;
    rom[9435] = 25'b0000000000011011111000110;
    rom[9436] = 25'b0000000000011011111001011;
    rom[9437] = 25'b0000000000011011111010000;
    rom[9438] = 25'b0000000000011011111010110;
    rom[9439] = 25'b0000000000011011111011100;
    rom[9440] = 25'b0000000000011011111100001;
    rom[9441] = 25'b0000000000011011111100110;
    rom[9442] = 25'b0000000000011011111101011;
    rom[9443] = 25'b0000000000011011111110001;
    rom[9444] = 25'b0000000000011011111110111;
    rom[9445] = 25'b0000000000011011111111100;
    rom[9446] = 25'b0000000000011100000000001;
    rom[9447] = 25'b0000000000011100000000110;
    rom[9448] = 25'b0000000000011100000001011;
    rom[9449] = 25'b0000000000011100000010001;
    rom[9450] = 25'b0000000000011100000010110;
    rom[9451] = 25'b0000000000011100000011011;
    rom[9452] = 25'b0000000000011100000100000;
    rom[9453] = 25'b0000000000011100000100110;
    rom[9454] = 25'b0000000000011100000101011;
    rom[9455] = 25'b0000000000011100000110000;
    rom[9456] = 25'b0000000000011100000110101;
    rom[9457] = 25'b0000000000011100000111011;
    rom[9458] = 25'b0000000000011100000111111;
    rom[9459] = 25'b0000000000011100001000100;
    rom[9460] = 25'b0000000000011100001001001;
    rom[9461] = 25'b0000000000011100001001111;
    rom[9462] = 25'b0000000000011100001010100;
    rom[9463] = 25'b0000000000011100001011000;
    rom[9464] = 25'b0000000000011100001011110;
    rom[9465] = 25'b0000000000011100001100011;
    rom[9466] = 25'b0000000000011100001100111;
    rom[9467] = 25'b0000000000011100001101101;
    rom[9468] = 25'b0000000000011100001110010;
    rom[9469] = 25'b0000000000011100001110110;
    rom[9470] = 25'b0000000000011100001111100;
    rom[9471] = 25'b0000000000011100010000000;
    rom[9472] = 25'b0000000000011100010000101;
    rom[9473] = 25'b0000000000011100010001010;
    rom[9474] = 25'b0000000000011100010001111;
    rom[9475] = 25'b0000000000011100010010011;
    rom[9476] = 25'b0000000000011100010011000;
    rom[9477] = 25'b0000000000011100010011101;
    rom[9478] = 25'b0000000000011100010100010;
    rom[9479] = 25'b0000000000011100010100111;
    rom[9480] = 25'b0000000000011100010101011;
    rom[9481] = 25'b0000000000011100010110000;
    rom[9482] = 25'b0000000000011100010110100;
    rom[9483] = 25'b0000000000011100010111010;
    rom[9484] = 25'b0000000000011100010111110;
    rom[9485] = 25'b0000000000011100011000011;
    rom[9486] = 25'b0000000000011100011000111;
    rom[9487] = 25'b0000000000011100011001011;
    rom[9488] = 25'b0000000000011100011010001;
    rom[9489] = 25'b0000000000011100011010101;
    rom[9490] = 25'b0000000000011100011011010;
    rom[9491] = 25'b0000000000011100011011110;
    rom[9492] = 25'b0000000000011100011100011;
    rom[9493] = 25'b0000000000011100011100111;
    rom[9494] = 25'b0000000000011100011101100;
    rom[9495] = 25'b0000000000011100011110000;
    rom[9496] = 25'b0000000000011100011110101;
    rom[9497] = 25'b0000000000011100011111001;
    rom[9498] = 25'b0000000000011100011111110;
    rom[9499] = 25'b0000000000011100100000001;
    rom[9500] = 25'b0000000000011100100000110;
    rom[9501] = 25'b0000000000011100100001010;
    rom[9502] = 25'b0000000000011100100001111;
    rom[9503] = 25'b0000000000011100100010011;
    rom[9504] = 25'b0000000000011100100010111;
    rom[9505] = 25'b0000000000011100100011011;
    rom[9506] = 25'b0000000000011100100100000;
    rom[9507] = 25'b0000000000011100100100100;
    rom[9508] = 25'b0000000000011100100101000;
    rom[9509] = 25'b0000000000011100100101101;
    rom[9510] = 25'b0000000000011100100110000;
    rom[9511] = 25'b0000000000011100100110101;
    rom[9512] = 25'b0000000000011100100111001;
    rom[9513] = 25'b0000000000011100100111101;
    rom[9514] = 25'b0000000000011100101000001;
    rom[9515] = 25'b0000000000011100101000101;
    rom[9516] = 25'b0000000000011100101001001;
    rom[9517] = 25'b0000000000011100101001101;
    rom[9518] = 25'b0000000000011100101010001;
    rom[9519] = 25'b0000000000011100101010110;
    rom[9520] = 25'b0000000000011100101011001;
    rom[9521] = 25'b0000000000011100101011101;
    rom[9522] = 25'b0000000000011100101100010;
    rom[9523] = 25'b0000000000011100101100101;
    rom[9524] = 25'b0000000000011100101101001;
    rom[9525] = 25'b0000000000011100101101101;
    rom[9526] = 25'b0000000000011100101110001;
    rom[9527] = 25'b0000000000011100101110101;
    rom[9528] = 25'b0000000000011100101111001;
    rom[9529] = 25'b0000000000011100101111101;
    rom[9530] = 25'b0000000000011100110000000;
    rom[9531] = 25'b0000000000011100110000100;
    rom[9532] = 25'b0000000000011100110001000;
    rom[9533] = 25'b0000000000011100110001011;
    rom[9534] = 25'b0000000000011100110001111;
    rom[9535] = 25'b0000000000011100110010011;
    rom[9536] = 25'b0000000000011100110010111;
    rom[9537] = 25'b0000000000011100110011010;
    rom[9538] = 25'b0000000000011100110011110;
    rom[9539] = 25'b0000000000011100110100010;
    rom[9540] = 25'b0000000000011100110100110;
    rom[9541] = 25'b0000000000011100110101001;
    rom[9542] = 25'b0000000000011100110101100;
    rom[9543] = 25'b0000000000011100110110000;
    rom[9544] = 25'b0000000000011100110110100;
    rom[9545] = 25'b0000000000011100110111000;
    rom[9546] = 25'b0000000000011100110111011;
    rom[9547] = 25'b0000000000011100110111110;
    rom[9548] = 25'b0000000000011100111000010;
    rom[9549] = 25'b0000000000011100111000101;
    rom[9550] = 25'b0000000000011100111001001;
    rom[9551] = 25'b0000000000011100111001100;
    rom[9552] = 25'b0000000000011100111001111;
    rom[9553] = 25'b0000000000011100111010011;
    rom[9554] = 25'b0000000000011100111010110;
    rom[9555] = 25'b0000000000011100111011001;
    rom[9556] = 25'b0000000000011100111011101;
    rom[9557] = 25'b0000000000011100111100000;
    rom[9558] = 25'b0000000000011100111100100;
    rom[9559] = 25'b0000000000011100111100111;
    rom[9560] = 25'b0000000000011100111101010;
    rom[9561] = 25'b0000000000011100111101101;
    rom[9562] = 25'b0000000000011100111110000;
    rom[9563] = 25'b0000000000011100111110011;
    rom[9564] = 25'b0000000000011100111110111;
    rom[9565] = 25'b0000000000011100111111010;
    rom[9566] = 25'b0000000000011100111111101;
    rom[9567] = 25'b0000000000011101000000000;
    rom[9568] = 25'b0000000000011101000000011;
    rom[9569] = 25'b0000000000011101000000110;
    rom[9570] = 25'b0000000000011101000001010;
    rom[9571] = 25'b0000000000011101000001101;
    rom[9572] = 25'b0000000000011101000010000;
    rom[9573] = 25'b0000000000011101000010011;
    rom[9574] = 25'b0000000000011101000010110;
    rom[9575] = 25'b0000000000011101000011001;
    rom[9576] = 25'b0000000000011101000011011;
    rom[9577] = 25'b0000000000011101000011110;
    rom[9578] = 25'b0000000000011101000100001;
    rom[9579] = 25'b0000000000011101000100100;
    rom[9580] = 25'b0000000000011101000100111;
    rom[9581] = 25'b0000000000011101000101010;
    rom[9582] = 25'b0000000000011101000101101;
    rom[9583] = 25'b0000000000011101000101111;
    rom[9584] = 25'b0000000000011101000110010;
    rom[9585] = 25'b0000000000011101000110101;
    rom[9586] = 25'b0000000000011101000110111;
    rom[9587] = 25'b0000000000011101000111010;
    rom[9588] = 25'b0000000000011101000111101;
    rom[9589] = 25'b0000000000011101001000000;
    rom[9590] = 25'b0000000000011101001000011;
    rom[9591] = 25'b0000000000011101001000101;
    rom[9592] = 25'b0000000000011101001001000;
    rom[9593] = 25'b0000000000011101001001010;
    rom[9594] = 25'b0000000000011101001001101;
    rom[9595] = 25'b0000000000011101001001111;
    rom[9596] = 25'b0000000000011101001010010;
    rom[9597] = 25'b0000000000011101001010100;
    rom[9598] = 25'b0000000000011101001010111;
    rom[9599] = 25'b0000000000011101001011010;
    rom[9600] = 25'b0000000000011101001011100;
    rom[9601] = 25'b0000000000011101001011110;
    rom[9602] = 25'b0000000000011101001100001;
    rom[9603] = 25'b0000000000011101001100011;
    rom[9604] = 25'b0000000000011101001100110;
    rom[9605] = 25'b0000000000011101001101000;
    rom[9606] = 25'b0000000000011101001101010;
    rom[9607] = 25'b0000000000011101001101100;
    rom[9608] = 25'b0000000000011101001101111;
    rom[9609] = 25'b0000000000011101001110010;
    rom[9610] = 25'b0000000000011101001110100;
    rom[9611] = 25'b0000000000011101001110110;
    rom[9612] = 25'b0000000000011101001111000;
    rom[9613] = 25'b0000000000011101001111011;
    rom[9614] = 25'b0000000000011101001111100;
    rom[9615] = 25'b0000000000011101001111110;
    rom[9616] = 25'b0000000000011101010000001;
    rom[9617] = 25'b0000000000011101010000011;
    rom[9618] = 25'b0000000000011101010000101;
    rom[9619] = 25'b0000000000011101010000111;
    rom[9620] = 25'b0000000000011101010001001;
    rom[9621] = 25'b0000000000011101010001011;
    rom[9622] = 25'b0000000000011101010001101;
    rom[9623] = 25'b0000000000011101010001111;
    rom[9624] = 25'b0000000000011101010010001;
    rom[9625] = 25'b0000000000011101010010011;
    rom[9626] = 25'b0000000000011101010010101;
    rom[9627] = 25'b0000000000011101010010111;
    rom[9628] = 25'b0000000000011101010011001;
    rom[9629] = 25'b0000000000011101010011011;
    rom[9630] = 25'b0000000000011101010011101;
    rom[9631] = 25'b0000000000011101010011110;
    rom[9632] = 25'b0000000000011101010100001;
    rom[9633] = 25'b0000000000011101010100010;
    rom[9634] = 25'b0000000000011101010100100;
    rom[9635] = 25'b0000000000011101010100110;
    rom[9636] = 25'b0000000000011101010100111;
    rom[9637] = 25'b0000000000011101010101001;
    rom[9638] = 25'b0000000000011101010101011;
    rom[9639] = 25'b0000000000011101010101101;
    rom[9640] = 25'b0000000000011101010101110;
    rom[9641] = 25'b0000000000011101010110000;
    rom[9642] = 25'b0000000000011101010110001;
    rom[9643] = 25'b0000000000011101010110011;
    rom[9644] = 25'b0000000000011101010110101;
    rom[9645] = 25'b0000000000011101010110110;
    rom[9646] = 25'b0000000000011101010111000;
    rom[9647] = 25'b0000000000011101010111001;
    rom[9648] = 25'b0000000000011101010111011;
    rom[9649] = 25'b0000000000011101010111100;
    rom[9650] = 25'b0000000000011101010111110;
    rom[9651] = 25'b0000000000011101010111111;
    rom[9652] = 25'b0000000000011101011000001;
    rom[9653] = 25'b0000000000011101011000010;
    rom[9654] = 25'b0000000000011101011000011;
    rom[9655] = 25'b0000000000011101011000101;
    rom[9656] = 25'b0000000000011101011000110;
    rom[9657] = 25'b0000000000011101011001000;
    rom[9658] = 25'b0000000000011101011001000;
    rom[9659] = 25'b0000000000011101011001010;
    rom[9660] = 25'b0000000000011101011001011;
    rom[9661] = 25'b0000000000011101011001100;
    rom[9662] = 25'b0000000000011101011001101;
    rom[9663] = 25'b0000000000011101011001111;
    rom[9664] = 25'b0000000000011101011010000;
    rom[9665] = 25'b0000000000011101011010001;
    rom[9666] = 25'b0000000000011101011010010;
    rom[9667] = 25'b0000000000011101011010011;
    rom[9668] = 25'b0000000000011101011010100;
    rom[9669] = 25'b0000000000011101011010101;
    rom[9670] = 25'b0000000000011101011010110;
    rom[9671] = 25'b0000000000011101011010111;
    rom[9672] = 25'b0000000000011101011011001;
    rom[9673] = 25'b0000000000011101011011001;
    rom[9674] = 25'b0000000000011101011011010;
    rom[9675] = 25'b0000000000011101011011011;
    rom[9676] = 25'b0000000000011101011011100;
    rom[9677] = 25'b0000000000011101011011101;
    rom[9678] = 25'b0000000000011101011011110;
    rom[9679] = 25'b0000000000011101011011111;
    rom[9680] = 25'b0000000000011101011011111;
    rom[9681] = 25'b0000000000011101011100000;
    rom[9682] = 25'b0000000000011101011100001;
    rom[9683] = 25'b0000000000011101011100010;
    rom[9684] = 25'b0000000000011101011100010;
    rom[9685] = 25'b0000000000011101011100011;
    rom[9686] = 25'b0000000000011101011100100;
    rom[9687] = 25'b0000000000011101011100101;
    rom[9688] = 25'b0000000000011101011100101;
    rom[9689] = 25'b0000000000011101011100110;
    rom[9690] = 25'b0000000000011101011100111;
    rom[9691] = 25'b0000000000011101011101000;
    rom[9692] = 25'b0000000000011101011101000;
    rom[9693] = 25'b0000000000011101011101000;
    rom[9694] = 25'b0000000000011101011101001;
    rom[9695] = 25'b0000000000011101011101001;
    rom[9696] = 25'b0000000000011101011101010;
    rom[9697] = 25'b0000000000011101011101011;
    rom[9698] = 25'b0000000000011101011101011;
    rom[9699] = 25'b0000000000011101011101011;
    rom[9700] = 25'b0000000000011101011101011;
    rom[9701] = 25'b0000000000011101011101100;
    rom[9702] = 25'b0000000000011101011101100;
    rom[9703] = 25'b0000000000011101011101101;
    rom[9704] = 25'b0000000000011101011101101;
    rom[9705] = 25'b0000000000011101011101110;
    rom[9706] = 25'b0000000000011101011101110;
    rom[9707] = 25'b0000000000011101011101110;
    rom[9708] = 25'b0000000000011101011101110;
    rom[9709] = 25'b0000000000011101011101110;
    rom[9710] = 25'b0000000000011101011101110;
    rom[9711] = 25'b0000000000011101011101110;
    rom[9712] = 25'b0000000000011101011101111;
    rom[9713] = 25'b0000000000011101011101111;
    rom[9714] = 25'b0000000000011101011101111;
    rom[9715] = 25'b0000000000011101011101111;
    rom[9716] = 25'b0000000000011101011101111;
    rom[9717] = 25'b0000000000011101011101111;
    rom[9718] = 25'b0000000000011101011101111;
    rom[9719] = 25'b0000000000011101011101111;
    rom[9720] = 25'b0000000000011101011101111;
    rom[9721] = 25'b0000000000011101011101111;
    rom[9722] = 25'b0000000000011101011101111;
    rom[9723] = 25'b0000000000011101011101111;
    rom[9724] = 25'b0000000000011101011101111;
    rom[9725] = 25'b0000000000011101011101110;
    rom[9726] = 25'b0000000000011101011101110;
    rom[9727] = 25'b0000000000011101011101110;
    rom[9728] = 25'b0000000000011101011101110;
    rom[9729] = 25'b0000000000011101011101110;
    rom[9730] = 25'b0000000000011101011101110;
    rom[9731] = 25'b0000000000011101011101110;
    rom[9732] = 25'b0000000000011101011101101;
    rom[9733] = 25'b0000000000011101011101101;
    rom[9734] = 25'b0000000000011101011101100;
    rom[9735] = 25'b0000000000011101011101100;
    rom[9736] = 25'b0000000000011101011101011;
    rom[9737] = 25'b0000000000011101011101011;
    rom[9738] = 25'b0000000000011101011101011;
    rom[9739] = 25'b0000000000011101011101011;
    rom[9740] = 25'b0000000000011101011101010;
    rom[9741] = 25'b0000000000011101011101001;
    rom[9742] = 25'b0000000000011101011101001;
    rom[9743] = 25'b0000000000011101011101000;
    rom[9744] = 25'b0000000000011101011101000;
    rom[9745] = 25'b0000000000011101011101000;
    rom[9746] = 25'b0000000000011101011100111;
    rom[9747] = 25'b0000000000011101011100110;
    rom[9748] = 25'b0000000000011101011100101;
    rom[9749] = 25'b0000000000011101011100101;
    rom[9750] = 25'b0000000000011101011100100;
    rom[9751] = 25'b0000000000011101011100011;
    rom[9752] = 25'b0000000000011101011100010;
    rom[9753] = 25'b0000000000011101011100010;
    rom[9754] = 25'b0000000000011101011100001;
    rom[9755] = 25'b0000000000011101011100000;
    rom[9756] = 25'b0000000000011101011011111;
    rom[9757] = 25'b0000000000011101011011111;
    rom[9758] = 25'b0000000000011101011011110;
    rom[9759] = 25'b0000000000011101011011101;
    rom[9760] = 25'b0000000000011101011011100;
    rom[9761] = 25'b0000000000011101011011011;
    rom[9762] = 25'b0000000000011101011011010;
    rom[9763] = 25'b0000000000011101011011001;
    rom[9764] = 25'b0000000000011101011011000;
    rom[9765] = 25'b0000000000011101011010111;
    rom[9766] = 25'b0000000000011101011010110;
    rom[9767] = 25'b0000000000011101011010101;
    rom[9768] = 25'b0000000000011101011010100;
    rom[9769] = 25'b0000000000011101011010011;
    rom[9770] = 25'b0000000000011101011010010;
    rom[9771] = 25'b0000000000011101011010000;
    rom[9772] = 25'b0000000000011101011001111;
    rom[9773] = 25'b0000000000011101011001110;
    rom[9774] = 25'b0000000000011101011001101;
    rom[9775] = 25'b0000000000011101011001011;
    rom[9776] = 25'b0000000000011101011001010;
    rom[9777] = 25'b0000000000011101011001001;
    rom[9778] = 25'b0000000000011101011001000;
    rom[9779] = 25'b0000000000011101011000110;
    rom[9780] = 25'b0000000000011101011000101;
    rom[9781] = 25'b0000000000011101011000100;
    rom[9782] = 25'b0000000000011101011000010;
    rom[9783] = 25'b0000000000011101011000001;
    rom[9784] = 25'b0000000000011101010111111;
    rom[9785] = 25'b0000000000011101010111110;
    rom[9786] = 25'b0000000000011101010111100;
    rom[9787] = 25'b0000000000011101010111011;
    rom[9788] = 25'b0000000000011101010111001;
    rom[9789] = 25'b0000000000011101010111000;
    rom[9790] = 25'b0000000000011101010110110;
    rom[9791] = 25'b0000000000011101010110101;
    rom[9792] = 25'b0000000000011101010110011;
    rom[9793] = 25'b0000000000011101010110001;
    rom[9794] = 25'b0000000000011101010110000;
    rom[9795] = 25'b0000000000011101010101110;
    rom[9796] = 25'b0000000000011101010101100;
    rom[9797] = 25'b0000000000011101010101010;
    rom[9798] = 25'b0000000000011101010101001;
    rom[9799] = 25'b0000000000011101010100111;
    rom[9800] = 25'b0000000000011101010100101;
    rom[9801] = 25'b0000000000011101010100011;
    rom[9802] = 25'b0000000000011101010100001;
    rom[9803] = 25'b0000000000011101010011111;
    rom[9804] = 25'b0000000000011101010011110;
    rom[9805] = 25'b0000000000011101010011011;
    rom[9806] = 25'b0000000000011101010011010;
    rom[9807] = 25'b0000000000011101010011000;
    rom[9808] = 25'b0000000000011101010010101;
    rom[9809] = 25'b0000000000011101010010100;
    rom[9810] = 25'b0000000000011101010010010;
    rom[9811] = 25'b0000000000011101010001111;
    rom[9812] = 25'b0000000000011101010001101;
    rom[9813] = 25'b0000000000011101010001100;
    rom[9814] = 25'b0000000000011101010001010;
    rom[9815] = 25'b0000000000011101010000111;
    rom[9816] = 25'b0000000000011101010000101;
    rom[9817] = 25'b0000000000011101010000011;
    rom[9818] = 25'b0000000000011101010000001;
    rom[9819] = 25'b0000000000011101001111110;
    rom[9820] = 25'b0000000000011101001111100;
    rom[9821] = 25'b0000000000011101001111010;
    rom[9822] = 25'b0000000000011101001111000;
    rom[9823] = 25'b0000000000011101001110101;
    rom[9824] = 25'b0000000000011101001110010;
    rom[9825] = 25'b0000000000011101001110000;
    rom[9826] = 25'b0000000000011101001101110;
    rom[9827] = 25'b0000000000011101001101100;
    rom[9828] = 25'b0000000000011101001101001;
    rom[9829] = 25'b0000000000011101001100110;
    rom[9830] = 25'b0000000000011101001100100;
    rom[9831] = 25'b0000000000011101001100001;
    rom[9832] = 25'b0000000000011101001011111;
    rom[9833] = 25'b0000000000011101001011100;
    rom[9834] = 25'b0000000000011101001011010;
    rom[9835] = 25'b0000000000011101001010111;
    rom[9836] = 25'b0000000000011101001010100;
    rom[9837] = 25'b0000000000011101001010001;
    rom[9838] = 25'b0000000000011101001001111;
    rom[9839] = 25'b0000000000011101001001100;
    rom[9840] = 25'b0000000000011101001001001;
    rom[9841] = 25'b0000000000011101001000111;
    rom[9842] = 25'b0000000000011101001000100;
    rom[9843] = 25'b0000000000011101001000001;
    rom[9844] = 25'b0000000000011101000111111;
    rom[9845] = 25'b0000000000011101000111100;
    rom[9846] = 25'b0000000000011101000111001;
    rom[9847] = 25'b0000000000011101000110110;
    rom[9848] = 25'b0000000000011101000110011;
    rom[9849] = 25'b0000000000011101000110000;
    rom[9850] = 25'b0000000000011101000101101;
    rom[9851] = 25'b0000000000011101000101010;
    rom[9852] = 25'b0000000000011101000100111;
    rom[9853] = 25'b0000000000011101000100100;
    rom[9854] = 25'b0000000000011101000100001;
    rom[9855] = 25'b0000000000011101000011110;
    rom[9856] = 25'b0000000000011101000011011;
    rom[9857] = 25'b0000000000011101000010111;
    rom[9858] = 25'b0000000000011101000010100;
    rom[9859] = 25'b0000000000011101000010001;
    rom[9860] = 25'b0000000000011101000001110;
    rom[9861] = 25'b0000000000011101000001010;
    rom[9862] = 25'b0000000000011101000001000;
    rom[9863] = 25'b0000000000011101000000101;
    rom[9864] = 25'b0000000000011101000000001;
    rom[9865] = 25'b0000000000011100111111110;
    rom[9866] = 25'b0000000000011100111111010;
    rom[9867] = 25'b0000000000011100111110111;
    rom[9868] = 25'b0000000000011100111110011;
    rom[9869] = 25'b0000000000011100111110000;
    rom[9870] = 25'b0000000000011100111101101;
    rom[9871] = 25'b0000000000011100111101001;
    rom[9872] = 25'b0000000000011100111100110;
    rom[9873] = 25'b0000000000011100111100010;
    rom[9874] = 25'b0000000000011100111011110;
    rom[9875] = 25'b0000000000011100111011011;
    rom[9876] = 25'b0000000000011100111011000;
    rom[9877] = 25'b0000000000011100111010100;
    rom[9878] = 25'b0000000000011100111010000;
    rom[9879] = 25'b0000000000011100111001100;
    rom[9880] = 25'b0000000000011100111001001;
    rom[9881] = 25'b0000000000011100111000101;
    rom[9882] = 25'b0000000000011100111000001;
    rom[9883] = 25'b0000000000011100110111110;
    rom[9884] = 25'b0000000000011100110111010;
    rom[9885] = 25'b0000000000011100110110110;
    rom[9886] = 25'b0000000000011100110110010;
    rom[9887] = 25'b0000000000011100110101111;
    rom[9888] = 25'b0000000000011100110101011;
    rom[9889] = 25'b0000000000011100110100110;
    rom[9890] = 25'b0000000000011100110100011;
    rom[9891] = 25'b0000000000011100110011111;
    rom[9892] = 25'b0000000000011100110011011;
    rom[9893] = 25'b0000000000011100110010111;
    rom[9894] = 25'b0000000000011100110010011;
    rom[9895] = 25'b0000000000011100110001110;
    rom[9896] = 25'b0000000000011100110001011;
    rom[9897] = 25'b0000000000011100110000111;
    rom[9898] = 25'b0000000000011100110000011;
    rom[9899] = 25'b0000000000011100101111111;
    rom[9900] = 25'b0000000000011100101111010;
    rom[9901] = 25'b0000000000011100101110110;
    rom[9902] = 25'b0000000000011100101110010;
    rom[9903] = 25'b0000000000011100101101110;
    rom[9904] = 25'b0000000000011100101101001;
    rom[9905] = 25'b0000000000011100101100101;
    rom[9906] = 25'b0000000000011100101100001;
    rom[9907] = 25'b0000000000011100101011100;
    rom[9908] = 25'b0000000000011100101011000;
    rom[9909] = 25'b0000000000011100101010011;
    rom[9910] = 25'b0000000000011100101010000;
    rom[9911] = 25'b0000000000011100101001011;
    rom[9912] = 25'b0000000000011100101000111;
    rom[9913] = 25'b0000000000011100101000010;
    rom[9914] = 25'b0000000000011100100111110;
    rom[9915] = 25'b0000000000011100100111001;
    rom[9916] = 25'b0000000000011100100110101;
    rom[9917] = 25'b0000000000011100100110000;
    rom[9918] = 25'b0000000000011100100101011;
    rom[9919] = 25'b0000000000011100100100111;
    rom[9920] = 25'b0000000000011100100100010;
    rom[9921] = 25'b0000000000011100100011110;
    rom[9922] = 25'b0000000000011100100011000;
    rom[9923] = 25'b0000000000011100100010100;
    rom[9924] = 25'b0000000000011100100001111;
    rom[9925] = 25'b0000000000011100100001010;
    rom[9926] = 25'b0000000000011100100000110;
    rom[9927] = 25'b0000000000011100100000001;
    rom[9928] = 25'b0000000000011100011111100;
    rom[9929] = 25'b0000000000011100011111000;
    rom[9930] = 25'b0000000000011100011110010;
    rom[9931] = 25'b0000000000011100011101110;
    rom[9932] = 25'b0000000000011100011101001;
    rom[9933] = 25'b0000000000011100011100011;
    rom[9934] = 25'b0000000000011100011011111;
    rom[9935] = 25'b0000000000011100011011010;
    rom[9936] = 25'b0000000000011100011010100;
    rom[9937] = 25'b0000000000011100011001111;
    rom[9938] = 25'b0000000000011100011001011;
    rom[9939] = 25'b0000000000011100011000110;
    rom[9940] = 25'b0000000000011100011000000;
    rom[9941] = 25'b0000000000011100010111011;
    rom[9942] = 25'b0000000000011100010110110;
    rom[9943] = 25'b0000000000011100010110001;
    rom[9944] = 25'b0000000000011100010101011;
    rom[9945] = 25'b0000000000011100010100110;
    rom[9946] = 25'b0000000000011100010100001;
    rom[9947] = 25'b0000000000011100010011100;
    rom[9948] = 25'b0000000000011100010010110;
    rom[9949] = 25'b0000000000011100010010001;
    rom[9950] = 25'b0000000000011100010001100;
    rom[9951] = 25'b0000000000011100010000110;
    rom[9952] = 25'b0000000000011100010000001;
    rom[9953] = 25'b0000000000011100001111100;
    rom[9954] = 25'b0000000000011100001110110;
    rom[9955] = 25'b0000000000011100001110000;
    rom[9956] = 25'b0000000000011100001101011;
    rom[9957] = 25'b0000000000011100001100101;
    rom[9958] = 25'b0000000000011100001100000;
    rom[9959] = 25'b0000000000011100001011011;
    rom[9960] = 25'b0000000000011100001010101;
    rom[9961] = 25'b0000000000011100001001111;
    rom[9962] = 25'b0000000000011100001001001;
    rom[9963] = 25'b0000000000011100001000100;
    rom[9964] = 25'b0000000000011100000111110;
    rom[9965] = 25'b0000000000011100000111000;
    rom[9966] = 25'b0000000000011100000110010;
    rom[9967] = 25'b0000000000011100000101101;
    rom[9968] = 25'b0000000000011100000100111;
    rom[9969] = 25'b0000000000011100000100001;
    rom[9970] = 25'b0000000000011100000011011;
    rom[9971] = 25'b0000000000011100000010101;
    rom[9972] = 25'b0000000000011100000001111;
    rom[9973] = 25'b0000000000011100000001001;
    rom[9974] = 25'b0000000000011100000000011;
    rom[9975] = 25'b0000000000011011111111101;
    rom[9976] = 25'b0000000000011011111110111;
    rom[9977] = 25'b0000000000011011111110001;
    rom[9978] = 25'b0000000000011011111101011;
    rom[9979] = 25'b0000000000011011111100101;
    rom[9980] = 25'b0000000000011011111011111;
    rom[9981] = 25'b0000000000011011111011001;
    rom[9982] = 25'b0000000000011011111010011;
    rom[9983] = 25'b0000000000011011111001101;
    rom[9984] = 25'b0000000000011011111000111;
    rom[9985] = 25'b0000000000011011111000001;
    rom[9986] = 25'b0000000000011011110111010;
    rom[9987] = 25'b0000000000011011110110100;
    rom[9988] = 25'b0000000000011011110101101;
    rom[9989] = 25'b0000000000011011110100111;
    rom[9990] = 25'b0000000000011011110100001;
    rom[9991] = 25'b0000000000011011110011011;
    rom[9992] = 25'b0000000000011011110010100;
    rom[9993] = 25'b0000000000011011110001110;
    rom[9994] = 25'b0000000000011011110000111;
    rom[9995] = 25'b0000000000011011110000001;
    rom[9996] = 25'b0000000000011011101111011;
    rom[9997] = 25'b0000000000011011101110100;
    rom[9998] = 25'b0000000000011011101101101;
    rom[9999] = 25'b0000000000011011101100110;
    rom[10000] = 25'b0000000000011011101100000;
    rom[10001] = 25'b0000000000011011101011010;
    rom[10002] = 25'b0000000000011011101010011;
    rom[10003] = 25'b0000000000011011101001100;
    rom[10004] = 25'b0000000000011011101000110;
    rom[10005] = 25'b0000000000011011100111111;
    rom[10006] = 25'b0000000000011011100111000;
    rom[10007] = 25'b0000000000011011100110001;
    rom[10008] = 25'b0000000000011011100101011;
    rom[10009] = 25'b0000000000011011100100100;
    rom[10010] = 25'b0000000000011011100011100;
    rom[10011] = 25'b0000000000011011100010110;
    rom[10012] = 25'b0000000000011011100001111;
    rom[10013] = 25'b0000000000011011100001000;
    rom[10014] = 25'b0000000000011011100000001;
    rom[10015] = 25'b0000000000011011011111010;
    rom[10016] = 25'b0000000000011011011110011;
    rom[10017] = 25'b0000000000011011011101100;
    rom[10018] = 25'b0000000000011011011100101;
    rom[10019] = 25'b0000000000011011011011110;
    rom[10020] = 25'b0000000000011011011010111;
    rom[10021] = 25'b0000000000011011011001111;
    rom[10022] = 25'b0000000000011011011001001;
    rom[10023] = 25'b0000000000011011011000001;
    rom[10024] = 25'b0000000000011011010111011;
    rom[10025] = 25'b0000000000011011010110011;
    rom[10026] = 25'b0000000000011011010101100;
    rom[10027] = 25'b0000000000011011010100101;
    rom[10028] = 25'b0000000000011011010011101;
    rom[10029] = 25'b0000000000011011010010110;
    rom[10030] = 25'b0000000000011011010001110;
    rom[10031] = 25'b0000000000011011010000111;
    rom[10032] = 25'b0000000000011011010000000;
    rom[10033] = 25'b0000000000011011001111000;
    rom[10034] = 25'b0000000000011011001110001;
    rom[10035] = 25'b0000000000011011001101010;
    rom[10036] = 25'b0000000000011011001100010;
    rom[10037] = 25'b0000000000011011001011010;
    rom[10038] = 25'b0000000000011011001010011;
    rom[10039] = 25'b0000000000011011001001011;
    rom[10040] = 25'b0000000000011011001000100;
    rom[10041] = 25'b0000000000011011000111100;
    rom[10042] = 25'b0000000000011011000110101;
    rom[10043] = 25'b0000000000011011000101101;
    rom[10044] = 25'b0000000000011011000100101;
    rom[10045] = 25'b0000000000011011000011110;
    rom[10046] = 25'b0000000000011011000010101;
    rom[10047] = 25'b0000000000011011000001110;
    rom[10048] = 25'b0000000000011011000000110;
    rom[10049] = 25'b0000000000011010111111110;
    rom[10050] = 25'b0000000000011010111110111;
    rom[10051] = 25'b0000000000011010111101111;
    rom[10052] = 25'b0000000000011010111100110;
    rom[10053] = 25'b0000000000011010111011111;
    rom[10054] = 25'b0000000000011010111010111;
    rom[10055] = 25'b0000000000011010111001111;
    rom[10056] = 25'b0000000000011010111000111;
    rom[10057] = 25'b0000000000011010110111111;
    rom[10058] = 25'b0000000000011010110110111;
    rom[10059] = 25'b0000000000011010110101110;
    rom[10060] = 25'b0000000000011010110100111;
    rom[10061] = 25'b0000000000011010110011111;
    rom[10062] = 25'b0000000000011010110010110;
    rom[10063] = 25'b0000000000011010110001110;
    rom[10064] = 25'b0000000000011010110000110;
    rom[10065] = 25'b0000000000011010101111110;
    rom[10066] = 25'b0000000000011010101110110;
    rom[10067] = 25'b0000000000011010101101101;
    rom[10068] = 25'b0000000000011010101100101;
    rom[10069] = 25'b0000000000011010101011101;
    rom[10070] = 25'b0000000000011010101010100;
    rom[10071] = 25'b0000000000011010101001100;
    rom[10072] = 25'b0000000000011010101000011;
    rom[10073] = 25'b0000000000011010100111011;
    rom[10074] = 25'b0000000000011010100110010;
    rom[10075] = 25'b0000000000011010100101010;
    rom[10076] = 25'b0000000000011010100100010;
    rom[10077] = 25'b0000000000011010100011001;
    rom[10078] = 25'b0000000000011010100010001;
    rom[10079] = 25'b0000000000011010100001000;
    rom[10080] = 25'b0000000000011010100000000;
    rom[10081] = 25'b0000000000011010011110111;
    rom[10082] = 25'b0000000000011010011101110;
    rom[10083] = 25'b0000000000011010011100101;
    rom[10084] = 25'b0000000000011010011011100;
    rom[10085] = 25'b0000000000011010011010100;
    rom[10086] = 25'b0000000000011010011001011;
    rom[10087] = 25'b0000000000011010011000010;
    rom[10088] = 25'b0000000000011010010111001;
    rom[10089] = 25'b0000000000011010010110001;
    rom[10090] = 25'b0000000000011010010101000;
    rom[10091] = 25'b0000000000011010010011111;
    rom[10092] = 25'b0000000000011010010010110;
    rom[10093] = 25'b0000000000011010010001101;
    rom[10094] = 25'b0000000000011010010000100;
    rom[10095] = 25'b0000000000011010001111011;
    rom[10096] = 25'b0000000000011010001110010;
    rom[10097] = 25'b0000000000011010001101001;
    rom[10098] = 25'b0000000000011010001100000;
    rom[10099] = 25'b0000000000011010001010111;
    rom[10100] = 25'b0000000000011010001001110;
    rom[10101] = 25'b0000000000011010001000101;
    rom[10102] = 25'b0000000000011010000111100;
    rom[10103] = 25'b0000000000011010000110011;
    rom[10104] = 25'b0000000000011010000101001;
    rom[10105] = 25'b0000000000011010000100000;
    rom[10106] = 25'b0000000000011010000010111;
    rom[10107] = 25'b0000000000011010000001101;
    rom[10108] = 25'b0000000000011010000000100;
    rom[10109] = 25'b0000000000011001111111011;
    rom[10110] = 25'b0000000000011001111110010;
    rom[10111] = 25'b0000000000011001111101000;
    rom[10112] = 25'b0000000000011001111011110;
    rom[10113] = 25'b0000000000011001111010101;
    rom[10114] = 25'b0000000000011001111001100;
    rom[10115] = 25'b0000000000011001111000010;
    rom[10116] = 25'b0000000000011001110111001;
    rom[10117] = 25'b0000000000011001110101111;
    rom[10118] = 25'b0000000000011001110100110;
    rom[10119] = 25'b0000000000011001110011100;
    rom[10120] = 25'b0000000000011001110010010;
    rom[10121] = 25'b0000000000011001110001001;
    rom[10122] = 25'b0000000000011001110000000;
    rom[10123] = 25'b0000000000011001101110110;
    rom[10124] = 25'b0000000000011001101101100;
    rom[10125] = 25'b0000000000011001101100010;
    rom[10126] = 25'b0000000000011001101011001;
    rom[10127] = 25'b0000000000011001101001110;
    rom[10128] = 25'b0000000000011001101000100;
    rom[10129] = 25'b0000000000011001100111011;
    rom[10130] = 25'b0000000000011001100110001;
    rom[10131] = 25'b0000000000011001100100111;
    rom[10132] = 25'b0000000000011001100011101;
    rom[10133] = 25'b0000000000011001100010011;
    rom[10134] = 25'b0000000000011001100001001;
    rom[10135] = 25'b0000000000011001011111111;
    rom[10136] = 25'b0000000000011001011110101;
    rom[10137] = 25'b0000000000011001011101011;
    rom[10138] = 25'b0000000000011001011100001;
    rom[10139] = 25'b0000000000011001011010111;
    rom[10140] = 25'b0000000000011001011001101;
    rom[10141] = 25'b0000000000011001011000010;
    rom[10142] = 25'b0000000000011001010111001;
    rom[10143] = 25'b0000000000011001010101110;
    rom[10144] = 25'b0000000000011001010100100;
    rom[10145] = 25'b0000000000011001010011010;
    rom[10146] = 25'b0000000000011001010010000;
    rom[10147] = 25'b0000000000011001010000101;
    rom[10148] = 25'b0000000000011001001111011;
    rom[10149] = 25'b0000000000011001001110000;
    rom[10150] = 25'b0000000000011001001100110;
    rom[10151] = 25'b0000000000011001001011100;
    rom[10152] = 25'b0000000000011001001010010;
    rom[10153] = 25'b0000000000011001001000111;
    rom[10154] = 25'b0000000000011001000111101;
    rom[10155] = 25'b0000000000011001000110010;
    rom[10156] = 25'b0000000000011001000100111;
    rom[10157] = 25'b0000000000011001000011101;
    rom[10158] = 25'b0000000000011001000010010;
    rom[10159] = 25'b0000000000011001000001000;
    rom[10160] = 25'b0000000000011000111111101;
    rom[10161] = 25'b0000000000011000111110010;
    rom[10162] = 25'b0000000000011000111101000;
    rom[10163] = 25'b0000000000011000111011101;
    rom[10164] = 25'b0000000000011000111010010;
    rom[10165] = 25'b0000000000011000111000111;
    rom[10166] = 25'b0000000000011000110111101;
    rom[10167] = 25'b0000000000011000110110010;
    rom[10168] = 25'b0000000000011000110100111;
    rom[10169] = 25'b0000000000011000110011100;
    rom[10170] = 25'b0000000000011000110010001;
    rom[10171] = 25'b0000000000011000110000110;
    rom[10172] = 25'b0000000000011000101111011;
    rom[10173] = 25'b0000000000011000101110001;
    rom[10174] = 25'b0000000000011000101100110;
    rom[10175] = 25'b0000000000011000101011010;
    rom[10176] = 25'b0000000000011000101001111;
    rom[10177] = 25'b0000000000011000101000101;
    rom[10178] = 25'b0000000000011000100111010;
    rom[10179] = 25'b0000000000011000100101110;
    rom[10180] = 25'b0000000000011000100100011;
    rom[10181] = 25'b0000000000011000100011000;
    rom[10182] = 25'b0000000000011000100001101;
    rom[10183] = 25'b0000000000011000100000001;
    rom[10184] = 25'b0000000000011000011110110;
    rom[10185] = 25'b0000000000011000011101011;
    rom[10186] = 25'b0000000000011000011100000;
    rom[10187] = 25'b0000000000011000011010100;
    rom[10188] = 25'b0000000000011000011001001;
    rom[10189] = 25'b0000000000011000010111101;
    rom[10190] = 25'b0000000000011000010110010;
    rom[10191] = 25'b0000000000011000010100111;
    rom[10192] = 25'b0000000000011000010011011;
    rom[10193] = 25'b0000000000011000010010000;
    rom[10194] = 25'b0000000000011000010000100;
    rom[10195] = 25'b0000000000011000001111001;
    rom[10196] = 25'b0000000000011000001101110;
    rom[10197] = 25'b0000000000011000001100010;
    rom[10198] = 25'b0000000000011000001010110;
    rom[10199] = 25'b0000000000011000001001010;
    rom[10200] = 25'b0000000000011000000111110;
    rom[10201] = 25'b0000000000011000000110011;
    rom[10202] = 25'b0000000000011000000100111;
    rom[10203] = 25'b0000000000011000000011011;
    rom[10204] = 25'b0000000000011000000010000;
    rom[10205] = 25'b0000000000011000000000100;
    rom[10206] = 25'b0000000000010111111111000;
    rom[10207] = 25'b0000000000010111111101100;
    rom[10208] = 25'b0000000000010111111100000;
    rom[10209] = 25'b0000000000010111111010100;
    rom[10210] = 25'b0000000000010111111001000;
    rom[10211] = 25'b0000000000010111110111101;
    rom[10212] = 25'b0000000000010111110110001;
    rom[10213] = 25'b0000000000010111110100101;
    rom[10214] = 25'b0000000000010111110011001;
    rom[10215] = 25'b0000000000010111110001101;
    rom[10216] = 25'b0000000000010111110000001;
    rom[10217] = 25'b0000000000010111101110101;
    rom[10218] = 25'b0000000000010111101101001;
    rom[10219] = 25'b0000000000010111101011100;
    rom[10220] = 25'b0000000000010111101010000;
    rom[10221] = 25'b0000000000010111101000100;
    rom[10222] = 25'b0000000000010111100111000;
    rom[10223] = 25'b0000000000010111100101100;
    rom[10224] = 25'b0000000000010111100100000;
    rom[10225] = 25'b0000000000010111100010011;
    rom[10226] = 25'b0000000000010111100000111;
    rom[10227] = 25'b0000000000010111011111010;
    rom[10228] = 25'b0000000000010111011101110;
    rom[10229] = 25'b0000000000010111011100010;
    rom[10230] = 25'b0000000000010111011010101;
    rom[10231] = 25'b0000000000010111011001001;
    rom[10232] = 25'b0000000000010111010111100;
    rom[10233] = 25'b0000000000010111010110000;
    rom[10234] = 25'b0000000000010111010100100;
    rom[10235] = 25'b0000000000010111010010111;
    rom[10236] = 25'b0000000000010111010001010;
    rom[10237] = 25'b0000000000010111001111101;
    rom[10238] = 25'b0000000000010111001110001;
    rom[10239] = 25'b0000000000010111001100100;
    rom[10240] = 25'b0000000000010111001010111;
    rom[10241] = 25'b0000000000010111001001011;
    rom[10242] = 25'b0000000000010111000111110;
    rom[10243] = 25'b0000000000010111000110001;
    rom[10244] = 25'b0000000000010111000100101;
    rom[10245] = 25'b0000000000010111000011000;
    rom[10246] = 25'b0000000000010111000001011;
    rom[10247] = 25'b0000000000010110111111110;
    rom[10248] = 25'b0000000000010110111110001;
    rom[10249] = 25'b0000000000010110111100100;
    rom[10250] = 25'b0000000000010110111011000;
    rom[10251] = 25'b0000000000010110111001011;
    rom[10252] = 25'b0000000000010110110111101;
    rom[10253] = 25'b0000000000010110110110001;
    rom[10254] = 25'b0000000000010110110100011;
    rom[10255] = 25'b0000000000010110110010111;
    rom[10256] = 25'b0000000000010110110001001;
    rom[10257] = 25'b0000000000010110101111100;
    rom[10258] = 25'b0000000000010110101101111;
    rom[10259] = 25'b0000000000010110101100010;
    rom[10260] = 25'b0000000000010110101010101;
    rom[10261] = 25'b0000000000010110101000111;
    rom[10262] = 25'b0000000000010110100111011;
    rom[10263] = 25'b0000000000010110100101101;
    rom[10264] = 25'b0000000000010110100100000;
    rom[10265] = 25'b0000000000010110100010010;
    rom[10266] = 25'b0000000000010110100000101;
    rom[10267] = 25'b0000000000010110011111000;
    rom[10268] = 25'b0000000000010110011101011;
    rom[10269] = 25'b0000000000010110011011101;
    rom[10270] = 25'b0000000000010110011010000;
    rom[10271] = 25'b0000000000010110011000010;
    rom[10272] = 25'b0000000000010110010110100;
    rom[10273] = 25'b0000000000010110010100111;
    rom[10274] = 25'b0000000000010110010011001;
    rom[10275] = 25'b0000000000010110010001100;
    rom[10276] = 25'b0000000000010110001111110;
    rom[10277] = 25'b0000000000010110001110001;
    rom[10278] = 25'b0000000000010110001100011;
    rom[10279] = 25'b0000000000010110001010101;
    rom[10280] = 25'b0000000000010110001001000;
    rom[10281] = 25'b0000000000010110000111010;
    rom[10282] = 25'b0000000000010110000101100;
    rom[10283] = 25'b0000000000010110000011111;
    rom[10284] = 25'b0000000000010110000010001;
    rom[10285] = 25'b0000000000010110000000011;
    rom[10286] = 25'b0000000000010101111110101;
    rom[10287] = 25'b0000000000010101111101000;
    rom[10288] = 25'b0000000000010101111011001;
    rom[10289] = 25'b0000000000010101111001011;
    rom[10290] = 25'b0000000000010101110111110;
    rom[10291] = 25'b0000000000010101110110000;
    rom[10292] = 25'b0000000000010101110100001;
    rom[10293] = 25'b0000000000010101110010011;
    rom[10294] = 25'b0000000000010101110000110;
    rom[10295] = 25'b0000000000010101101110111;
    rom[10296] = 25'b0000000000010101101101001;
    rom[10297] = 25'b0000000000010101101011011;
    rom[10298] = 25'b0000000000010101101001101;
    rom[10299] = 25'b0000000000010101100111111;
    rom[10300] = 25'b0000000000010101100110001;
    rom[10301] = 25'b0000000000010101100100010;
    rom[10302] = 25'b0000000000010101100010100;
    rom[10303] = 25'b0000000000010101100000110;
    rom[10304] = 25'b0000000000010101011111000;
    rom[10305] = 25'b0000000000010101011101010;
    rom[10306] = 25'b0000000000010101011011011;
    rom[10307] = 25'b0000000000010101011001100;
    rom[10308] = 25'b0000000000010101010111110;
    rom[10309] = 25'b0000000000010101010110000;
    rom[10310] = 25'b0000000000010101010100001;
    rom[10311] = 25'b0000000000010101010010011;
    rom[10312] = 25'b0000000000010101010000100;
    rom[10313] = 25'b0000000000010101001110110;
    rom[10314] = 25'b0000000000010101001100111;
    rom[10315] = 25'b0000000000010101001011001;
    rom[10316] = 25'b0000000000010101001001010;
    rom[10317] = 25'b0000000000010101000111011;
    rom[10318] = 25'b0000000000010101000101101;
    rom[10319] = 25'b0000000000010101000011110;
    rom[10320] = 25'b0000000000010101000001111;
    rom[10321] = 25'b0000000000010101000000000;
    rom[10322] = 25'b0000000000010100111110010;
    rom[10323] = 25'b0000000000010100111100011;
    rom[10324] = 25'b0000000000010100111010100;
    rom[10325] = 25'b0000000000010100111000101;
    rom[10326] = 25'b0000000000010100110110110;
    rom[10327] = 25'b0000000000010100110101000;
    rom[10328] = 25'b0000000000010100110011001;
    rom[10329] = 25'b0000000000010100110001010;
    rom[10330] = 25'b0000000000010100101111011;
    rom[10331] = 25'b0000000000010100101101100;
    rom[10332] = 25'b0000000000010100101011101;
    rom[10333] = 25'b0000000000010100101001110;
    rom[10334] = 25'b0000000000010100100111111;
    rom[10335] = 25'b0000000000010100100110000;
    rom[10336] = 25'b0000000000010100100100000;
    rom[10337] = 25'b0000000000010100100010001;
    rom[10338] = 25'b0000000000010100100000010;
    rom[10339] = 25'b0000000000010100011110011;
    rom[10340] = 25'b0000000000010100011100100;
    rom[10341] = 25'b0000000000010100011010101;
    rom[10342] = 25'b0000000000010100011000101;
    rom[10343] = 25'b0000000000010100010110110;
    rom[10344] = 25'b0000000000010100010100111;
    rom[10345] = 25'b0000000000010100010011000;
    rom[10346] = 25'b0000000000010100010001000;
    rom[10347] = 25'b0000000000010100001111001;
    rom[10348] = 25'b0000000000010100001101001;
    rom[10349] = 25'b0000000000010100001011010;
    rom[10350] = 25'b0000000000010100001001011;
    rom[10351] = 25'b0000000000010100000111011;
    rom[10352] = 25'b0000000000010100000101011;
    rom[10353] = 25'b0000000000010100000011100;
    rom[10354] = 25'b0000000000010100000001101;
    rom[10355] = 25'b0000000000010011111111101;
    rom[10356] = 25'b0000000000010011111101101;
    rom[10357] = 25'b0000000000010011111011110;
    rom[10358] = 25'b0000000000010011111001110;
    rom[10359] = 25'b0000000000010011110111110;
    rom[10360] = 25'b0000000000010011110101111;
    rom[10361] = 25'b0000000000010011110011111;
    rom[10362] = 25'b0000000000010011110001111;
    rom[10363] = 25'b0000000000010011101111111;
    rom[10364] = 25'b0000000000010011101101111;
    rom[10365] = 25'b0000000000010011101011111;
    rom[10366] = 25'b0000000000010011101010000;
    rom[10367] = 25'b0000000000010011101000000;
    rom[10368] = 25'b0000000000010011100110000;
    rom[10369] = 25'b0000000000010011100100000;
    rom[10370] = 25'b0000000000010011100010000;
    rom[10371] = 25'b0000000000010011100000000;
    rom[10372] = 25'b0000000000010011011110000;
    rom[10373] = 25'b0000000000010011011100000;
    rom[10374] = 25'b0000000000010011011010000;
    rom[10375] = 25'b0000000000010011010111111;
    rom[10376] = 25'b0000000000010011010110000;
    rom[10377] = 25'b0000000000010011010011111;
    rom[10378] = 25'b0000000000010011010010000;
    rom[10379] = 25'b0000000000010011001111111;
    rom[10380] = 25'b0000000000010011001101111;
    rom[10381] = 25'b0000000000010011001011111;
    rom[10382] = 25'b0000000000010011001001111;
    rom[10383] = 25'b0000000000010011000111110;
    rom[10384] = 25'b0000000000010011000101110;
    rom[10385] = 25'b0000000000010011000011101;
    rom[10386] = 25'b0000000000010011000001101;
    rom[10387] = 25'b0000000000010010111111100;
    rom[10388] = 25'b0000000000010010111101101;
    rom[10389] = 25'b0000000000010010111011100;
    rom[10390] = 25'b0000000000010010111001100;
    rom[10391] = 25'b0000000000010010110111011;
    rom[10392] = 25'b0000000000010010110101010;
    rom[10393] = 25'b0000000000010010110011010;
    rom[10394] = 25'b0000000000010010110001001;
    rom[10395] = 25'b0000000000010010101111001;
    rom[10396] = 25'b0000000000010010101101001;
    rom[10397] = 25'b0000000000010010101010111;
    rom[10398] = 25'b0000000000010010101000111;
    rom[10399] = 25'b0000000000010010100110110;
    rom[10400] = 25'b0000000000010010100100101;
    rom[10401] = 25'b0000000000010010100010101;
    rom[10402] = 25'b0000000000010010100000100;
    rom[10403] = 25'b0000000000010010011110011;
    rom[10404] = 25'b0000000000010010011100011;
    rom[10405] = 25'b0000000000010010011010010;
    rom[10406] = 25'b0000000000010010011000001;
    rom[10407] = 25'b0000000000010010010110000;
    rom[10408] = 25'b0000000000010010010011111;
    rom[10409] = 25'b0000000000010010010001110;
    rom[10410] = 25'b0000000000010010001111101;
    rom[10411] = 25'b0000000000010010001101100;
    rom[10412] = 25'b0000000000010010001011011;
    rom[10413] = 25'b0000000000010010001001010;
    rom[10414] = 25'b0000000000010010000111001;
    rom[10415] = 25'b0000000000010010000101000;
    rom[10416] = 25'b0000000000010010000010111;
    rom[10417] = 25'b0000000000010010000000110;
    rom[10418] = 25'b0000000000010001111110100;
    rom[10419] = 25'b0000000000010001111100011;
    rom[10420] = 25'b0000000000010001111010010;
    rom[10421] = 25'b0000000000010001111000001;
    rom[10422] = 25'b0000000000010001110110000;
    rom[10423] = 25'b0000000000010001110011111;
    rom[10424] = 25'b0000000000010001110001101;
    rom[10425] = 25'b0000000000010001101111100;
    rom[10426] = 25'b0000000000010001101101010;
    rom[10427] = 25'b0000000000010001101011001;
    rom[10428] = 25'b0000000000010001101001000;
    rom[10429] = 25'b0000000000010001100110111;
    rom[10430] = 25'b0000000000010001100100101;
    rom[10431] = 25'b0000000000010001100010100;
    rom[10432] = 25'b0000000000010001100000010;
    rom[10433] = 25'b0000000000010001011110000;
    rom[10434] = 25'b0000000000010001011011111;
    rom[10435] = 25'b0000000000010001011001101;
    rom[10436] = 25'b0000000000010001010111011;
    rom[10437] = 25'b0000000000010001010101010;
    rom[10438] = 25'b0000000000010001010011000;
    rom[10439] = 25'b0000000000010001010000111;
    rom[10440] = 25'b0000000000010001001110101;
    rom[10441] = 25'b0000000000010001001100011;
    rom[10442] = 25'b0000000000010001001010001;
    rom[10443] = 25'b0000000000010001001000000;
    rom[10444] = 25'b0000000000010001000101110;
    rom[10445] = 25'b0000000000010001000011100;
    rom[10446] = 25'b0000000000010001000001010;
    rom[10447] = 25'b0000000000010000111111000;
    rom[10448] = 25'b0000000000010000111100111;
    rom[10449] = 25'b0000000000010000111010101;
    rom[10450] = 25'b0000000000010000111000011;
    rom[10451] = 25'b0000000000010000110110001;
    rom[10452] = 25'b0000000000010000110011111;
    rom[10453] = 25'b0000000000010000110001101;
    rom[10454] = 25'b0000000000010000101111011;
    rom[10455] = 25'b0000000000010000101101001;
    rom[10456] = 25'b0000000000010000101010111;
    rom[10457] = 25'b0000000000010000101000100;
    rom[10458] = 25'b0000000000010000100110010;
    rom[10459] = 25'b0000000000010000100100001;
    rom[10460] = 25'b0000000000010000100001111;
    rom[10461] = 25'b0000000000010000011111100;
    rom[10462] = 25'b0000000000010000011101010;
    rom[10463] = 25'b0000000000010000011010111;
    rom[10464] = 25'b0000000000010000011000101;
    rom[10465] = 25'b0000000000010000010110011;
    rom[10466] = 25'b0000000000010000010100001;
    rom[10467] = 25'b0000000000010000010001110;
    rom[10468] = 25'b0000000000010000001111100;
    rom[10469] = 25'b0000000000010000001101001;
    rom[10470] = 25'b0000000000010000001011000;
    rom[10471] = 25'b0000000000010000001000101;
    rom[10472] = 25'b0000000000010000000110010;
    rom[10473] = 25'b0000000000010000000100000;
    rom[10474] = 25'b0000000000010000000001110;
    rom[10475] = 25'b0000000000001111111111011;
    rom[10476] = 25'b0000000000001111111101000;
    rom[10477] = 25'b0000000000001111111010110;
    rom[10478] = 25'b0000000000001111111000011;
    rom[10479] = 25'b0000000000001111110110000;
    rom[10480] = 25'b0000000000001111110011110;
    rom[10481] = 25'b0000000000001111110001011;
    rom[10482] = 25'b0000000000001111101111000;
    rom[10483] = 25'b0000000000001111101100110;
    rom[10484] = 25'b0000000000001111101010011;
    rom[10485] = 25'b0000000000001111101000000;
    rom[10486] = 25'b0000000000001111100101101;
    rom[10487] = 25'b0000000000001111100011011;
    rom[10488] = 25'b0000000000001111100000111;
    rom[10489] = 25'b0000000000001111011110101;
    rom[10490] = 25'b0000000000001111011100010;
    rom[10491] = 25'b0000000000001111011001111;
    rom[10492] = 25'b0000000000001111010111100;
    rom[10493] = 25'b0000000000001111010101001;
    rom[10494] = 25'b0000000000001111010010110;
    rom[10495] = 25'b0000000000001111010000011;
    rom[10496] = 25'b0000000000001111001110000;
    rom[10497] = 25'b0000000000001111001011101;
    rom[10498] = 25'b0000000000001111001001010;
    rom[10499] = 25'b0000000000001111000110111;
    rom[10500] = 25'b0000000000001111000100100;
    rom[10501] = 25'b0000000000001111000010000;
    rom[10502] = 25'b0000000000001110111111101;
    rom[10503] = 25'b0000000000001110111101010;
    rom[10504] = 25'b0000000000001110111010111;
    rom[10505] = 25'b0000000000001110111000100;
    rom[10506] = 25'b0000000000001110110110000;
    rom[10507] = 25'b0000000000001110110011101;
    rom[10508] = 25'b0000000000001110110001010;
    rom[10509] = 25'b0000000000001110101110110;
    rom[10510] = 25'b0000000000001110101100011;
    rom[10511] = 25'b0000000000001110101001111;
    rom[10512] = 25'b0000000000001110100111100;
    rom[10513] = 25'b0000000000001110100101000;
    rom[10514] = 25'b0000000000001110100010101;
    rom[10515] = 25'b0000000000001110100000010;
    rom[10516] = 25'b0000000000001110011101110;
    rom[10517] = 25'b0000000000001110011011011;
    rom[10518] = 25'b0000000000001110011000111;
    rom[10519] = 25'b0000000000001110010110100;
    rom[10520] = 25'b0000000000001110010100000;
    rom[10521] = 25'b0000000000001110010001100;
    rom[10522] = 25'b0000000000001110001111001;
    rom[10523] = 25'b0000000000001110001100101;
    rom[10524] = 25'b0000000000001110001010001;
    rom[10525] = 25'b0000000000001110000111110;
    rom[10526] = 25'b0000000000001110000101010;
    rom[10527] = 25'b0000000000001110000010110;
    rom[10528] = 25'b0000000000001110000000010;
    rom[10529] = 25'b0000000000001101111101111;
    rom[10530] = 25'b0000000000001101111011011;
    rom[10531] = 25'b0000000000001101111000111;
    rom[10532] = 25'b0000000000001101110110011;
    rom[10533] = 25'b0000000000001101110011111;
    rom[10534] = 25'b0000000000001101110001011;
    rom[10535] = 25'b0000000000001101101110111;
    rom[10536] = 25'b0000000000001101101100011;
    rom[10537] = 25'b0000000000001101101001111;
    rom[10538] = 25'b0000000000001101100111011;
    rom[10539] = 25'b0000000000001101100100111;
    rom[10540] = 25'b0000000000001101100010011;
    rom[10541] = 25'b0000000000001101011111111;
    rom[10542] = 25'b0000000000001101011101011;
    rom[10543] = 25'b0000000000001101011010111;
    rom[10544] = 25'b0000000000001101011000010;
    rom[10545] = 25'b0000000000001101010101110;
    rom[10546] = 25'b0000000000001101010011010;
    rom[10547] = 25'b0000000000001101010000110;
    rom[10548] = 25'b0000000000001101001110010;
    rom[10549] = 25'b0000000000001101001011110;
    rom[10550] = 25'b0000000000001101001001001;
    rom[10551] = 25'b0000000000001101000110100;
    rom[10552] = 25'b0000000000001101000100000;
    rom[10553] = 25'b0000000000001101000001100;
    rom[10554] = 25'b0000000000001100111111000;
    rom[10555] = 25'b0000000000001100111100011;
    rom[10556] = 25'b0000000000001100111001111;
    rom[10557] = 25'b0000000000001100110111010;
    rom[10558] = 25'b0000000000001100110100110;
    rom[10559] = 25'b0000000000001100110010010;
    rom[10560] = 25'b0000000000001100101111101;
    rom[10561] = 25'b0000000000001100101101000;
    rom[10562] = 25'b0000000000001100101010100;
    rom[10563] = 25'b0000000000001100100111111;
    rom[10564] = 25'b0000000000001100100101010;
    rom[10565] = 25'b0000000000001100100010110;
    rom[10566] = 25'b0000000000001100100000001;
    rom[10567] = 25'b0000000000001100011101100;
    rom[10568] = 25'b0000000000001100011011000;
    rom[10569] = 25'b0000000000001100011000011;
    rom[10570] = 25'b0000000000001100010101110;
    rom[10571] = 25'b0000000000001100010011010;
    rom[10572] = 25'b0000000000001100010000101;
    rom[10573] = 25'b0000000000001100001110000;
    rom[10574] = 25'b0000000000001100001011011;
    rom[10575] = 25'b0000000000001100001000110;
    rom[10576] = 25'b0000000000001100000110001;
    rom[10577] = 25'b0000000000001100000011100;
    rom[10578] = 25'b0000000000001100000000111;
    rom[10579] = 25'b0000000000001011111110010;
    rom[10580] = 25'b0000000000001011111011101;
    rom[10581] = 25'b0000000000001011111001000;
    rom[10582] = 25'b0000000000001011110110011;
    rom[10583] = 25'b0000000000001011110011110;
    rom[10584] = 25'b0000000000001011110001001;
    rom[10585] = 25'b0000000000001011101110100;
    rom[10586] = 25'b0000000000001011101011111;
    rom[10587] = 25'b0000000000001011101001010;
    rom[10588] = 25'b0000000000001011100110100;
    rom[10589] = 25'b0000000000001011100011111;
    rom[10590] = 25'b0000000000001011100001010;
    rom[10591] = 25'b0000000000001011011110101;
    rom[10592] = 25'b0000000000001011011100000;
    rom[10593] = 25'b0000000000001011011001010;
    rom[10594] = 25'b0000000000001011010110101;
    rom[10595] = 25'b0000000000001011010100000;
    rom[10596] = 25'b0000000000001011010001010;
    rom[10597] = 25'b0000000000001011001110101;
    rom[10598] = 25'b0000000000001011001011111;
    rom[10599] = 25'b0000000000001011001001011;
    rom[10600] = 25'b0000000000001011000110101;
    rom[10601] = 25'b0000000000001011000011111;
    rom[10602] = 25'b0000000000001011000001010;
    rom[10603] = 25'b0000000000001010111110101;
    rom[10604] = 25'b0000000000001010111011111;
    rom[10605] = 25'b0000000000001010111001001;
    rom[10606] = 25'b0000000000001010110110100;
    rom[10607] = 25'b0000000000001010110011110;
    rom[10608] = 25'b0000000000001010110001000;
    rom[10609] = 25'b0000000000001010101110011;
    rom[10610] = 25'b0000000000001010101011101;
    rom[10611] = 25'b0000000000001010101000111;
    rom[10612] = 25'b0000000000001010100110010;
    rom[10613] = 25'b0000000000001010100011100;
    rom[10614] = 25'b0000000000001010100000110;
    rom[10615] = 25'b0000000000001010011110001;
    rom[10616] = 25'b0000000000001010011011011;
    rom[10617] = 25'b0000000000001010011000101;
    rom[10618] = 25'b0000000000001010010101111;
    rom[10619] = 25'b0000000000001010010011001;
    rom[10620] = 25'b0000000000001010010000100;
    rom[10621] = 25'b0000000000001010001101110;
    rom[10622] = 25'b0000000000001010001011000;
    rom[10623] = 25'b0000000000001010001000010;
    rom[10624] = 25'b0000000000001010000101011;
    rom[10625] = 25'b0000000000001010000010110;
    rom[10626] = 25'b0000000000001001111111111;
    rom[10627] = 25'b0000000000001001111101010;
    rom[10628] = 25'b0000000000001001111010011;
    rom[10629] = 25'b0000000000001001110111110;
    rom[10630] = 25'b0000000000001001110100111;
    rom[10631] = 25'b0000000000001001110010010;
    rom[10632] = 25'b0000000000001001101111011;
    rom[10633] = 25'b0000000000001001101100101;
    rom[10634] = 25'b0000000000001001101001111;
    rom[10635] = 25'b0000000000001001100111001;
    rom[10636] = 25'b0000000000001001100100010;
    rom[10637] = 25'b0000000000001001100001101;
    rom[10638] = 25'b0000000000001001011110110;
    rom[10639] = 25'b0000000000001001011100000;
    rom[10640] = 25'b0000000000001001011001001;
    rom[10641] = 25'b0000000000001001010110011;
    rom[10642] = 25'b0000000000001001010011100;
    rom[10643] = 25'b0000000000001001010000110;
    rom[10644] = 25'b0000000000001001001110000;
    rom[10645] = 25'b0000000000001001001011001;
    rom[10646] = 25'b0000000000001001001000011;
    rom[10647] = 25'b0000000000001001000101100;
    rom[10648] = 25'b0000000000001001000010110;
    rom[10649] = 25'b0000000000001001000000000;
    rom[10650] = 25'b0000000000001000111101001;
    rom[10651] = 25'b0000000000001000111010011;
    rom[10652] = 25'b0000000000001000110111100;
    rom[10653] = 25'b0000000000001000110100101;
    rom[10654] = 25'b0000000000001000110001111;
    rom[10655] = 25'b0000000000001000101111000;
    rom[10656] = 25'b0000000000001000101100001;
    rom[10657] = 25'b0000000000001000101001011;
    rom[10658] = 25'b0000000000001000100110100;
    rom[10659] = 25'b0000000000001000100011101;
    rom[10660] = 25'b0000000000001000100000111;
    rom[10661] = 25'b0000000000001000011110000;
    rom[10662] = 25'b0000000000001000011011001;
    rom[10663] = 25'b0000000000001000011000010;
    rom[10664] = 25'b0000000000001000010101100;
    rom[10665] = 25'b0000000000001000010010101;
    rom[10666] = 25'b0000000000001000001111101;
    rom[10667] = 25'b0000000000001000001100111;
    rom[10668] = 25'b0000000000001000001010000;
    rom[10669] = 25'b0000000000001000000111001;
    rom[10670] = 25'b0000000000001000000100010;
    rom[10671] = 25'b0000000000001000000001011;
    rom[10672] = 25'b0000000000000111111110100;
    rom[10673] = 25'b0000000000000111111011101;
    rom[10674] = 25'b0000000000000111111000110;
    rom[10675] = 25'b0000000000000111110101111;
    rom[10676] = 25'b0000000000000111110011000;
    rom[10677] = 25'b0000000000000111110000001;
    rom[10678] = 25'b0000000000000111101101010;
    rom[10679] = 25'b0000000000000111101010011;
    rom[10680] = 25'b0000000000000111100111011;
    rom[10681] = 25'b0000000000000111100100100;
    rom[10682] = 25'b0000000000000111100001101;
    rom[10683] = 25'b0000000000000111011110110;
    rom[10684] = 25'b0000000000000111011011111;
    rom[10685] = 25'b0000000000000111011000111;
    rom[10686] = 25'b0000000000000111010110000;
    rom[10687] = 25'b0000000000000111010011000;
    rom[10688] = 25'b0000000000000111010000001;
    rom[10689] = 25'b0000000000000111001101010;
    rom[10690] = 25'b0000000000000111001010010;
    rom[10691] = 25'b0000000000000111000111011;
    rom[10692] = 25'b0000000000000111000100100;
    rom[10693] = 25'b0000000000000111000001100;
    rom[10694] = 25'b0000000000000110111110101;
    rom[10695] = 25'b0000000000000110111011101;
    rom[10696] = 25'b0000000000000110111000110;
    rom[10697] = 25'b0000000000000110110101111;
    rom[10698] = 25'b0000000000000110110010111;
    rom[10699] = 25'b0000000000000110110000000;
    rom[10700] = 25'b0000000000000110101101000;
    rom[10701] = 25'b0000000000000110101010000;
    rom[10702] = 25'b0000000000000110100111001;
    rom[10703] = 25'b0000000000000110100100001;
    rom[10704] = 25'b0000000000000110100001001;
    rom[10705] = 25'b0000000000000110011110010;
    rom[10706] = 25'b0000000000000110011011010;
    rom[10707] = 25'b0000000000000110011000010;
    rom[10708] = 25'b0000000000000110010101011;
    rom[10709] = 25'b0000000000000110010010011;
    rom[10710] = 25'b0000000000000110001111011;
    rom[10711] = 25'b0000000000000110001100011;
    rom[10712] = 25'b0000000000000110001001011;
    rom[10713] = 25'b0000000000000110000110011;
    rom[10714] = 25'b0000000000000110000011011;
    rom[10715] = 25'b0000000000000110000000011;
    rom[10716] = 25'b0000000000000101111101011;
    rom[10717] = 25'b0000000000000101111010011;
    rom[10718] = 25'b0000000000000101110111100;
    rom[10719] = 25'b0000000000000101110100100;
    rom[10720] = 25'b0000000000000101110001100;
    rom[10721] = 25'b0000000000000101101110100;
    rom[10722] = 25'b0000000000000101101011100;
    rom[10723] = 25'b0000000000000101101000100;
    rom[10724] = 25'b0000000000000101100101100;
    rom[10725] = 25'b0000000000000101100010011;
    rom[10726] = 25'b0000000000000101011111100;
    rom[10727] = 25'b0000000000000101011100100;
    rom[10728] = 25'b0000000000000101011001011;
    rom[10729] = 25'b0000000000000101010110011;
    rom[10730] = 25'b0000000000000101010011011;
    rom[10731] = 25'b0000000000000101010000011;
    rom[10732] = 25'b0000000000000101001101011;
    rom[10733] = 25'b0000000000000101001010011;
    rom[10734] = 25'b0000000000000101000111010;
    rom[10735] = 25'b0000000000000101000100010;
    rom[10736] = 25'b0000000000000101000001010;
    rom[10737] = 25'b0000000000000100111110001;
    rom[10738] = 25'b0000000000000100111011001;
    rom[10739] = 25'b0000000000000100111000000;
    rom[10740] = 25'b0000000000000100110101000;
    rom[10741] = 25'b0000000000000100110010000;
    rom[10742] = 25'b0000000000000100101110111;
    rom[10743] = 25'b0000000000000100101011111;
    rom[10744] = 25'b0000000000000100101000111;
    rom[10745] = 25'b0000000000000100100101110;
    rom[10746] = 25'b0000000000000100100010101;
    rom[10747] = 25'b0000000000000100011111101;
    rom[10748] = 25'b0000000000000100011100101;
    rom[10749] = 25'b0000000000000100011001100;
    rom[10750] = 25'b0000000000000100010110011;
    rom[10751] = 25'b0000000000000100010011011;
    rom[10752] = 25'b0000000000000100010000010;
    rom[10753] = 25'b0000000000000100001101001;
    rom[10754] = 25'b0000000000000100001010001;
    rom[10755] = 25'b0000000000000100000111000;
    rom[10756] = 25'b0000000000000100000011111;
    rom[10757] = 25'b0000000000000100000000111;
    rom[10758] = 25'b0000000000000011111101110;
    rom[10759] = 25'b0000000000000011111010101;
    rom[10760] = 25'b0000000000000011110111101;
    rom[10761] = 25'b0000000000000011110100100;
    rom[10762] = 25'b0000000000000011110001011;
    rom[10763] = 25'b0000000000000011101110010;
    rom[10764] = 25'b0000000000000011101011001;
    rom[10765] = 25'b0000000000000011101000001;
    rom[10766] = 25'b0000000000000011100100111;
    rom[10767] = 25'b0000000000000011100001111;
    rom[10768] = 25'b0000000000000011011110110;
    rom[10769] = 25'b0000000000000011011011101;
    rom[10770] = 25'b0000000000000011011000100;
    rom[10771] = 25'b0000000000000011010101011;
    rom[10772] = 25'b0000000000000011010010010;
    rom[10773] = 25'b0000000000000011001111001;
    rom[10774] = 25'b0000000000000011001100000;
    rom[10775] = 25'b0000000000000011001000111;
    rom[10776] = 25'b0000000000000011000101110;
    rom[10777] = 25'b0000000000000011000010100;
    rom[10778] = 25'b0000000000000010111111100;
    rom[10779] = 25'b0000000000000010111100010;
    rom[10780] = 25'b0000000000000010111001010;
    rom[10781] = 25'b0000000000000010110110000;
    rom[10782] = 25'b0000000000000010110010111;
    rom[10783] = 25'b0000000000000010101111110;
    rom[10784] = 25'b0000000000000010101100101;
    rom[10785] = 25'b0000000000000010101001011;
    rom[10786] = 25'b0000000000000010100110010;
    rom[10787] = 25'b0000000000000010100011001;
    rom[10788] = 25'b0000000000000010100000000;
    rom[10789] = 25'b0000000000000010011100111;
    rom[10790] = 25'b0000000000000010011001101;
    rom[10791] = 25'b0000000000000010010110100;
    rom[10792] = 25'b0000000000000010010011010;
    rom[10793] = 25'b0000000000000010010000001;
    rom[10794] = 25'b0000000000000010001101000;
    rom[10795] = 25'b0000000000000010001001110;
    rom[10796] = 25'b0000000000000010000110101;
    rom[10797] = 25'b0000000000000010000011011;
    rom[10798] = 25'b0000000000000010000000010;
    rom[10799] = 25'b0000000000000001111101001;
    rom[10800] = 25'b0000000000000001111001110;
    rom[10801] = 25'b0000000000000001110110101;
    rom[10802] = 25'b0000000000000001110011100;
    rom[10803] = 25'b0000000000000001110000010;
    rom[10804] = 25'b0000000000000001101101001;
    rom[10805] = 25'b0000000000000001101001111;
    rom[10806] = 25'b0000000000000001100110101;
    rom[10807] = 25'b0000000000000001100011100;
    rom[10808] = 25'b0000000000000001100000010;
    rom[10809] = 25'b0000000000000001011101000;
    rom[10810] = 25'b0000000000000001011001111;
    rom[10811] = 25'b0000000000000001010110101;
    rom[10812] = 25'b0000000000000001010011011;
    rom[10813] = 25'b0000000000000001010000001;
    rom[10814] = 25'b0000000000000001001101000;
    rom[10815] = 25'b0000000000000001001001110;
    rom[10816] = 25'b0000000000000001000110100;
    rom[10817] = 25'b0000000000000001000011010;
    rom[10818] = 25'b0000000000000001000000001;
    rom[10819] = 25'b0000000000000000111100111;
    rom[10820] = 25'b0000000000000000111001101;
    rom[10821] = 25'b0000000000000000110110011;
    rom[10822] = 25'b0000000000000000110011001;
    rom[10823] = 25'b0000000000000000110000000;
    rom[10824] = 25'b0000000000000000101100101;
    rom[10825] = 25'b0000000000000000101001011;
    rom[10826] = 25'b0000000000000000100110001;
    rom[10827] = 25'b0000000000000000100011000;
    rom[10828] = 25'b0000000000000000011111110;
    rom[10829] = 25'b0000000000000000011100011;
    rom[10830] = 25'b0000000000000000011001001;
    rom[10831] = 25'b0000000000000000010101111;
    rom[10832] = 25'b0000000000000000010010101;
    rom[10833] = 25'b0000000000000000001111100;
    rom[10834] = 25'b0000000000000000001100001;
    rom[10835] = 25'b0000000000000000001000111;
    rom[10836] = 25'b0000000000000000000101101;
    rom[10837] = 25'b0000000000000000000010011;
    rom[10838] = 25'b1111111111111111111111010;
    rom[10839] = 25'b1111111111111111111011111;
    rom[10840] = 25'b1111111111111111111000100;
    rom[10841] = 25'b1111111111111111110101010;
    rom[10842] = 25'b1111111111111111110010000;
    rom[10843] = 25'b1111111111111111101110110;
    rom[10844] = 25'b1111111111111111101011100;
    rom[10845] = 25'b1111111111111111101000010;
    rom[10846] = 25'b1111111111111111100100111;
    rom[10847] = 25'b1111111111111111100001101;
    rom[10848] = 25'b1111111111111111011110011;
    rom[10849] = 25'b1111111111111111011011000;
    rom[10850] = 25'b1111111111111111010111110;
    rom[10851] = 25'b1111111111111111010100011;
    rom[10852] = 25'b1111111111111111010001001;
    rom[10853] = 25'b1111111111111111001101110;
    rom[10854] = 25'b1111111111111111001010100;
    rom[10855] = 25'b1111111111111111000111010;
    rom[10856] = 25'b1111111111111111000011111;
    rom[10857] = 25'b1111111111111111000000101;
    rom[10858] = 25'b1111111111111110111101010;
    rom[10859] = 25'b1111111111111110111010000;
    rom[10860] = 25'b1111111111111110110110101;
    rom[10861] = 25'b1111111111111110110011011;
    rom[10862] = 25'b1111111111111110110000000;
    rom[10863] = 25'b1111111111111110101100101;
    rom[10864] = 25'b1111111111111110101001011;
    rom[10865] = 25'b1111111111111110100110000;
    rom[10866] = 25'b1111111111111110100010101;
    rom[10867] = 25'b1111111111111110011111011;
    rom[10868] = 25'b1111111111111110011100000;
    rom[10869] = 25'b1111111111111110011000101;
    rom[10870] = 25'b1111111111111110010101011;
    rom[10871] = 25'b1111111111111110010010000;
    rom[10872] = 25'b1111111111111110001110101;
    rom[10873] = 25'b1111111111111110001011010;
    rom[10874] = 25'b1111111111111110000111111;
    rom[10875] = 25'b1111111111111110000100101;
    rom[10876] = 25'b1111111111111110000001010;
    rom[10877] = 25'b1111111111111101111110000;
    rom[10878] = 25'b1111111111111101111010101;
    rom[10879] = 25'b1111111111111101110111010;
    rom[10880] = 25'b1111111111111101110011111;
    rom[10881] = 25'b1111111111111101110000100;
    rom[10882] = 25'b1111111111111101101101001;
    rom[10883] = 25'b1111111111111101101001110;
    rom[10884] = 25'b1111111111111101100110011;
    rom[10885] = 25'b1111111111111101100011000;
    rom[10886] = 25'b1111111111111101011111101;
    rom[10887] = 25'b1111111111111101011100011;
    rom[10888] = 25'b1111111111111101011000111;
    rom[10889] = 25'b1111111111111101010101100;
    rom[10890] = 25'b1111111111111101010010001;
    rom[10891] = 25'b1111111111111101001110110;
    rom[10892] = 25'b1111111111111101001011011;
    rom[10893] = 25'b1111111111111101001000000;
    rom[10894] = 25'b1111111111111101000100101;
    rom[10895] = 25'b1111111111111101000001010;
    rom[10896] = 25'b1111111111111100111101111;
    rom[10897] = 25'b1111111111111100111010011;
    rom[10898] = 25'b1111111111111100110111000;
    rom[10899] = 25'b1111111111111100110011110;
    rom[10900] = 25'b1111111111111100110000010;
    rom[10901] = 25'b1111111111111100101100111;
    rom[10902] = 25'b1111111111111100101001011;
    rom[10903] = 25'b1111111111111100100110001;
    rom[10904] = 25'b1111111111111100100010101;
    rom[10905] = 25'b1111111111111100011111010;
    rom[10906] = 25'b1111111111111100011011110;
    rom[10907] = 25'b1111111111111100011000011;
    rom[10908] = 25'b1111111111111100010101000;
    rom[10909] = 25'b1111111111111100010001101;
    rom[10910] = 25'b1111111111111100001110001;
    rom[10911] = 25'b1111111111111100001010110;
    rom[10912] = 25'b1111111111111100000111011;
    rom[10913] = 25'b1111111111111100000011111;
    rom[10914] = 25'b1111111111111100000000100;
    rom[10915] = 25'b1111111111111011111101001;
    rom[10916] = 25'b1111111111111011111001101;
    rom[10917] = 25'b1111111111111011110110010;
    rom[10918] = 25'b1111111111111011110010110;
    rom[10919] = 25'b1111111111111011101111011;
    rom[10920] = 25'b1111111111111011101011111;
    rom[10921] = 25'b1111111111111011101000011;
    rom[10922] = 25'b1111111111111011100101001;
    rom[10923] = 25'b1111111111111011100001101;
    rom[10924] = 25'b1111111111111011011110001;
    rom[10925] = 25'b1111111111111011011010110;
    rom[10926] = 25'b1111111111111011010111010;
    rom[10927] = 25'b1111111111111011010011110;
    rom[10928] = 25'b1111111111111011010000011;
    rom[10929] = 25'b1111111111111011001100111;
    rom[10930] = 25'b1111111111111011001001011;
    rom[10931] = 25'b1111111111111011000110000;
    rom[10932] = 25'b1111111111111011000010100;
    rom[10933] = 25'b1111111111111010111111000;
    rom[10934] = 25'b1111111111111010111011101;
    rom[10935] = 25'b1111111111111010111000001;
    rom[10936] = 25'b1111111111111010110100110;
    rom[10937] = 25'b1111111111111010110001010;
    rom[10938] = 25'b1111111111111010101101110;
    rom[10939] = 25'b1111111111111010101010011;
    rom[10940] = 25'b1111111111111010100110110;
    rom[10941] = 25'b1111111111111010100011011;
    rom[10942] = 25'b1111111111111010011111111;
    rom[10943] = 25'b1111111111111010011100011;
    rom[10944] = 25'b1111111111111010011001000;
    rom[10945] = 25'b1111111111111010010101011;
    rom[10946] = 25'b1111111111111010010010000;
    rom[10947] = 25'b1111111111111010001110100;
    rom[10948] = 25'b1111111111111010001011000;
    rom[10949] = 25'b1111111111111010000111100;
    rom[10950] = 25'b1111111111111010000100000;
    rom[10951] = 25'b1111111111111010000000100;
    rom[10952] = 25'b1111111111111001111101000;
    rom[10953] = 25'b1111111111111001111001100;
    rom[10954] = 25'b1111111111111001110110000;
    rom[10955] = 25'b1111111111111001110010101;
    rom[10956] = 25'b1111111111111001101111000;
    rom[10957] = 25'b1111111111111001101011101;
    rom[10958] = 25'b1111111111111001101000000;
    rom[10959] = 25'b1111111111111001100100101;
    rom[10960] = 25'b1111111111111001100001000;
    rom[10961] = 25'b1111111111111001011101100;
    rom[10962] = 25'b1111111111111001011010000;
    rom[10963] = 25'b1111111111111001010110100;
    rom[10964] = 25'b1111111111111001010011000;
    rom[10965] = 25'b1111111111111001001111100;
    rom[10966] = 25'b1111111111111001001011111;
    rom[10967] = 25'b1111111111111001001000100;
    rom[10968] = 25'b1111111111111001000100111;
    rom[10969] = 25'b1111111111111001000001011;
    rom[10970] = 25'b1111111111111000111101111;
    rom[10971] = 25'b1111111111111000111010011;
    rom[10972] = 25'b1111111111111000110110110;
    rom[10973] = 25'b1111111111111000110011010;
    rom[10974] = 25'b1111111111111000101111110;
    rom[10975] = 25'b1111111111111000101100010;
    rom[10976] = 25'b1111111111111000101000110;
    rom[10977] = 25'b1111111111111000100101001;
    rom[10978] = 25'b1111111111111000100001101;
    rom[10979] = 25'b1111111111111000011110000;
    rom[10980] = 25'b1111111111111000011010100;
    rom[10981] = 25'b1111111111111000010111000;
    rom[10982] = 25'b1111111111111000010011100;
    rom[10983] = 25'b1111111111111000010000000;
    rom[10984] = 25'b1111111111111000001100011;
    rom[10985] = 25'b1111111111111000001000111;
    rom[10986] = 25'b1111111111111000000101011;
    rom[10987] = 25'b1111111111111000000001110;
    rom[10988] = 25'b1111111111110111111110010;
    rom[10989] = 25'b1111111111110111111010101;
    rom[10990] = 25'b1111111111110111110111000;
    rom[10991] = 25'b1111111111110111110011100;
    rom[10992] = 25'b1111111111110111101111111;
    rom[10993] = 25'b1111111111110111101100011;
    rom[10994] = 25'b1111111111110111101000111;
    rom[10995] = 25'b1111111111110111100101010;
    rom[10996] = 25'b1111111111110111100001110;
    rom[10997] = 25'b1111111111110111011110001;
    rom[10998] = 25'b1111111111110111011010100;
    rom[10999] = 25'b1111111111110111010111000;
    rom[11000] = 25'b1111111111110111010011100;
    rom[11001] = 25'b1111111111110111001111111;
    rom[11002] = 25'b1111111111110111001100010;
    rom[11003] = 25'b1111111111110111001000110;
    rom[11004] = 25'b1111111111110111000101001;
    rom[11005] = 25'b1111111111110111000001100;
    rom[11006] = 25'b1111111111110110111110000;
    rom[11007] = 25'b1111111111110110111010011;
    rom[11008] = 25'b1111111111110110110110110;
    rom[11009] = 25'b1111111111110110110011010;
    rom[11010] = 25'b1111111111110110101111101;
    rom[11011] = 25'b1111111111110110101100000;
    rom[11012] = 25'b1111111111110110101000100;
    rom[11013] = 25'b1111111111110110100100111;
    rom[11014] = 25'b1111111111110110100001010;
    rom[11015] = 25'b1111111111110110011101101;
    rom[11016] = 25'b1111111111110110011010001;
    rom[11017] = 25'b1111111111110110010110100;
    rom[11018] = 25'b1111111111110110010010111;
    rom[11019] = 25'b1111111111110110001111010;
    rom[11020] = 25'b1111111111110110001011110;
    rom[11021] = 25'b1111111111110110001000001;
    rom[11022] = 25'b1111111111110110000100100;
    rom[11023] = 25'b1111111111110110000000111;
    rom[11024] = 25'b1111111111110101111101010;
    rom[11025] = 25'b1111111111110101111001110;
    rom[11026] = 25'b1111111111110101110110000;
    rom[11027] = 25'b1111111111110101110010011;
    rom[11028] = 25'b1111111111110101101110111;
    rom[11029] = 25'b1111111111110101101011010;
    rom[11030] = 25'b1111111111110101100111101;
    rom[11031] = 25'b1111111111110101100100000;
    rom[11032] = 25'b1111111111110101100000011;
    rom[11033] = 25'b1111111111110101011100110;
    rom[11034] = 25'b1111111111110101011001001;
    rom[11035] = 25'b1111111111110101010101100;
    rom[11036] = 25'b1111111111110101010001111;
    rom[11037] = 25'b1111111111110101001110010;
    rom[11038] = 25'b1111111111110101001010101;
    rom[11039] = 25'b1111111111110101000111000;
    rom[11040] = 25'b1111111111110101000011011;
    rom[11041] = 25'b1111111111110100111111110;
    rom[11042] = 25'b1111111111110100111100001;
    rom[11043] = 25'b1111111111110100111000100;
    rom[11044] = 25'b1111111111110100110100111;
    rom[11045] = 25'b1111111111110100110001010;
    rom[11046] = 25'b1111111111110100101101101;
    rom[11047] = 25'b1111111111110100101010000;
    rom[11048] = 25'b1111111111110100100110010;
    rom[11049] = 25'b1111111111110100100010101;
    rom[11050] = 25'b1111111111110100011111000;
    rom[11051] = 25'b1111111111110100011011011;
    rom[11052] = 25'b1111111111110100010111110;
    rom[11053] = 25'b1111111111110100010100001;
    rom[11054] = 25'b1111111111110100010000100;
    rom[11055] = 25'b1111111111110100001100110;
    rom[11056] = 25'b1111111111110100001001001;
    rom[11057] = 25'b1111111111110100000101100;
    rom[11058] = 25'b1111111111110100000001111;
    rom[11059] = 25'b1111111111110011111110010;
    rom[11060] = 25'b1111111111110011111010100;
    rom[11061] = 25'b1111111111110011110110111;
    rom[11062] = 25'b1111111111110011110011010;
    rom[11063] = 25'b1111111111110011101111101;
    rom[11064] = 25'b1111111111110011101100000;
    rom[11065] = 25'b1111111111110011101000010;
    rom[11066] = 25'b1111111111110011100100100;
    rom[11067] = 25'b1111111111110011100000111;
    rom[11068] = 25'b1111111111110011011101010;
    rom[11069] = 25'b1111111111110011011001101;
    rom[11070] = 25'b1111111111110011010101111;
    rom[11071] = 25'b1111111111110011010010010;
    rom[11072] = 25'b1111111111110011001110101;
    rom[11073] = 25'b1111111111110011001010111;
    rom[11074] = 25'b1111111111110011000111010;
    rom[11075] = 25'b1111111111110011000011101;
    rom[11076] = 25'b1111111111110010111111111;
    rom[11077] = 25'b1111111111110010111100010;
    rom[11078] = 25'b1111111111110010111000101;
    rom[11079] = 25'b1111111111110010110100111;
    rom[11080] = 25'b1111111111110010110001010;
    rom[11081] = 25'b1111111111110010101101100;
    rom[11082] = 25'b1111111111110010101001111;
    rom[11083] = 25'b1111111111110010100110001;
    rom[11084] = 25'b1111111111110010100010100;
    rom[11085] = 25'b1111111111110010011110110;
    rom[11086] = 25'b1111111111110010011011001;
    rom[11087] = 25'b1111111111110010010111011;
    rom[11088] = 25'b1111111111110010010011101;
    rom[11089] = 25'b1111111111110010010000000;
    rom[11090] = 25'b1111111111110010001100010;
    rom[11091] = 25'b1111111111110010001000101;
    rom[11092] = 25'b1111111111110010000100111;
    rom[11093] = 25'b1111111111110010000001010;
    rom[11094] = 25'b1111111111110001111101100;
    rom[11095] = 25'b1111111111110001111001111;
    rom[11096] = 25'b1111111111110001110110001;
    rom[11097] = 25'b1111111111110001110010100;
    rom[11098] = 25'b1111111111110001101110110;
    rom[11099] = 25'b1111111111110001101011001;
    rom[11100] = 25'b1111111111110001100111011;
    rom[11101] = 25'b1111111111110001100011101;
    rom[11102] = 25'b1111111111110001100000000;
    rom[11103] = 25'b1111111111110001011100010;
    rom[11104] = 25'b1111111111110001011000101;
    rom[11105] = 25'b1111111111110001010100111;
    rom[11106] = 25'b1111111111110001010001001;
    rom[11107] = 25'b1111111111110001001101100;
    rom[11108] = 25'b1111111111110001001001110;
    rom[11109] = 25'b1111111111110001000110000;
    rom[11110] = 25'b1111111111110001000010010;
    rom[11111] = 25'b1111111111110000111110101;
    rom[11112] = 25'b1111111111110000111010111;
    rom[11113] = 25'b1111111111110000110111001;
    rom[11114] = 25'b1111111111110000110011011;
    rom[11115] = 25'b1111111111110000101111101;
    rom[11116] = 25'b1111111111110000101100000;
    rom[11117] = 25'b1111111111110000101000010;
    rom[11118] = 25'b1111111111110000100100100;
    rom[11119] = 25'b1111111111110000100000111;
    rom[11120] = 25'b1111111111110000011101001;
    rom[11121] = 25'b1111111111110000011001011;
    rom[11122] = 25'b1111111111110000010101101;
    rom[11123] = 25'b1111111111110000010010000;
    rom[11124] = 25'b1111111111110000001110010;
    rom[11125] = 25'b1111111111110000001010100;
    rom[11126] = 25'b1111111111110000000110110;
    rom[11127] = 25'b1111111111110000000011000;
    rom[11128] = 25'b1111111111101111111111010;
    rom[11129] = 25'b1111111111101111111011100;
    rom[11130] = 25'b1111111111101111110111111;
    rom[11131] = 25'b1111111111101111110100001;
    rom[11132] = 25'b1111111111101111110000011;
    rom[11133] = 25'b1111111111101111101100101;
    rom[11134] = 25'b1111111111101111101000111;
    rom[11135] = 25'b1111111111101111100101001;
    rom[11136] = 25'b1111111111101111100001011;
    rom[11137] = 25'b1111111111101111011101101;
    rom[11138] = 25'b1111111111101111011010000;
    rom[11139] = 25'b1111111111101111010110010;
    rom[11140] = 25'b1111111111101111010010100;
    rom[11141] = 25'b1111111111101111001110110;
    rom[11142] = 25'b1111111111101111001011000;
    rom[11143] = 25'b1111111111101111000111010;
    rom[11144] = 25'b1111111111101111000011011;
    rom[11145] = 25'b1111111111101110111111110;
    rom[11146] = 25'b1111111111101110111100000;
    rom[11147] = 25'b1111111111101110111000010;
    rom[11148] = 25'b1111111111101110110100100;
    rom[11149] = 25'b1111111111101110110000110;
    rom[11150] = 25'b1111111111101110101101000;
    rom[11151] = 25'b1111111111101110101001010;
    rom[11152] = 25'b1111111111101110100101100;
    rom[11153] = 25'b1111111111101110100001110;
    rom[11154] = 25'b1111111111101110011110000;
    rom[11155] = 25'b1111111111101110011010010;
    rom[11156] = 25'b1111111111101110010110100;
    rom[11157] = 25'b1111111111101110010010101;
    rom[11158] = 25'b1111111111101110001111000;
    rom[11159] = 25'b1111111111101110001011010;
    rom[11160] = 25'b1111111111101110000111100;
    rom[11161] = 25'b1111111111101110000011101;
    rom[11162] = 25'b1111111111101101111111111;
    rom[11163] = 25'b1111111111101101111100001;
    rom[11164] = 25'b1111111111101101111000100;
    rom[11165] = 25'b1111111111101101110100101;
    rom[11166] = 25'b1111111111101101110000111;
    rom[11167] = 25'b1111111111101101101101001;
    rom[11168] = 25'b1111111111101101101001011;
    rom[11169] = 25'b1111111111101101100101101;
    rom[11170] = 25'b1111111111101101100001111;
    rom[11171] = 25'b1111111111101101011110000;
    rom[11172] = 25'b1111111111101101011010010;
    rom[11173] = 25'b1111111111101101010110100;
    rom[11174] = 25'b1111111111101101010010110;
    rom[11175] = 25'b1111111111101101001111000;
    rom[11176] = 25'b1111111111101101001011010;
    rom[11177] = 25'b1111111111101101000111011;
    rom[11178] = 25'b1111111111101101000011101;
    rom[11179] = 25'b1111111111101100111111111;
    rom[11180] = 25'b1111111111101100111100001;
    rom[11181] = 25'b1111111111101100111000011;
    rom[11182] = 25'b1111111111101100110100100;
    rom[11183] = 25'b1111111111101100110000111;
    rom[11184] = 25'b1111111111101100101101000;
    rom[11185] = 25'b1111111111101100101001010;
    rom[11186] = 25'b1111111111101100100101011;
    rom[11187] = 25'b1111111111101100100001110;
    rom[11188] = 25'b1111111111101100011101111;
    rom[11189] = 25'b1111111111101100011010001;
    rom[11190] = 25'b1111111111101100010110011;
    rom[11191] = 25'b1111111111101100010010100;
    rom[11192] = 25'b1111111111101100001110111;
    rom[11193] = 25'b1111111111101100001011000;
    rom[11194] = 25'b1111111111101100000111010;
    rom[11195] = 25'b1111111111101100000011011;
    rom[11196] = 25'b1111111111101011111111110;
    rom[11197] = 25'b1111111111101011111011111;
    rom[11198] = 25'b1111111111101011111000000;
    rom[11199] = 25'b1111111111101011110100010;
    rom[11200] = 25'b1111111111101011110000100;
    rom[11201] = 25'b1111111111101011101100110;
    rom[11202] = 25'b1111111111101011101000111;
    rom[11203] = 25'b1111111111101011100101001;
    rom[11204] = 25'b1111111111101011100001011;
    rom[11205] = 25'b1111111111101011011101101;
    rom[11206] = 25'b1111111111101011011001110;
    rom[11207] = 25'b1111111111101011010110000;
    rom[11208] = 25'b1111111111101011010010010;
    rom[11209] = 25'b1111111111101011001110011;
    rom[11210] = 25'b1111111111101011001010101;
    rom[11211] = 25'b1111111111101011000110111;
    rom[11212] = 25'b1111111111101011000011000;
    rom[11213] = 25'b1111111111101010111111010;
    rom[11214] = 25'b1111111111101010111011011;
    rom[11215] = 25'b1111111111101010110111101;
    rom[11216] = 25'b1111111111101010110011111;
    rom[11217] = 25'b1111111111101010110000000;
    rom[11218] = 25'b1111111111101010101100010;
    rom[11219] = 25'b1111111111101010101000100;
    rom[11220] = 25'b1111111111101010100100101;
    rom[11221] = 25'b1111111111101010100000111;
    rom[11222] = 25'b1111111111101010011101001;
    rom[11223] = 25'b1111111111101010011001010;
    rom[11224] = 25'b1111111111101010010101011;
    rom[11225] = 25'b1111111111101010010001101;
    rom[11226] = 25'b1111111111101010001101111;
    rom[11227] = 25'b1111111111101010001010000;
    rom[11228] = 25'b1111111111101010000110010;
    rom[11229] = 25'b1111111111101010000010100;
    rom[11230] = 25'b1111111111101001111110101;
    rom[11231] = 25'b1111111111101001111010111;
    rom[11232] = 25'b1111111111101001110111001;
    rom[11233] = 25'b1111111111101001110011010;
    rom[11234] = 25'b1111111111101001101111011;
    rom[11235] = 25'b1111111111101001101011101;
    rom[11236] = 25'b1111111111101001100111111;
    rom[11237] = 25'b1111111111101001100100000;
    rom[11238] = 25'b1111111111101001100000010;
    rom[11239] = 25'b1111111111101001011100100;
    rom[11240] = 25'b1111111111101001011000101;
    rom[11241] = 25'b1111111111101001010100110;
    rom[11242] = 25'b1111111111101001010001000;
    rom[11243] = 25'b1111111111101001001101010;
    rom[11244] = 25'b1111111111101001001001011;
    rom[11245] = 25'b1111111111101001000101101;
    rom[11246] = 25'b1111111111101001000001110;
    rom[11247] = 25'b1111111111101000111110000;
    rom[11248] = 25'b1111111111101000111010001;
    rom[11249] = 25'b1111111111101000110110011;
    rom[11250] = 25'b1111111111101000110010100;
    rom[11251] = 25'b1111111111101000101110110;
    rom[11252] = 25'b1111111111101000101011000;
    rom[11253] = 25'b1111111111101000100111001;
    rom[11254] = 25'b1111111111101000100011010;
    rom[11255] = 25'b1111111111101000011111100;
    rom[11256] = 25'b1111111111101000011011101;
    rom[11257] = 25'b1111111111101000010111111;
    rom[11258] = 25'b1111111111101000010100001;
    rom[11259] = 25'b1111111111101000010000010;
    rom[11260] = 25'b1111111111101000001100011;
    rom[11261] = 25'b1111111111101000001000101;
    rom[11262] = 25'b1111111111101000000100110;
    rom[11263] = 25'b1111111111101000000000111;
    rom[11264] = 25'b1111111111100111111101010;
    rom[11265] = 25'b1111111111100111111001011;
    rom[11266] = 25'b1111111111100111110101100;
    rom[11267] = 25'b1111111111100111110001110;
    rom[11268] = 25'b1111111111100111101101111;
    rom[11269] = 25'b1111111111100111101010000;
    rom[11270] = 25'b1111111111100111100110011;
    rom[11271] = 25'b1111111111100111100010100;
    rom[11272] = 25'b1111111111100111011110101;
    rom[11273] = 25'b1111111111100111011010111;
    rom[11274] = 25'b1111111111100111010111000;
    rom[11275] = 25'b1111111111100111010011001;
    rom[11276] = 25'b1111111111100111001111011;
    rom[11277] = 25'b1111111111100111001011100;
    rom[11278] = 25'b1111111111100111000111110;
    rom[11279] = 25'b1111111111100111000100000;
    rom[11280] = 25'b1111111111100111000000001;
    rom[11281] = 25'b1111111111100110111100010;
    rom[11282] = 25'b1111111111100110111000100;
    rom[11283] = 25'b1111111111100110110100101;
    rom[11284] = 25'b1111111111100110110000110;
    rom[11285] = 25'b1111111111100110101101000;
    rom[11286] = 25'b1111111111100110101001010;
    rom[11287] = 25'b1111111111100110100101011;
    rom[11288] = 25'b1111111111100110100001101;
    rom[11289] = 25'b1111111111100110011101110;
    rom[11290] = 25'b1111111111100110011001111;
    rom[11291] = 25'b1111111111100110010110001;
    rom[11292] = 25'b1111111111100110010010010;
    rom[11293] = 25'b1111111111100110001110100;
    rom[11294] = 25'b1111111111100110001010101;
    rom[11295] = 25'b1111111111100110000110110;
    rom[11296] = 25'b1111111111100110000011000;
    rom[11297] = 25'b1111111111100101111111010;
    rom[11298] = 25'b1111111111100101111011011;
    rom[11299] = 25'b1111111111100101110111101;
    rom[11300] = 25'b1111111111100101110011110;
    rom[11301] = 25'b1111111111100101101111111;
    rom[11302] = 25'b1111111111100101101100001;
    rom[11303] = 25'b1111111111100101101000010;
    rom[11304] = 25'b1111111111100101100100011;
    rom[11305] = 25'b1111111111100101100000101;
    rom[11306] = 25'b1111111111100101011100110;
    rom[11307] = 25'b1111111111100101011001000;
    rom[11308] = 25'b1111111111100101010101010;
    rom[11309] = 25'b1111111111100101010001011;
    rom[11310] = 25'b1111111111100101001101100;
    rom[11311] = 25'b1111111111100101001001110;
    rom[11312] = 25'b1111111111100101000101111;
    rom[11313] = 25'b1111111111100101000010000;
    rom[11314] = 25'b1111111111100100111110010;
    rom[11315] = 25'b1111111111100100111010011;
    rom[11316] = 25'b1111111111100100110110101;
    rom[11317] = 25'b1111111111100100110010110;
    rom[11318] = 25'b1111111111100100101111000;
    rom[11319] = 25'b1111111111100100101011001;
    rom[11320] = 25'b1111111111100100100111011;
    rom[11321] = 25'b1111111111100100100011100;
    rom[11322] = 25'b1111111111100100011111101;
    rom[11323] = 25'b1111111111100100011011111;
    rom[11324] = 25'b1111111111100100011000000;
    rom[11325] = 25'b1111111111100100010100010;
    rom[11326] = 25'b1111111111100100010000011;
    rom[11327] = 25'b1111111111100100001100100;
    rom[11328] = 25'b1111111111100100001000110;
    rom[11329] = 25'b1111111111100100000101000;
    rom[11330] = 25'b1111111111100100000001001;
    rom[11331] = 25'b1111111111100011111101011;
    rom[11332] = 25'b1111111111100011111001100;
    rom[11333] = 25'b1111111111100011110101101;
    rom[11334] = 25'b1111111111100011110001111;
    rom[11335] = 25'b1111111111100011101110000;
    rom[11336] = 25'b1111111111100011101010001;
    rom[11337] = 25'b1111111111100011100110011;
    rom[11338] = 25'b1111111111100011100010101;
    rom[11339] = 25'b1111111111100011011110110;
    rom[11340] = 25'b1111111111100011011011000;
    rom[11341] = 25'b1111111111100011010111001;
    rom[11342] = 25'b1111111111100011010011010;
    rom[11343] = 25'b1111111111100011001111100;
    rom[11344] = 25'b1111111111100011001011101;
    rom[11345] = 25'b1111111111100011000111110;
    rom[11346] = 25'b1111111111100011000100000;
    rom[11347] = 25'b1111111111100011000000010;
    rom[11348] = 25'b1111111111100010111100011;
    rom[11349] = 25'b1111111111100010111000101;
    rom[11350] = 25'b1111111111100010110100110;
    rom[11351] = 25'b1111111111100010110000111;
    rom[11352] = 25'b1111111111100010101101001;
    rom[11353] = 25'b1111111111100010101001010;
    rom[11354] = 25'b1111111111100010100101100;
    rom[11355] = 25'b1111111111100010100001110;
    rom[11356] = 25'b1111111111100010011101111;
    rom[11357] = 25'b1111111111100010011010000;
    rom[11358] = 25'b1111111111100010010110010;
    rom[11359] = 25'b1111111111100010010010011;
    rom[11360] = 25'b1111111111100010001110100;
    rom[11361] = 25'b1111111111100010001010111;
    rom[11362] = 25'b1111111111100010000111000;
    rom[11363] = 25'b1111111111100010000011001;
    rom[11364] = 25'b1111111111100001111111011;
    rom[11365] = 25'b1111111111100001111011100;
    rom[11366] = 25'b1111111111100001110111101;
    rom[11367] = 25'b1111111111100001110100000;
    rom[11368] = 25'b1111111111100001110000001;
    rom[11369] = 25'b1111111111100001101100010;
    rom[11370] = 25'b1111111111100001101000100;
    rom[11371] = 25'b1111111111100001100100101;
    rom[11372] = 25'b1111111111100001100000111;
    rom[11373] = 25'b1111111111100001011101001;
    rom[11374] = 25'b1111111111100001011001010;
    rom[11375] = 25'b1111111111100001010101011;
    rom[11376] = 25'b1111111111100001010001101;
    rom[11377] = 25'b1111111111100001001101111;
    rom[11378] = 25'b1111111111100001001010000;
    rom[11379] = 25'b1111111111100001000110001;
    rom[11380] = 25'b1111111111100001000010011;
    rom[11381] = 25'b1111111111100000111110100;
    rom[11382] = 25'b1111111111100000111010110;
    rom[11383] = 25'b1111111111100000110111000;
    rom[11384] = 25'b1111111111100000110011001;
    rom[11385] = 25'b1111111111100000101111010;
    rom[11386] = 25'b1111111111100000101011101;
    rom[11387] = 25'b1111111111100000100111110;
    rom[11388] = 25'b1111111111100000100011111;
    rom[11389] = 25'b1111111111100000100000001;
    rom[11390] = 25'b1111111111100000011100011;
    rom[11391] = 25'b1111111111100000011000100;
    rom[11392] = 25'b1111111111100000010100110;
    rom[11393] = 25'b1111111111100000010001000;
    rom[11394] = 25'b1111111111100000001101001;
    rom[11395] = 25'b1111111111100000001001010;
    rom[11396] = 25'b1111111111100000000101100;
    rom[11397] = 25'b1111111111100000000001110;
    rom[11398] = 25'b1111111111011111111101111;
    rom[11399] = 25'b1111111111011111111010001;
    rom[11400] = 25'b1111111111011111110110011;
    rom[11401] = 25'b1111111111011111110010100;
    rom[11402] = 25'b1111111111011111101110101;
    rom[11403] = 25'b1111111111011111101011000;
    rom[11404] = 25'b1111111111011111100111001;
    rom[11405] = 25'b1111111111011111100011010;
    rom[11406] = 25'b1111111111011111011111100;
    rom[11407] = 25'b1111111111011111011011110;
    rom[11408] = 25'b1111111111011111010111111;
    rom[11409] = 25'b1111111111011111010100001;
    rom[11410] = 25'b1111111111011111010000011;
    rom[11411] = 25'b1111111111011111001100101;
    rom[11412] = 25'b1111111111011111001000110;
    rom[11413] = 25'b1111111111011111000101000;
    rom[11414] = 25'b1111111111011111000001010;
    rom[11415] = 25'b1111111111011110111101011;
    rom[11416] = 25'b1111111111011110111001101;
    rom[11417] = 25'b1111111111011110110101110;
    rom[11418] = 25'b1111111111011110110010000;
    rom[11419] = 25'b1111111111011110101110010;
    rom[11420] = 25'b1111111111011110101010011;
    rom[11421] = 25'b1111111111011110100110101;
    rom[11422] = 25'b1111111111011110100010111;
    rom[11423] = 25'b1111111111011110011111001;
    rom[11424] = 25'b1111111111011110011011010;
    rom[11425] = 25'b1111111111011110010111100;
    rom[11426] = 25'b1111111111011110010011110;
    rom[11427] = 25'b1111111111011110010000000;
    rom[11428] = 25'b1111111111011110001100001;
    rom[11429] = 25'b1111111111011110001000011;
    rom[11430] = 25'b1111111111011110000100101;
    rom[11431] = 25'b1111111111011110000000111;
    rom[11432] = 25'b1111111111011101111101000;
    rom[11433] = 25'b1111111111011101111001010;
    rom[11434] = 25'b1111111111011101110101100;
    rom[11435] = 25'b1111111111011101110001110;
    rom[11436] = 25'b1111111111011101101101111;
    rom[11437] = 25'b1111111111011101101010001;
    rom[11438] = 25'b1111111111011101100110011;
    rom[11439] = 25'b1111111111011101100010101;
    rom[11440] = 25'b1111111111011101011110111;
    rom[11441] = 25'b1111111111011101011011000;
    rom[11442] = 25'b1111111111011101010111010;
    rom[11443] = 25'b1111111111011101010011100;
    rom[11444] = 25'b1111111111011101001111110;
    rom[11445] = 25'b1111111111011101001100000;
    rom[11446] = 25'b1111111111011101001000001;
    rom[11447] = 25'b1111111111011101000100100;
    rom[11448] = 25'b1111111111011101000000110;
    rom[11449] = 25'b1111111111011100111100111;
    rom[11450] = 25'b1111111111011100111001001;
    rom[11451] = 25'b1111111111011100110101011;
    rom[11452] = 25'b1111111111011100110001101;
    rom[11453] = 25'b1111111111011100101101111;
    rom[11454] = 25'b1111111111011100101010001;
    rom[11455] = 25'b1111111111011100100110010;
    rom[11456] = 25'b1111111111011100100010100;
    rom[11457] = 25'b1111111111011100011110110;
    rom[11458] = 25'b1111111111011100011011000;
    rom[11459] = 25'b1111111111011100010111010;
    rom[11460] = 25'b1111111111011100010011100;
    rom[11461] = 25'b1111111111011100001111110;
    rom[11462] = 25'b1111111111011100001100000;
    rom[11463] = 25'b1111111111011100001000010;
    rom[11464] = 25'b1111111111011100000100100;
    rom[11465] = 25'b1111111111011100000000110;
    rom[11466] = 25'b1111111111011011111101000;
    rom[11467] = 25'b1111111111011011111001001;
    rom[11468] = 25'b1111111111011011110101011;
    rom[11469] = 25'b1111111111011011110001110;
    rom[11470] = 25'b1111111111011011101110000;
    rom[11471] = 25'b1111111111011011101010010;
    rom[11472] = 25'b1111111111011011100110100;
    rom[11473] = 25'b1111111111011011100010110;
    rom[11474] = 25'b1111111111011011011110111;
    rom[11475] = 25'b1111111111011011011011010;
    rom[11476] = 25'b1111111111011011010111100;
    rom[11477] = 25'b1111111111011011010011110;
    rom[11478] = 25'b1111111111011011010000000;
    rom[11479] = 25'b1111111111011011001100010;
    rom[11480] = 25'b1111111111011011001000100;
    rom[11481] = 25'b1111111111011011000100110;
    rom[11482] = 25'b1111111111011011000001000;
    rom[11483] = 25'b1111111111011010111101010;
    rom[11484] = 25'b1111111111011010111001101;
    rom[11485] = 25'b1111111111011010110101111;
    rom[11486] = 25'b1111111111011010110010001;
    rom[11487] = 25'b1111111111011010101110011;
    rom[11488] = 25'b1111111111011010101010101;
    rom[11489] = 25'b1111111111011010100110111;
    rom[11490] = 25'b1111111111011010100011001;
    rom[11491] = 25'b1111111111011010011111011;
    rom[11492] = 25'b1111111111011010011011110;
    rom[11493] = 25'b1111111111011010011000000;
    rom[11494] = 25'b1111111111011010010100010;
    rom[11495] = 25'b1111111111011010010000100;
    rom[11496] = 25'b1111111111011010001100111;
    rom[11497] = 25'b1111111111011010001001001;
    rom[11498] = 25'b1111111111011010000101011;
    rom[11499] = 25'b1111111111011010000001101;
    rom[11500] = 25'b1111111111011001111101111;
    rom[11501] = 25'b1111111111011001111010001;
    rom[11502] = 25'b1111111111011001110110100;
    rom[11503] = 25'b1111111111011001110010110;
    rom[11504] = 25'b1111111111011001101111000;
    rom[11505] = 25'b1111111111011001101011011;
    rom[11506] = 25'b1111111111011001100111101;
    rom[11507] = 25'b1111111111011001100011111;
    rom[11508] = 25'b1111111111011001100000010;
    rom[11509] = 25'b1111111111011001011100100;
    rom[11510] = 25'b1111111111011001011000111;
    rom[11511] = 25'b1111111111011001010101001;
    rom[11512] = 25'b1111111111011001010001011;
    rom[11513] = 25'b1111111111011001001101101;
    rom[11514] = 25'b1111111111011001001010000;
    rom[11515] = 25'b1111111111011001000110010;
    rom[11516] = 25'b1111111111011001000010100;
    rom[11517] = 25'b1111111111011000111110111;
    rom[11518] = 25'b1111111111011000111011001;
    rom[11519] = 25'b1111111111011000110111100;
    rom[11520] = 25'b1111111111011000110011110;
    rom[11521] = 25'b1111111111011000110000000;
    rom[11522] = 25'b1111111111011000101100011;
    rom[11523] = 25'b1111111111011000101000101;
    rom[11524] = 25'b1111111111011000100101000;
    rom[11525] = 25'b1111111111011000100001010;
    rom[11526] = 25'b1111111111011000011101101;
    rom[11527] = 25'b1111111111011000011001111;
    rom[11528] = 25'b1111111111011000010110010;
    rom[11529] = 25'b1111111111011000010010100;
    rom[11530] = 25'b1111111111011000001110111;
    rom[11531] = 25'b1111111111011000001011001;
    rom[11532] = 25'b1111111111011000000111100;
    rom[11533] = 25'b1111111111011000000011111;
    rom[11534] = 25'b1111111111011000000000001;
    rom[11535] = 25'b1111111111010111111100100;
    rom[11536] = 25'b1111111111010111111000110;
    rom[11537] = 25'b1111111111010111110101001;
    rom[11538] = 25'b1111111111010111110001100;
    rom[11539] = 25'b1111111111010111101101110;
    rom[11540] = 25'b1111111111010111101010001;
    rom[11541] = 25'b1111111111010111100110011;
    rom[11542] = 25'b1111111111010111100010110;
    rom[11543] = 25'b1111111111010111011111000;
    rom[11544] = 25'b1111111111010111011011011;
    rom[11545] = 25'b1111111111010111010111110;
    rom[11546] = 25'b1111111111010111010100001;
    rom[11547] = 25'b1111111111010111010000011;
    rom[11548] = 25'b1111111111010111001100110;
    rom[11549] = 25'b1111111111010111001001001;
    rom[11550] = 25'b1111111111010111000101100;
    rom[11551] = 25'b1111111111010111000001111;
    rom[11552] = 25'b1111111111010110111110001;
    rom[11553] = 25'b1111111111010110111010100;
    rom[11554] = 25'b1111111111010110110110110;
    rom[11555] = 25'b1111111111010110110011001;
    rom[11556] = 25'b1111111111010110101111100;
    rom[11557] = 25'b1111111111010110101011111;
    rom[11558] = 25'b1111111111010110101000010;
    rom[11559] = 25'b1111111111010110100100101;
    rom[11560] = 25'b1111111111010110100001000;
    rom[11561] = 25'b1111111111010110011101010;
    rom[11562] = 25'b1111111111010110011001101;
    rom[11563] = 25'b1111111111010110010110000;
    rom[11564] = 25'b1111111111010110010010011;
    rom[11565] = 25'b1111111111010110001110110;
    rom[11566] = 25'b1111111111010110001011001;
    rom[11567] = 25'b1111111111010110000111100;
    rom[11568] = 25'b1111111111010110000011110;
    rom[11569] = 25'b1111111111010110000000010;
    rom[11570] = 25'b1111111111010101111100101;
    rom[11571] = 25'b1111111111010101111001000;
    rom[11572] = 25'b1111111111010101110101011;
    rom[11573] = 25'b1111111111010101110001110;
    rom[11574] = 25'b1111111111010101101110000;
    rom[11575] = 25'b1111111111010101101010100;
    rom[11576] = 25'b1111111111010101100110111;
    rom[11577] = 25'b1111111111010101100011010;
    rom[11578] = 25'b1111111111010101011111101;
    rom[11579] = 25'b1111111111010101011100000;
    rom[11580] = 25'b1111111111010101011000011;
    rom[11581] = 25'b1111111111010101010100110;
    rom[11582] = 25'b1111111111010101010001010;
    rom[11583] = 25'b1111111111010101001101100;
    rom[11584] = 25'b1111111111010101001001111;
    rom[11585] = 25'b1111111111010101000110011;
    rom[11586] = 25'b1111111111010101000010110;
    rom[11587] = 25'b1111111111010100111111001;
    rom[11588] = 25'b1111111111010100111011100;
    rom[11589] = 25'b1111111111010100111000000;
    rom[11590] = 25'b1111111111010100110100011;
    rom[11591] = 25'b1111111111010100110000110;
    rom[11592] = 25'b1111111111010100101101001;
    rom[11593] = 25'b1111111111010100101001101;
    rom[11594] = 25'b1111111111010100100110000;
    rom[11595] = 25'b1111111111010100100010011;
    rom[11596] = 25'b1111111111010100011110110;
    rom[11597] = 25'b1111111111010100011011010;
    rom[11598] = 25'b1111111111010100010111101;
    rom[11599] = 25'b1111111111010100010100000;
    rom[11600] = 25'b1111111111010100010000100;
    rom[11601] = 25'b1111111111010100001100111;
    rom[11602] = 25'b1111111111010100001001010;
    rom[11603] = 25'b1111111111010100000101110;
    rom[11604] = 25'b1111111111010100000010001;
    rom[11605] = 25'b1111111111010011111110100;
    rom[11606] = 25'b1111111111010011111011000;
    rom[11607] = 25'b1111111111010011110111100;
    rom[11608] = 25'b1111111111010011110011111;
    rom[11609] = 25'b1111111111010011110000011;
    rom[11610] = 25'b1111111111010011101100110;
    rom[11611] = 25'b1111111111010011101001001;
    rom[11612] = 25'b1111111111010011100101101;
    rom[11613] = 25'b1111111111010011100010000;
    rom[11614] = 25'b1111111111010011011110100;
    rom[11615] = 25'b1111111111010011011011000;
    rom[11616] = 25'b1111111111010011010111011;
    rom[11617] = 25'b1111111111010011010011111;
    rom[11618] = 25'b1111111111010011010000011;
    rom[11619] = 25'b1111111111010011001100110;
    rom[11620] = 25'b1111111111010011001001010;
    rom[11621] = 25'b1111111111010011000101101;
    rom[11622] = 25'b1111111111010011000010001;
    rom[11623] = 25'b1111111111010010111110101;
    rom[11624] = 25'b1111111111010010111011000;
    rom[11625] = 25'b1111111111010010110111101;
    rom[11626] = 25'b1111111111010010110100000;
    rom[11627] = 25'b1111111111010010110000100;
    rom[11628] = 25'b1111111111010010101100111;
    rom[11629] = 25'b1111111111010010101001011;
    rom[11630] = 25'b1111111111010010100101111;
    rom[11631] = 25'b1111111111010010100010011;
    rom[11632] = 25'b1111111111010010011110111;
    rom[11633] = 25'b1111111111010010011011010;
    rom[11634] = 25'b1111111111010010010111111;
    rom[11635] = 25'b1111111111010010010100010;
    rom[11636] = 25'b1111111111010010010000110;
    rom[11637] = 25'b1111111111010010001101010;
    rom[11638] = 25'b1111111111010010001001110;
    rom[11639] = 25'b1111111111010010000110010;
    rom[11640] = 25'b1111111111010010000010110;
    rom[11641] = 25'b1111111111010001111111010;
    rom[11642] = 25'b1111111111010001111011110;
    rom[11643] = 25'b1111111111010001111000010;
    rom[11644] = 25'b1111111111010001110100110;
    rom[11645] = 25'b1111111111010001110001010;
    rom[11646] = 25'b1111111111010001101101110;
    rom[11647] = 25'b1111111111010001101010010;
    rom[11648] = 25'b1111111111010001100110110;
    rom[11649] = 25'b1111111111010001100011010;
    rom[11650] = 25'b1111111111010001011111110;
    rom[11651] = 25'b1111111111010001011100010;
    rom[11652] = 25'b1111111111010001011000110;
    rom[11653] = 25'b1111111111010001010101011;
    rom[11654] = 25'b1111111111010001010001111;
    rom[11655] = 25'b1111111111010001001110011;
    rom[11656] = 25'b1111111111010001001010111;
    rom[11657] = 25'b1111111111010001000111011;
    rom[11658] = 25'b1111111111010001000100000;
    rom[11659] = 25'b1111111111010001000000100;
    rom[11660] = 25'b1111111111010000111101000;
    rom[11661] = 25'b1111111111010000111001100;
    rom[11662] = 25'b1111111111010000110110000;
    rom[11663] = 25'b1111111111010000110010101;
    rom[11664] = 25'b1111111111010000101111001;
    rom[11665] = 25'b1111111111010000101011101;
    rom[11666] = 25'b1111111111010000101000010;
    rom[11667] = 25'b1111111111010000100100110;
    rom[11668] = 25'b1111111111010000100001010;
    rom[11669] = 25'b1111111111010000011101111;
    rom[11670] = 25'b1111111111010000011010100;
    rom[11671] = 25'b1111111111010000010111000;
    rom[11672] = 25'b1111111111010000010011101;
    rom[11673] = 25'b1111111111010000010000001;
    rom[11674] = 25'b1111111111010000001100101;
    rom[11675] = 25'b1111111111010000001001010;
    rom[11676] = 25'b1111111111010000000101111;
    rom[11677] = 25'b1111111111010000000010011;
    rom[11678] = 25'b1111111111001111111111000;
    rom[11679] = 25'b1111111111001111111011101;
    rom[11680] = 25'b1111111111001111111000001;
    rom[11681] = 25'b1111111111001111110100101;
    rom[11682] = 25'b1111111111001111110001010;
    rom[11683] = 25'b1111111111001111101101111;
    rom[11684] = 25'b1111111111001111101010100;
    rom[11685] = 25'b1111111111001111100111000;
    rom[11686] = 25'b1111111111001111100011101;
    rom[11687] = 25'b1111111111001111100000010;
    rom[11688] = 25'b1111111111001111011100110;
    rom[11689] = 25'b1111111111001111011001011;
    rom[11690] = 25'b1111111111001111010110000;
    rom[11691] = 25'b1111111111001111010010101;
    rom[11692] = 25'b1111111111001111001111010;
    rom[11693] = 25'b1111111111001111001011111;
    rom[11694] = 25'b1111111111001111001000011;
    rom[11695] = 25'b1111111111001111000101000;
    rom[11696] = 25'b1111111111001111000001101;
    rom[11697] = 25'b1111111111001110111110010;
    rom[11698] = 25'b1111111111001110111010111;
    rom[11699] = 25'b1111111111001110110111100;
    rom[11700] = 25'b1111111111001110110100001;
    rom[11701] = 25'b1111111111001110110000110;
    rom[11702] = 25'b1111111111001110101101011;
    rom[11703] = 25'b1111111111001110101010000;
    rom[11704] = 25'b1111111111001110100110101;
    rom[11705] = 25'b1111111111001110100011010;
    rom[11706] = 25'b1111111111001110011111111;
    rom[11707] = 25'b1111111111001110011100100;
    rom[11708] = 25'b1111111111001110011001001;
    rom[11709] = 25'b1111111111001110010101110;
    rom[11710] = 25'b1111111111001110010010011;
    rom[11711] = 25'b1111111111001110001111001;
    rom[11712] = 25'b1111111111001110001011110;
    rom[11713] = 25'b1111111111001110001000011;
    rom[11714] = 25'b1111111111001110000101001;
    rom[11715] = 25'b1111111111001110000001110;
    rom[11716] = 25'b1111111111001101111110011;
    rom[11717] = 25'b1111111111001101111011001;
    rom[11718] = 25'b1111111111001101110111110;
    rom[11719] = 25'b1111111111001101110100011;
    rom[11720] = 25'b1111111111001101110001001;
    rom[11721] = 25'b1111111111001101101101110;
    rom[11722] = 25'b1111111111001101101010011;
    rom[11723] = 25'b1111111111001101100111001;
    rom[11724] = 25'b1111111111001101100011110;
    rom[11725] = 25'b1111111111001101100000100;
    rom[11726] = 25'b1111111111001101011101001;
    rom[11727] = 25'b1111111111001101011001111;
    rom[11728] = 25'b1111111111001101010110100;
    rom[11729] = 25'b1111111111001101010011010;
    rom[11730] = 25'b1111111111001101001111111;
    rom[11731] = 25'b1111111111001101001100101;
    rom[11732] = 25'b1111111111001101001001010;
    rom[11733] = 25'b1111111111001101000110000;
    rom[11734] = 25'b1111111111001101000010101;
    rom[11735] = 25'b1111111111001100111111011;
    rom[11736] = 25'b1111111111001100111100001;
    rom[11737] = 25'b1111111111001100111000111;
    rom[11738] = 25'b1111111111001100110101100;
    rom[11739] = 25'b1111111111001100110010010;
    rom[11740] = 25'b1111111111001100101111000;
    rom[11741] = 25'b1111111111001100101011110;
    rom[11742] = 25'b1111111111001100101000011;
    rom[11743] = 25'b1111111111001100100101001;
    rom[11744] = 25'b1111111111001100100001111;
    rom[11745] = 25'b1111111111001100011110101;
    rom[11746] = 25'b1111111111001100011011011;
    rom[11747] = 25'b1111111111001100011000001;
    rom[11748] = 25'b1111111111001100010100111;
    rom[11749] = 25'b1111111111001100010001100;
    rom[11750] = 25'b1111111111001100001110010;
    rom[11751] = 25'b1111111111001100001011001;
    rom[11752] = 25'b1111111111001100000111111;
    rom[11753] = 25'b1111111111001100000100101;
    rom[11754] = 25'b1111111111001100000001010;
    rom[11755] = 25'b1111111111001011111110001;
    rom[11756] = 25'b1111111111001011111010111;
    rom[11757] = 25'b1111111111001011110111101;
    rom[11758] = 25'b1111111111001011110100011;
    rom[11759] = 25'b1111111111001011110001001;
    rom[11760] = 25'b1111111111001011101110000;
    rom[11761] = 25'b1111111111001011101010110;
    rom[11762] = 25'b1111111111001011100111100;
    rom[11763] = 25'b1111111111001011100100010;
    rom[11764] = 25'b1111111111001011100001001;
    rom[11765] = 25'b1111111111001011011101111;
    rom[11766] = 25'b1111111111001011011010101;
    rom[11767] = 25'b1111111111001011010111100;
    rom[11768] = 25'b1111111111001011010100010;
    rom[11769] = 25'b1111111111001011010001000;
    rom[11770] = 25'b1111111111001011001101111;
    rom[11771] = 25'b1111111111001011001010101;
    rom[11772] = 25'b1111111111001011000111011;
    rom[11773] = 25'b1111111111001011000100010;
    rom[11774] = 25'b1111111111001011000001000;
    rom[11775] = 25'b1111111111001010111101111;
    rom[11776] = 25'b1111111111001010111010110;
    rom[11777] = 25'b1111111111001010110111100;
    rom[11778] = 25'b1111111111001010110100011;
    rom[11779] = 25'b1111111111001010110001001;
    rom[11780] = 25'b1111111111001010101110000;
    rom[11781] = 25'b1111111111001010101010111;
    rom[11782] = 25'b1111111111001010100111101;
    rom[11783] = 25'b1111111111001010100100100;
    rom[11784] = 25'b1111111111001010100001010;
    rom[11785] = 25'b1111111111001010011110010;
    rom[11786] = 25'b1111111111001010011011000;
    rom[11787] = 25'b1111111111001010010111111;
    rom[11788] = 25'b1111111111001010010100110;
    rom[11789] = 25'b1111111111001010010001101;
    rom[11790] = 25'b1111111111001010001110100;
    rom[11791] = 25'b1111111111001010001011010;
    rom[11792] = 25'b1111111111001010001000001;
    rom[11793] = 25'b1111111111001010000101000;
    rom[11794] = 25'b1111111111001010000001111;
    rom[11795] = 25'b1111111111001001111110110;
    rom[11796] = 25'b1111111111001001111011101;
    rom[11797] = 25'b1111111111001001111000100;
    rom[11798] = 25'b1111111111001001110101011;
    rom[11799] = 25'b1111111111001001110010011;
    rom[11800] = 25'b1111111111001001101111001;
    rom[11801] = 25'b1111111111001001101100001;
    rom[11802] = 25'b1111111111001001101001000;
    rom[11803] = 25'b1111111111001001100101111;
    rom[11804] = 25'b1111111111001001100010110;
    rom[11805] = 25'b1111111111001001011111101;
    rom[11806] = 25'b1111111111001001011100101;
    rom[11807] = 25'b1111111111001001011001100;
    rom[11808] = 25'b1111111111001001010110011;
    rom[11809] = 25'b1111111111001001010011011;
    rom[11810] = 25'b1111111111001001010000010;
    rom[11811] = 25'b1111111111001001001101001;
    rom[11812] = 25'b1111111111001001001010001;
    rom[11813] = 25'b1111111111001001000111000;
    rom[11814] = 25'b1111111111001001000011111;
    rom[11815] = 25'b1111111111001001000000111;
    rom[11816] = 25'b1111111111001000111101110;
    rom[11817] = 25'b1111111111001000111010110;
    rom[11818] = 25'b1111111111001000110111101;
    rom[11819] = 25'b1111111111001000110100101;
    rom[11820] = 25'b1111111111001000110001100;
    rom[11821] = 25'b1111111111001000101110100;
    rom[11822] = 25'b1111111111001000101011100;
    rom[11823] = 25'b1111111111001000101000100;
    rom[11824] = 25'b1111111111001000100101011;
    rom[11825] = 25'b1111111111001000100010011;
    rom[11826] = 25'b1111111111001000011111010;
    rom[11827] = 25'b1111111111001000011100011;
    rom[11828] = 25'b1111111111001000011001010;
    rom[11829] = 25'b1111111111001000010110010;
    rom[11830] = 25'b1111111111001000010011001;
    rom[11831] = 25'b1111111111001000010000001;
    rom[11832] = 25'b1111111111001000001101010;
    rom[11833] = 25'b1111111111001000001010010;
    rom[11834] = 25'b1111111111001000000111001;
    rom[11835] = 25'b1111111111001000000100001;
    rom[11836] = 25'b1111111111001000000001001;
    rom[11837] = 25'b1111111111000111111110001;
    rom[11838] = 25'b1111111111000111111011001;
    rom[11839] = 25'b1111111111000111111000001;
    rom[11840] = 25'b1111111111000111110101010;
    rom[11841] = 25'b1111111111000111110010010;
    rom[11842] = 25'b1111111111000111101111010;
    rom[11843] = 25'b1111111111000111101100010;
    rom[11844] = 25'b1111111111000111101001010;
    rom[11845] = 25'b1111111111000111100110010;
    rom[11846] = 25'b1111111111000111100011011;
    rom[11847] = 25'b1111111111000111100000011;
    rom[11848] = 25'b1111111111000111011101011;
    rom[11849] = 25'b1111111111000111011010011;
    rom[11850] = 25'b1111111111000111010111100;
    rom[11851] = 25'b1111111111000111010100100;
    rom[11852] = 25'b1111111111000111010001101;
    rom[11853] = 25'b1111111111000111001110101;
    rom[11854] = 25'b1111111111000111001011101;
    rom[11855] = 25'b1111111111000111001000110;
    rom[11856] = 25'b1111111111000111000101111;
    rom[11857] = 25'b1111111111000111000010111;
    rom[11858] = 25'b1111111111000111000000000;
    rom[11859] = 25'b1111111111000110111101000;
    rom[11860] = 25'b1111111111000110111010001;
    rom[11861] = 25'b1111111111000110110111001;
    rom[11862] = 25'b1111111111000110110100010;
    rom[11863] = 25'b1111111111000110110001010;
    rom[11864] = 25'b1111111111000110101110011;
    rom[11865] = 25'b1111111111000110101011100;
    rom[11866] = 25'b1111111111000110101000101;
    rom[11867] = 25'b1111111111000110100101110;
    rom[11868] = 25'b1111111111000110100010111;
    rom[11869] = 25'b1111111111000110011111111;
    rom[11870] = 25'b1111111111000110011101000;
    rom[11871] = 25'b1111111111000110011010001;
    rom[11872] = 25'b1111111111000110010111010;
    rom[11873] = 25'b1111111111000110010100100;
    rom[11874] = 25'b1111111111000110010001100;
    rom[11875] = 25'b1111111111000110001110101;
    rom[11876] = 25'b1111111111000110001011110;
    rom[11877] = 25'b1111111111000110001001000;
    rom[11878] = 25'b1111111111000110000110000;
    rom[11879] = 25'b1111111111000110000011001;
    rom[11880] = 25'b1111111111000110000000011;
    rom[11881] = 25'b1111111111000101111101100;
    rom[11882] = 25'b1111111111000101111010101;
    rom[11883] = 25'b1111111111000101110111110;
    rom[11884] = 25'b1111111111000101110101000;
    rom[11885] = 25'b1111111111000101110010001;
    rom[11886] = 25'b1111111111000101101111010;
    rom[11887] = 25'b1111111111000101101100100;
    rom[11888] = 25'b1111111111000101101001101;
    rom[11889] = 25'b1111111111000101100110110;
    rom[11890] = 25'b1111111111000101100100000;
    rom[11891] = 25'b1111111111000101100001001;
    rom[11892] = 25'b1111111111000101011110011;
    rom[11893] = 25'b1111111111000101011011101;
    rom[11894] = 25'b1111111111000101011000110;
    rom[11895] = 25'b1111111111000101010110000;
    rom[11896] = 25'b1111111111000101010011001;
    rom[11897] = 25'b1111111111000101010000011;
    rom[11898] = 25'b1111111111000101001101100;
    rom[11899] = 25'b1111111111000101001010110;
    rom[11900] = 25'b1111111111000101001000000;
    rom[11901] = 25'b1111111111000101000101010;
    rom[11902] = 25'b1111111111000101000010100;
    rom[11903] = 25'b1111111111000100111111101;
    rom[11904] = 25'b1111111111000100111101000;
    rom[11905] = 25'b1111111111000100111010001;
    rom[11906] = 25'b1111111111000100110111011;
    rom[11907] = 25'b1111111111000100110100101;
    rom[11908] = 25'b1111111111000100110001111;
    rom[11909] = 25'b1111111111000100101111001;
    rom[11910] = 25'b1111111111000100101100011;
    rom[11911] = 25'b1111111111000100101001101;
    rom[11912] = 25'b1111111111000100100110111;
    rom[11913] = 25'b1111111111000100100100001;
    rom[11914] = 25'b1111111111000100100001011;
    rom[11915] = 25'b1111111111000100011110101;
    rom[11916] = 25'b1111111111000100011100000;
    rom[11917] = 25'b1111111111000100011001010;
    rom[11918] = 25'b1111111111000100010110100;
    rom[11919] = 25'b1111111111000100010011110;
    rom[11920] = 25'b1111111111000100010001000;
    rom[11921] = 25'b1111111111000100001110011;
    rom[11922] = 25'b1111111111000100001011101;
    rom[11923] = 25'b1111111111000100001001000;
    rom[11924] = 25'b1111111111000100000110010;
    rom[11925] = 25'b1111111111000100000011101;
    rom[11926] = 25'b1111111111000100000000111;
    rom[11927] = 25'b1111111111000011111110001;
    rom[11928] = 25'b1111111111000011111011101;
    rom[11929] = 25'b1111111111000011111000111;
    rom[11930] = 25'b1111111111000011110110001;
    rom[11931] = 25'b1111111111000011110011100;
    rom[11932] = 25'b1111111111000011110000111;
    rom[11933] = 25'b1111111111000011101110010;
    rom[11934] = 25'b1111111111000011101011100;
    rom[11935] = 25'b1111111111000011101000111;
    rom[11936] = 25'b1111111111000011100110010;
    rom[11937] = 25'b1111111111000011100011101;
    rom[11938] = 25'b1111111111000011100001000;
    rom[11939] = 25'b1111111111000011011110011;
    rom[11940] = 25'b1111111111000011011011101;
    rom[11941] = 25'b1111111111000011011001000;
    rom[11942] = 25'b1111111111000011010110011;
    rom[11943] = 25'b1111111111000011010011110;
    rom[11944] = 25'b1111111111000011010001001;
    rom[11945] = 25'b1111111111000011001110100;
    rom[11946] = 25'b1111111111000011001100000;
    rom[11947] = 25'b1111111111000011001001011;
    rom[11948] = 25'b1111111111000011000110110;
    rom[11949] = 25'b1111111111000011000100001;
    rom[11950] = 25'b1111111111000011000001101;
    rom[11951] = 25'b1111111111000010111111000;
    rom[11952] = 25'b1111111111000010111100011;
    rom[11953] = 25'b1111111111000010111001110;
    rom[11954] = 25'b1111111111000010110111010;
    rom[11955] = 25'b1111111111000010110100101;
    rom[11956] = 25'b1111111111000010110010001;
    rom[11957] = 25'b1111111111000010101111100;
    rom[11958] = 25'b1111111111000010101100111;
    rom[11959] = 25'b1111111111000010101010011;
    rom[11960] = 25'b1111111111000010100111110;
    rom[11961] = 25'b1111111111000010100101010;
    rom[11962] = 25'b1111111111000010100010101;
    rom[11963] = 25'b1111111111000010100000001;
    rom[11964] = 25'b1111111111000010011101101;
    rom[11965] = 25'b1111111111000010011011001;
    rom[11966] = 25'b1111111111000010011000101;
    rom[11967] = 25'b1111111111000010010110000;
    rom[11968] = 25'b1111111111000010010011100;
    rom[11969] = 25'b1111111111000010010001000;
    rom[11970] = 25'b1111111111000010001110100;
    rom[11971] = 25'b1111111111000010001100000;
    rom[11972] = 25'b1111111111000010001001100;
    rom[11973] = 25'b1111111111000010000110111;
    rom[11974] = 25'b1111111111000010000100011;
    rom[11975] = 25'b1111111111000010000010000;
    rom[11976] = 25'b1111111111000001111111100;
    rom[11977] = 25'b1111111111000001111100111;
    rom[11978] = 25'b1111111111000001111010100;
    rom[11979] = 25'b1111111111000001111000000;
    rom[11980] = 25'b1111111111000001110101100;
    rom[11981] = 25'b1111111111000001110011000;
    rom[11982] = 25'b1111111111000001110000101;
    rom[11983] = 25'b1111111111000001101110001;
    rom[11984] = 25'b1111111111000001101011101;
    rom[11985] = 25'b1111111111000001101001010;
    rom[11986] = 25'b1111111111000001100110110;
    rom[11987] = 25'b1111111111000001100100010;
    rom[11988] = 25'b1111111111000001100001111;
    rom[11989] = 25'b1111111111000001011111011;
    rom[11990] = 25'b1111111111000001011101000;
    rom[11991] = 25'b1111111111000001011010101;
    rom[11992] = 25'b1111111111000001011000001;
    rom[11993] = 25'b1111111111000001010101110;
    rom[11994] = 25'b1111111111000001010011010;
    rom[11995] = 25'b1111111111000001010000111;
    rom[11996] = 25'b1111111111000001001110011;
    rom[11997] = 25'b1111111111000001001100001;
    rom[11998] = 25'b1111111111000001001001101;
    rom[11999] = 25'b1111111111000001000111010;
    rom[12000] = 25'b1111111111000001000100111;
    rom[12001] = 25'b1111111111000001000010100;
    rom[12002] = 25'b1111111111000001000000001;
    rom[12003] = 25'b1111111111000000111101110;
    rom[12004] = 25'b1111111111000000111011011;
    rom[12005] = 25'b1111111111000000111001000;
    rom[12006] = 25'b1111111111000000110110101;
    rom[12007] = 25'b1111111111000000110100010;
    rom[12008] = 25'b1111111111000000110001111;
    rom[12009] = 25'b1111111111000000101111100;
    rom[12010] = 25'b1111111111000000101101001;
    rom[12011] = 25'b1111111111000000101010111;
    rom[12012] = 25'b1111111111000000101000100;
    rom[12013] = 25'b1111111111000000100110001;
    rom[12014] = 25'b1111111111000000100011111;
    rom[12015] = 25'b1111111111000000100001100;
    rom[12016] = 25'b1111111111000000011111001;
    rom[12017] = 25'b1111111111000000011100111;
    rom[12018] = 25'b1111111111000000011010100;
    rom[12019] = 25'b1111111111000000011000010;
    rom[12020] = 25'b1111111111000000010101111;
    rom[12021] = 25'b1111111111000000010011101;
    rom[12022] = 25'b1111111111000000010001011;
    rom[12023] = 25'b1111111111000000001111000;
    rom[12024] = 25'b1111111111000000001100110;
    rom[12025] = 25'b1111111111000000001010100;
    rom[12026] = 25'b1111111111000000001000010;
    rom[12027] = 25'b1111111111000000000101111;
    rom[12028] = 25'b1111111111000000000011101;
    rom[12029] = 25'b1111111111000000000001011;
    rom[12030] = 25'b1111111110111111111111001;
    rom[12031] = 25'b1111111110111111111100110;
    rom[12032] = 25'b1111111110111111111010101;
    rom[12033] = 25'b1111111110111111111000011;
    rom[12034] = 25'b1111111110111111110110001;
    rom[12035] = 25'b1111111110111111110011111;
    rom[12036] = 25'b1111111110111111110001101;
    rom[12037] = 25'b1111111110111111101111011;
    rom[12038] = 25'b1111111110111111101101010;
    rom[12039] = 25'b1111111110111111101011000;
    rom[12040] = 25'b1111111110111111101000110;
    rom[12041] = 25'b1111111110111111100110100;
    rom[12042] = 25'b1111111110111111100100011;
    rom[12043] = 25'b1111111110111111100010001;
    rom[12044] = 25'b1111111110111111011111111;
    rom[12045] = 25'b1111111110111111011101110;
    rom[12046] = 25'b1111111110111111011011100;
    rom[12047] = 25'b1111111110111111011001011;
    rom[12048] = 25'b1111111110111111010111001;
    rom[12049] = 25'b1111111110111111010100111;
    rom[12050] = 25'b1111111110111111010010110;
    rom[12051] = 25'b1111111110111111010000101;
    rom[12052] = 25'b1111111110111111001110100;
    rom[12053] = 25'b1111111110111111001100011;
    rom[12054] = 25'b1111111110111111001010001;
    rom[12055] = 25'b1111111110111111001000000;
    rom[12056] = 25'b1111111110111111000101110;
    rom[12057] = 25'b1111111110111111000011101;
    rom[12058] = 25'b1111111110111111000001101;
    rom[12059] = 25'b1111111110111110111111100;
    rom[12060] = 25'b1111111110111110111101010;
    rom[12061] = 25'b1111111110111110111011001;
    rom[12062] = 25'b1111111110111110111001001;
    rom[12063] = 25'b1111111110111110110111000;
    rom[12064] = 25'b1111111110111110110100110;
    rom[12065] = 25'b1111111110111110110010110;
    rom[12066] = 25'b1111111110111110110000101;
    rom[12067] = 25'b1111111110111110101110100;
    rom[12068] = 25'b1111111110111110101100011;
    rom[12069] = 25'b1111111110111110101010011;
    rom[12070] = 25'b1111111110111110101000010;
    rom[12071] = 25'b1111111110111110100110010;
    rom[12072] = 25'b1111111110111110100100001;
    rom[12073] = 25'b1111111110111110100010000;
    rom[12074] = 25'b1111111110111110100000000;
    rom[12075] = 25'b1111111110111110011101111;
    rom[12076] = 25'b1111111110111110011011111;
    rom[12077] = 25'b1111111110111110011001111;
    rom[12078] = 25'b1111111110111110010111110;
    rom[12079] = 25'b1111111110111110010101110;
    rom[12080] = 25'b1111111110111110010011110;
    rom[12081] = 25'b1111111110111110010001110;
    rom[12082] = 25'b1111111110111110001111101;
    rom[12083] = 25'b1111111110111110001101101;
    rom[12084] = 25'b1111111110111110001011101;
    rom[12085] = 25'b1111111110111110001001101;
    rom[12086] = 25'b1111111110111110000111101;
    rom[12087] = 25'b1111111110111110000101101;
    rom[12088] = 25'b1111111110111110000011101;
    rom[12089] = 25'b1111111110111110000001101;
    rom[12090] = 25'b1111111110111101111111101;
    rom[12091] = 25'b1111111110111101111101101;
    rom[12092] = 25'b1111111110111101111011101;
    rom[12093] = 25'b1111111110111101111001110;
    rom[12094] = 25'b1111111110111101110111110;
    rom[12095] = 25'b1111111110111101110101110;
    rom[12096] = 25'b1111111110111101110011110;
    rom[12097] = 25'b1111111110111101110001111;
    rom[12098] = 25'b1111111110111101101111111;
    rom[12099] = 25'b1111111110111101101101111;
    rom[12100] = 25'b1111111110111101101100000;
    rom[12101] = 25'b1111111110111101101010001;
    rom[12102] = 25'b1111111110111101101000001;
    rom[12103] = 25'b1111111110111101100110001;
    rom[12104] = 25'b1111111110111101100100010;
    rom[12105] = 25'b1111111110111101100010011;
    rom[12106] = 25'b1111111110111101100000100;
    rom[12107] = 25'b1111111110111101011110101;
    rom[12108] = 25'b1111111110111101011100101;
    rom[12109] = 25'b1111111110111101011010110;
    rom[12110] = 25'b1111111110111101011000111;
    rom[12111] = 25'b1111111110111101010111000;
    rom[12112] = 25'b1111111110111101010101001;
    rom[12113] = 25'b1111111110111101010011010;
    rom[12114] = 25'b1111111110111101010001011;
    rom[12115] = 25'b1111111110111101001111100;
    rom[12116] = 25'b1111111110111101001101101;
    rom[12117] = 25'b1111111110111101001011110;
    rom[12118] = 25'b1111111110111101001001111;
    rom[12119] = 25'b1111111110111101001000001;
    rom[12120] = 25'b1111111110111101000110010;
    rom[12121] = 25'b1111111110111101000100011;
    rom[12122] = 25'b1111111110111101000010101;
    rom[12123] = 25'b1111111110111101000000110;
    rom[12124] = 25'b1111111110111100111111000;
    rom[12125] = 25'b1111111110111100111101001;
    rom[12126] = 25'b1111111110111100111011010;
    rom[12127] = 25'b1111111110111100111001100;
    rom[12128] = 25'b1111111110111100110111101;
    rom[12129] = 25'b1111111110111100110101111;
    rom[12130] = 25'b1111111110111100110100001;
    rom[12131] = 25'b1111111110111100110010010;
    rom[12132] = 25'b1111111110111100110000100;
    rom[12133] = 25'b1111111110111100101110110;
    rom[12134] = 25'b1111111110111100101100111;
    rom[12135] = 25'b1111111110111100101011001;
    rom[12136] = 25'b1111111110111100101001100;
    rom[12137] = 25'b1111111110111100100111110;
    rom[12138] = 25'b1111111110111100100101111;
    rom[12139] = 25'b1111111110111100100100001;
    rom[12140] = 25'b1111111110111100100010100;
    rom[12141] = 25'b1111111110111100100000110;
    rom[12142] = 25'b1111111110111100011110111;
    rom[12143] = 25'b1111111110111100011101010;
    rom[12144] = 25'b1111111110111100011011100;
    rom[12145] = 25'b1111111110111100011001110;
    rom[12146] = 25'b1111111110111100011000001;
    rom[12147] = 25'b1111111110111100010110011;
    rom[12148] = 25'b1111111110111100010100101;
    rom[12149] = 25'b1111111110111100010011000;
    rom[12150] = 25'b1111111110111100010001010;
    rom[12151] = 25'b1111111110111100001111101;
    rom[12152] = 25'b1111111110111100001101111;
    rom[12153] = 25'b1111111110111100001100010;
    rom[12154] = 25'b1111111110111100001010100;
    rom[12155] = 25'b1111111110111100001000111;
    rom[12156] = 25'b1111111110111100000111010;
    rom[12157] = 25'b1111111110111100000101101;
    rom[12158] = 25'b1111111110111100000011111;
    rom[12159] = 25'b1111111110111100000010010;
    rom[12160] = 25'b1111111110111100000000101;
    rom[12161] = 25'b1111111110111011111111000;
    rom[12162] = 25'b1111111110111011111101011;
    rom[12163] = 25'b1111111110111011111011110;
    rom[12164] = 25'b1111111110111011111010001;
    rom[12165] = 25'b1111111110111011111000100;
    rom[12166] = 25'b1111111110111011110111000;
    rom[12167] = 25'b1111111110111011110101010;
    rom[12168] = 25'b1111111110111011110011101;
    rom[12169] = 25'b1111111110111011110010001;
    rom[12170] = 25'b1111111110111011110000100;
    rom[12171] = 25'b1111111110111011101110111;
    rom[12172] = 25'b1111111110111011101101011;
    rom[12173] = 25'b1111111110111011101011111;
    rom[12174] = 25'b1111111110111011101010010;
    rom[12175] = 25'b1111111110111011101000101;
    rom[12176] = 25'b1111111110111011100111001;
    rom[12177] = 25'b1111111110111011100101101;
    rom[12178] = 25'b1111111110111011100100000;
    rom[12179] = 25'b1111111110111011100010100;
    rom[12180] = 25'b1111111110111011100000111;
    rom[12181] = 25'b1111111110111011011111011;
    rom[12182] = 25'b1111111110111011011101111;
    rom[12183] = 25'b1111111110111011011100011;
    rom[12184] = 25'b1111111110111011011010111;
    rom[12185] = 25'b1111111110111011011001011;
    rom[12186] = 25'b1111111110111011010111111;
    rom[12187] = 25'b1111111110111011010110011;
    rom[12188] = 25'b1111111110111011010100111;
    rom[12189] = 25'b1111111110111011010011011;
    rom[12190] = 25'b1111111110111011010001111;
    rom[12191] = 25'b1111111110111011010000011;
    rom[12192] = 25'b1111111110111011001110111;
    rom[12193] = 25'b1111111110111011001101100;
    rom[12194] = 25'b1111111110111011001100000;
    rom[12195] = 25'b1111111110111011001010100;
    rom[12196] = 25'b1111111110111011001001001;
    rom[12197] = 25'b1111111110111011000111101;
    rom[12198] = 25'b1111111110111011000110010;
    rom[12199] = 25'b1111111110111011000100110;
    rom[12200] = 25'b1111111110111011000011010;
    rom[12201] = 25'b1111111110111011000001111;
    rom[12202] = 25'b1111111110111011000000100;
    rom[12203] = 25'b1111111110111010111111001;
    rom[12204] = 25'b1111111110111010111101101;
    rom[12205] = 25'b1111111110111010111100010;
    rom[12206] = 25'b1111111110111010111010111;
    rom[12207] = 25'b1111111110111010111001100;
    rom[12208] = 25'b1111111110111010111000001;
    rom[12209] = 25'b1111111110111010110110110;
    rom[12210] = 25'b1111111110111010110101010;
    rom[12211] = 25'b1111111110111010110100000;
    rom[12212] = 25'b1111111110111010110010101;
    rom[12213] = 25'b1111111110111010110001010;
    rom[12214] = 25'b1111111110111010101111111;
    rom[12215] = 25'b1111111110111010101110100;
    rom[12216] = 25'b1111111110111010101101001;
    rom[12217] = 25'b1111111110111010101011111;
    rom[12218] = 25'b1111111110111010101010100;
    rom[12219] = 25'b1111111110111010101001001;
    rom[12220] = 25'b1111111110111010100111111;
    rom[12221] = 25'b1111111110111010100110100;
    rom[12222] = 25'b1111111110111010100101010;
    rom[12223] = 25'b1111111110111010100011111;
    rom[12224] = 25'b1111111110111010100010101;
    rom[12225] = 25'b1111111110111010100001011;
    rom[12226] = 25'b1111111110111010100000000;
    rom[12227] = 25'b1111111110111010011110110;
    rom[12228] = 25'b1111111110111010011101100;
    rom[12229] = 25'b1111111110111010011100001;
    rom[12230] = 25'b1111111110111010011011000;
    rom[12231] = 25'b1111111110111010011001101;
    rom[12232] = 25'b1111111110111010011000100;
    rom[12233] = 25'b1111111110111010010111010;
    rom[12234] = 25'b1111111110111010010101111;
    rom[12235] = 25'b1111111110111010010100110;
    rom[12236] = 25'b1111111110111010010011100;
    rom[12237] = 25'b1111111110111010010010010;
    rom[12238] = 25'b1111111110111010010001001;
    rom[12239] = 25'b1111111110111010001111111;
    rom[12240] = 25'b1111111110111010001110101;
    rom[12241] = 25'b1111111110111010001101011;
    rom[12242] = 25'b1111111110111010001100010;
    rom[12243] = 25'b1111111110111010001011000;
    rom[12244] = 25'b1111111110111010001001110;
    rom[12245] = 25'b1111111110111010001000101;
    rom[12246] = 25'b1111111110111010000111100;
    rom[12247] = 25'b1111111110111010000110011;
    rom[12248] = 25'b1111111110111010000101001;
    rom[12249] = 25'b1111111110111010000100000;
    rom[12250] = 25'b1111111110111010000010110;
    rom[12251] = 25'b1111111110111010000001101;
    rom[12252] = 25'b1111111110111010000000100;
    rom[12253] = 25'b1111111110111001111111011;
    rom[12254] = 25'b1111111110111001111110010;
    rom[12255] = 25'b1111111110111001111101001;
    rom[12256] = 25'b1111111110111001111100000;
    rom[12257] = 25'b1111111110111001111010111;
    rom[12258] = 25'b1111111110111001111001110;
    rom[12259] = 25'b1111111110111001111000110;
    rom[12260] = 25'b1111111110111001110111101;
    rom[12261] = 25'b1111111110111001110110100;
    rom[12262] = 25'b1111111110111001110101011;
    rom[12263] = 25'b1111111110111001110100010;
    rom[12264] = 25'b1111111110111001110011010;
    rom[12265] = 25'b1111111110111001110010001;
    rom[12266] = 25'b1111111110111001110001001;
    rom[12267] = 25'b1111111110111001110000001;
    rom[12268] = 25'b1111111110111001101111000;
    rom[12269] = 25'b1111111110111001101110000;
    rom[12270] = 25'b1111111110111001101100111;
    rom[12271] = 25'b1111111110111001101011111;
    rom[12272] = 25'b1111111110111001101010111;
    rom[12273] = 25'b1111111110111001101001111;
    rom[12274] = 25'b1111111110111001101000111;
    rom[12275] = 25'b1111111110111001100111110;
    rom[12276] = 25'b1111111110111001100110110;
    rom[12277] = 25'b1111111110111001100101111;
    rom[12278] = 25'b1111111110111001100100110;
    rom[12279] = 25'b1111111110111001100011110;
    rom[12280] = 25'b1111111110111001100010111;
    rom[12281] = 25'b1111111110111001100001110;
    rom[12282] = 25'b1111111110111001100000111;
    rom[12283] = 25'b1111111110111001100000000;
    rom[12284] = 25'b1111111110111001011110111;
    rom[12285] = 25'b1111111110111001011110000;
    rom[12286] = 25'b1111111110111001011101000;
    rom[12287] = 25'b1111111110111001011100001;
    rom[12288] = 25'b1111111110111001011011001;
    rom[12289] = 25'b1111111110111001011010010;
    rom[12290] = 25'b1111111110111001011001011;
    rom[12291] = 25'b1111111110111001011000011;
    rom[12292] = 25'b1111111110111001010111100;
    rom[12293] = 25'b1111111110111001010110101;
    rom[12294] = 25'b1111111110111001010101101;
    rom[12295] = 25'b1111111110111001010100111;
    rom[12296] = 25'b1111111110111001010011111;
    rom[12297] = 25'b1111111110111001010011000;
    rom[12298] = 25'b1111111110111001010010001;
    rom[12299] = 25'b1111111110111001010001010;
    rom[12300] = 25'b1111111110111001010000100;
    rom[12301] = 25'b1111111110111001001111100;
    rom[12302] = 25'b1111111110111001001110101;
    rom[12303] = 25'b1111111110111001001101111;
    rom[12304] = 25'b1111111110111001001101000;
    rom[12305] = 25'b1111111110111001001100001;
    rom[12306] = 25'b1111111110111001001011010;
    rom[12307] = 25'b1111111110111001001010100;
    rom[12308] = 25'b1111111110111001001001110;
    rom[12309] = 25'b1111111110111001001000111;
    rom[12310] = 25'b1111111110111001001000000;
    rom[12311] = 25'b1111111110111001000111010;
    rom[12312] = 25'b1111111110111001000110100;
    rom[12313] = 25'b1111111110111001000101110;
    rom[12314] = 25'b1111111110111001000100111;
    rom[12315] = 25'b1111111110111001000100001;
    rom[12316] = 25'b1111111110111001000011011;
    rom[12317] = 25'b1111111110111001000010101;
    rom[12318] = 25'b1111111110111001000001111;
    rom[12319] = 25'b1111111110111001000001000;
    rom[12320] = 25'b1111111110111001000000011;
    rom[12321] = 25'b1111111110111000111111101;
    rom[12322] = 25'b1111111110111000111110111;
    rom[12323] = 25'b1111111110111000111110001;
    rom[12324] = 25'b1111111110111000111101011;
    rom[12325] = 25'b1111111110111000111100101;
    rom[12326] = 25'b1111111110111000111100000;
    rom[12327] = 25'b1111111110111000111011010;
    rom[12328] = 25'b1111111110111000111010101;
    rom[12329] = 25'b1111111110111000111001111;
    rom[12330] = 25'b1111111110111000111001010;
    rom[12331] = 25'b1111111110111000111000100;
    rom[12332] = 25'b1111111110111000110111111;
    rom[12333] = 25'b1111111110111000110111001;
    rom[12334] = 25'b1111111110111000110110100;
    rom[12335] = 25'b1111111110111000110101111;
    rom[12336] = 25'b1111111110111000110101001;
    rom[12337] = 25'b1111111110111000110100100;
    rom[12338] = 25'b1111111110111000110100000;
    rom[12339] = 25'b1111111110111000110011010;
    rom[12340] = 25'b1111111110111000110010101;
    rom[12341] = 25'b1111111110111000110010000;
    rom[12342] = 25'b1111111110111000110001011;
    rom[12343] = 25'b1111111110111000110000110;
    rom[12344] = 25'b1111111110111000110000010;
    rom[12345] = 25'b1111111110111000101111101;
    rom[12346] = 25'b1111111110111000101111000;
    rom[12347] = 25'b1111111110111000101110100;
    rom[12348] = 25'b1111111110111000101101111;
    rom[12349] = 25'b1111111110111000101101011;
    rom[12350] = 25'b1111111110111000101100110;
    rom[12351] = 25'b1111111110111000101100010;
    rom[12352] = 25'b1111111110111000101011101;
    rom[12353] = 25'b1111111110111000101011001;
    rom[12354] = 25'b1111111110111000101010100;
    rom[12355] = 25'b1111111110111000101010000;
    rom[12356] = 25'b1111111110111000101001100;
    rom[12357] = 25'b1111111110111000101001000;
    rom[12358] = 25'b1111111110111000101000100;
    rom[12359] = 25'b1111111110111000100111111;
    rom[12360] = 25'b1111111110111000100111100;
    rom[12361] = 25'b1111111110111000100110111;
    rom[12362] = 25'b1111111110111000100110011;
    rom[12363] = 25'b1111111110111000100110000;
    rom[12364] = 25'b1111111110111000100101100;
    rom[12365] = 25'b1111111110111000100101000;
    rom[12366] = 25'b1111111110111000100100100;
    rom[12367] = 25'b1111111110111000100100001;
    rom[12368] = 25'b1111111110111000100011101;
    rom[12369] = 25'b1111111110111000100011001;
    rom[12370] = 25'b1111111110111000100010101;
    rom[12371] = 25'b1111111110111000100010010;
    rom[12372] = 25'b1111111110111000100001111;
    rom[12373] = 25'b1111111110111000100001100;
    rom[12374] = 25'b1111111110111000100001000;
    rom[12375] = 25'b1111111110111000100000101;
    rom[12376] = 25'b1111111110111000100000001;
    rom[12377] = 25'b1111111110111000011111110;
    rom[12378] = 25'b1111111110111000011111011;
    rom[12379] = 25'b1111111110111000011111000;
    rom[12380] = 25'b1111111110111000011110101;
    rom[12381] = 25'b1111111110111000011110010;
    rom[12382] = 25'b1111111110111000011101111;
    rom[12383] = 25'b1111111110111000011101100;
    rom[12384] = 25'b1111111110111000011101001;
    rom[12385] = 25'b1111111110111000011100111;
    rom[12386] = 25'b1111111110111000011100100;
    rom[12387] = 25'b1111111110111000011100001;
    rom[12388] = 25'b1111111110111000011011111;
    rom[12389] = 25'b1111111110111000011011100;
    rom[12390] = 25'b1111111110111000011011010;
    rom[12391] = 25'b1111111110111000011010111;
    rom[12392] = 25'b1111111110111000011010100;
    rom[12393] = 25'b1111111110111000011010010;
    rom[12394] = 25'b1111111110111000011010000;
    rom[12395] = 25'b1111111110111000011001110;
    rom[12396] = 25'b1111111110111000011001011;
    rom[12397] = 25'b1111111110111000011001001;
    rom[12398] = 25'b1111111110111000011000111;
    rom[12399] = 25'b1111111110111000011000110;
    rom[12400] = 25'b1111111110111000011000011;
    rom[12401] = 25'b1111111110111000011000001;
    rom[12402] = 25'b1111111110111000011000000;
    rom[12403] = 25'b1111111110111000010111101;
    rom[12404] = 25'b1111111110111000010111100;
    rom[12405] = 25'b1111111110111000010111010;
    rom[12406] = 25'b1111111110111000010111000;
    rom[12407] = 25'b1111111110111000010110111;
    rom[12408] = 25'b1111111110111000010110101;
    rom[12409] = 25'b1111111110111000010110011;
    rom[12410] = 25'b1111111110111000010110001;
    rom[12411] = 25'b1111111110111000010110000;
    rom[12412] = 25'b1111111110111000010101111;
    rom[12413] = 25'b1111111110111000010101110;
    rom[12414] = 25'b1111111110111000010101100;
    rom[12415] = 25'b1111111110111000010101011;
    rom[12416] = 25'b1111111110111000010101010;
    rom[12417] = 25'b1111111110111000010101000;
    rom[12418] = 25'b1111111110111000010101000;
    rom[12419] = 25'b1111111110111000010100110;
    rom[12420] = 25'b1111111110111000010100101;
    rom[12421] = 25'b1111111110111000010100101;
    rom[12422] = 25'b1111111110111000010100011;
    rom[12423] = 25'b1111111110111000010100010;
    rom[12424] = 25'b1111111110111000010100010;
    rom[12425] = 25'b1111111110111000010100001;
    rom[12426] = 25'b1111111110111000010100000;
    rom[12427] = 25'b1111111110111000010100000;
    rom[12428] = 25'b1111111110111000010011111;
    rom[12429] = 25'b1111111110111000010011111;
    rom[12430] = 25'b1111111110111000010011110;
    rom[12431] = 25'b1111111110111000010011110;
    rom[12432] = 25'b1111111110111000010011101;
    rom[12433] = 25'b1111111110111000010011101;
    rom[12434] = 25'b1111111110111000010011100;
    rom[12435] = 25'b1111111110111000010011100;
    rom[12436] = 25'b1111111110111000010011100;
    rom[12437] = 25'b1111111110111000010011100;
    rom[12438] = 25'b1111111110111000010011100;
    rom[12439] = 25'b1111111110111000010011100;
    rom[12440] = 25'b1111111110111000010011100;
    rom[12441] = 25'b1111111110111000010011100;
    rom[12442] = 25'b1111111110111000010011100;
    rom[12443] = 25'b1111111110111000010011100;
    rom[12444] = 25'b1111111110111000010011101;
    rom[12445] = 25'b1111111110111000010011101;
    rom[12446] = 25'b1111111110111000010011101;
    rom[12447] = 25'b1111111110111000010011110;
    rom[12448] = 25'b1111111110111000010011111;
    rom[12449] = 25'b1111111110111000010011111;
    rom[12450] = 25'b1111111110111000010011111;
    rom[12451] = 25'b1111111110111000010100000;
    rom[12452] = 25'b1111111110111000010100001;
    rom[12453] = 25'b1111111110111000010100010;
    rom[12454] = 25'b1111111110111000010100010;
    rom[12455] = 25'b1111111110111000010100011;
    rom[12456] = 25'b1111111110111000010100100;
    rom[12457] = 25'b1111111110111000010100101;
    rom[12458] = 25'b1111111110111000010100110;
    rom[12459] = 25'b1111111110111000010100111;
    rom[12460] = 25'b1111111110111000010101000;
    rom[12461] = 25'b1111111110111000010101001;
    rom[12462] = 25'b1111111110111000010101010;
    rom[12463] = 25'b1111111110111000010101011;
    rom[12464] = 25'b1111111110111000010101101;
    rom[12465] = 25'b1111111110111000010101110;
    rom[12466] = 25'b1111111110111000010110000;
    rom[12467] = 25'b1111111110111000010110001;
    rom[12468] = 25'b1111111110111000010110011;
    rom[12469] = 25'b1111111110111000010110100;
    rom[12470] = 25'b1111111110111000010110110;
    rom[12471] = 25'b1111111110111000010110111;
    rom[12472] = 25'b1111111110111000010111001;
    rom[12473] = 25'b1111111110111000010111011;
    rom[12474] = 25'b1111111110111000010111101;
    rom[12475] = 25'b1111111110111000010111111;
    rom[12476] = 25'b1111111110111000011000000;
    rom[12477] = 25'b1111111110111000011000011;
    rom[12478] = 25'b1111111110111000011000101;
    rom[12479] = 25'b1111111110111000011000110;
    rom[12480] = 25'b1111111110111000011001001;
    rom[12481] = 25'b1111111110111000011001011;
    rom[12482] = 25'b1111111110111000011001101;
    rom[12483] = 25'b1111111110111000011001111;
    rom[12484] = 25'b1111111110111000011010010;
    rom[12485] = 25'b1111111110111000011010100;
    rom[12486] = 25'b1111111110111000011010111;
    rom[12487] = 25'b1111111110111000011011001;
    rom[12488] = 25'b1111111110111000011011100;
    rom[12489] = 25'b1111111110111000011011110;
    rom[12490] = 25'b1111111110111000011100001;
    rom[12491] = 25'b1111111110111000011100100;
    rom[12492] = 25'b1111111110111000011100110;
    rom[12493] = 25'b1111111110111000011101001;
    rom[12494] = 25'b1111111110111000011101100;
    rom[12495] = 25'b1111111110111000011101111;
    rom[12496] = 25'b1111111110111000011110010;
    rom[12497] = 25'b1111111110111000011110101;
    rom[12498] = 25'b1111111110111000011111000;
    rom[12499] = 25'b1111111110111000011111011;
    rom[12500] = 25'b1111111110111000011111111;
    rom[12501] = 25'b1111111110111000100000010;
    rom[12502] = 25'b1111111110111000100000110;
    rom[12503] = 25'b1111111110111000100001001;
    rom[12504] = 25'b1111111110111000100001100;
    rom[12505] = 25'b1111111110111000100001111;
    rom[12506] = 25'b1111111110111000100010011;
    rom[12507] = 25'b1111111110111000100010111;
    rom[12508] = 25'b1111111110111000100011011;
    rom[12509] = 25'b1111111110111000100011110;
    rom[12510] = 25'b1111111110111000100100010;
    rom[12511] = 25'b1111111110111000100100110;
    rom[12512] = 25'b1111111110111000100101010;
    rom[12513] = 25'b1111111110111000100101101;
    rom[12514] = 25'b1111111110111000100110010;
    rom[12515] = 25'b1111111110111000100110110;
    rom[12516] = 25'b1111111110111000100111010;
    rom[12517] = 25'b1111111110111000100111110;
    rom[12518] = 25'b1111111110111000101000010;
    rom[12519] = 25'b1111111110111000101000110;
    rom[12520] = 25'b1111111110111000101001010;
    rom[12521] = 25'b1111111110111000101001111;
    rom[12522] = 25'b1111111110111000101010011;
    rom[12523] = 25'b1111111110111000101011000;
    rom[12524] = 25'b1111111110111000101011100;
    rom[12525] = 25'b1111111110111000101100001;
    rom[12526] = 25'b1111111110111000101100101;
    rom[12527] = 25'b1111111110111000101101011;
    rom[12528] = 25'b1111111110111000101101111;
    rom[12529] = 25'b1111111110111000101110100;
    rom[12530] = 25'b1111111110111000101111001;
    rom[12531] = 25'b1111111110111000101111101;
    rom[12532] = 25'b1111111110111000110000011;
    rom[12533] = 25'b1111111110111000110001000;
    rom[12534] = 25'b1111111110111000110001101;
    rom[12535] = 25'b1111111110111000110010001;
    rom[12536] = 25'b1111111110111000110010111;
    rom[12537] = 25'b1111111110111000110011100;
    rom[12538] = 25'b1111111110111000110100001;
    rom[12539] = 25'b1111111110111000110100111;
    rom[12540] = 25'b1111111110111000110101100;
    rom[12541] = 25'b1111111110111000110110010;
    rom[12542] = 25'b1111111110111000110110111;
    rom[12543] = 25'b1111111110111000110111101;
    rom[12544] = 25'b1111111110111000111000010;
    rom[12545] = 25'b1111111110111000111001000;
    rom[12546] = 25'b1111111110111000111001110;
    rom[12547] = 25'b1111111110111000111010011;
    rom[12548] = 25'b1111111110111000111011001;
    rom[12549] = 25'b1111111110111000111011111;
    rom[12550] = 25'b1111111110111000111100101;
    rom[12551] = 25'b1111111110111000111101011;
    rom[12552] = 25'b1111111110111000111110001;
    rom[12553] = 25'b1111111110111000111110111;
    rom[12554] = 25'b1111111110111000111111110;
    rom[12555] = 25'b1111111110111001000000100;
    rom[12556] = 25'b1111111110111001000001010;
    rom[12557] = 25'b1111111110111001000010000;
    rom[12558] = 25'b1111111110111001000010111;
    rom[12559] = 25'b1111111110111001000011101;
    rom[12560] = 25'b1111111110111001000100100;
    rom[12561] = 25'b1111111110111001000101011;
    rom[12562] = 25'b1111111110111001000110001;
    rom[12563] = 25'b1111111110111001000110111;
    rom[12564] = 25'b1111111110111001000111110;
    rom[12565] = 25'b1111111110111001001000110;
    rom[12566] = 25'b1111111110111001001001100;
    rom[12567] = 25'b1111111110111001001010011;
    rom[12568] = 25'b1111111110111001001011010;
    rom[12569] = 25'b1111111110111001001100001;
    rom[12570] = 25'b1111111110111001001101000;
    rom[12571] = 25'b1111111110111001001101111;
    rom[12572] = 25'b1111111110111001001110110;
    rom[12573] = 25'b1111111110111001001111110;
    rom[12574] = 25'b1111111110111001010000101;
    rom[12575] = 25'b1111111110111001010001100;
    rom[12576] = 25'b1111111110111001010010011;
    rom[12577] = 25'b1111111110111001010011011;
    rom[12578] = 25'b1111111110111001010100010;
    rom[12579] = 25'b1111111110111001010101010;
    rom[12580] = 25'b1111111110111001010110010;
    rom[12581] = 25'b1111111110111001010111001;
    rom[12582] = 25'b1111111110111001011000001;
    rom[12583] = 25'b1111111110111001011001001;
    rom[12584] = 25'b1111111110111001011010000;
    rom[12585] = 25'b1111111110111001011011001;
    rom[12586] = 25'b1111111110111001011100000;
    rom[12587] = 25'b1111111110111001011101000;
    rom[12588] = 25'b1111111110111001011110001;
    rom[12589] = 25'b1111111110111001011111001;
    rom[12590] = 25'b1111111110111001100000001;
    rom[12591] = 25'b1111111110111001100001001;
    rom[12592] = 25'b1111111110111001100010001;
    rom[12593] = 25'b1111111110111001100011010;
    rom[12594] = 25'b1111111110111001100100010;
    rom[12595] = 25'b1111111110111001100101011;
    rom[12596] = 25'b1111111110111001100110011;
    rom[12597] = 25'b1111111110111001100111100;
    rom[12598] = 25'b1111111110111001101000100;
    rom[12599] = 25'b1111111110111001101001101;
    rom[12600] = 25'b1111111110111001101010110;
    rom[12601] = 25'b1111111110111001101011110;
    rom[12602] = 25'b1111111110111001101100111;
    rom[12603] = 25'b1111111110111001101110000;
    rom[12604] = 25'b1111111110111001101111001;
    rom[12605] = 25'b1111111110111001110000010;
    rom[12606] = 25'b1111111110111001110001011;
    rom[12607] = 25'b1111111110111001110010101;
    rom[12608] = 25'b1111111110111001110011110;
    rom[12609] = 25'b1111111110111001110100111;
    rom[12610] = 25'b1111111110111001110110001;
    rom[12611] = 25'b1111111110111001110111010;
    rom[12612] = 25'b1111111110111001111000011;
    rom[12613] = 25'b1111111110111001111001101;
    rom[12614] = 25'b1111111110111001111010110;
    rom[12615] = 25'b1111111110111001111100000;
    rom[12616] = 25'b1111111110111001111101001;
    rom[12617] = 25'b1111111110111001111110011;
    rom[12618] = 25'b1111111110111001111111101;
    rom[12619] = 25'b1111111110111010000000111;
    rom[12620] = 25'b1111111110111010000010001;
    rom[12621] = 25'b1111111110111010000011011;
    rom[12622] = 25'b1111111110111010000100100;
    rom[12623] = 25'b1111111110111010000101111;
    rom[12624] = 25'b1111111110111010000111001;
    rom[12625] = 25'b1111111110111010001000011;
    rom[12626] = 25'b1111111110111010001001110;
    rom[12627] = 25'b1111111110111010001010111;
    rom[12628] = 25'b1111111110111010001100010;
    rom[12629] = 25'b1111111110111010001101100;
    rom[12630] = 25'b1111111110111010001110111;
    rom[12631] = 25'b1111111110111010010000001;
    rom[12632] = 25'b1111111110111010010001100;
    rom[12633] = 25'b1111111110111010010010111;
    rom[12634] = 25'b1111111110111010010100001;
    rom[12635] = 25'b1111111110111010010101100;
    rom[12636] = 25'b1111111110111010010110111;
    rom[12637] = 25'b1111111110111010011000001;
    rom[12638] = 25'b1111111110111010011001101;
    rom[12639] = 25'b1111111110111010011010111;
    rom[12640] = 25'b1111111110111010011100010;
    rom[12641] = 25'b1111111110111010011101101;
    rom[12642] = 25'b1111111110111010011111001;
    rom[12643] = 25'b1111111110111010100000100;
    rom[12644] = 25'b1111111110111010100001111;
    rom[12645] = 25'b1111111110111010100011010;
    rom[12646] = 25'b1111111110111010100100101;
    rom[12647] = 25'b1111111110111010100110001;
    rom[12648] = 25'b1111111110111010100111101;
    rom[12649] = 25'b1111111110111010101001000;
    rom[12650] = 25'b1111111110111010101010100;
    rom[12651] = 25'b1111111110111010101100000;
    rom[12652] = 25'b1111111110111010101101011;
    rom[12653] = 25'b1111111110111010101110111;
    rom[12654] = 25'b1111111110111010110000011;
    rom[12655] = 25'b1111111110111010110001111;
    rom[12656] = 25'b1111111110111010110011011;
    rom[12657] = 25'b1111111110111010110100111;
    rom[12658] = 25'b1111111110111010110110011;
    rom[12659] = 25'b1111111110111010110111111;
    rom[12660] = 25'b1111111110111010111001011;
    rom[12661] = 25'b1111111110111010111010111;
    rom[12662] = 25'b1111111110111010111100011;
    rom[12663] = 25'b1111111110111010111110000;
    rom[12664] = 25'b1111111110111010111111100;
    rom[12665] = 25'b1111111110111011000001001;
    rom[12666] = 25'b1111111110111011000010101;
    rom[12667] = 25'b1111111110111011000100010;
    rom[12668] = 25'b1111111110111011000101111;
    rom[12669] = 25'b1111111110111011000111011;
    rom[12670] = 25'b1111111110111011001001000;
    rom[12671] = 25'b1111111110111011001010101;
    rom[12672] = 25'b1111111110111011001100001;
    rom[12673] = 25'b1111111110111011001101110;
    rom[12674] = 25'b1111111110111011001111100;
    rom[12675] = 25'b1111111110111011010001000;
    rom[12676] = 25'b1111111110111011010010110;
    rom[12677] = 25'b1111111110111011010100010;
    rom[12678] = 25'b1111111110111011010110000;
    rom[12679] = 25'b1111111110111011010111101;
    rom[12680] = 25'b1111111110111011011001011;
    rom[12681] = 25'b1111111110111011011010111;
    rom[12682] = 25'b1111111110111011011100101;
    rom[12683] = 25'b1111111110111011011110011;
    rom[12684] = 25'b1111111110111011100000001;
    rom[12685] = 25'b1111111110111011100001110;
    rom[12686] = 25'b1111111110111011100011011;
    rom[12687] = 25'b1111111110111011100101010;
    rom[12688] = 25'b1111111110111011100110111;
    rom[12689] = 25'b1111111110111011101000101;
    rom[12690] = 25'b1111111110111011101010011;
    rom[12691] = 25'b1111111110111011101100001;
    rom[12692] = 25'b1111111110111011101101111;
    rom[12693] = 25'b1111111110111011101111101;
    rom[12694] = 25'b1111111110111011110001100;
    rom[12695] = 25'b1111111110111011110011010;
    rom[12696] = 25'b1111111110111011110101000;
    rom[12697] = 25'b1111111110111011110110110;
    rom[12698] = 25'b1111111110111011111000100;
    rom[12699] = 25'b1111111110111011111010010;
    rom[12700] = 25'b1111111110111011111100001;
    rom[12701] = 25'b1111111110111011111110000;
    rom[12702] = 25'b1111111110111011111111111;
    rom[12703] = 25'b1111111110111100000001101;
    rom[12704] = 25'b1111111110111100000011100;
    rom[12705] = 25'b1111111110111100000101011;
    rom[12706] = 25'b1111111110111100000111010;
    rom[12707] = 25'b1111111110111100001001001;
    rom[12708] = 25'b1111111110111100001010111;
    rom[12709] = 25'b1111111110111100001100110;
    rom[12710] = 25'b1111111110111100001110101;
    rom[12711] = 25'b1111111110111100010000100;
    rom[12712] = 25'b1111111110111100010010100;
    rom[12713] = 25'b1111111110111100010100011;
    rom[12714] = 25'b1111111110111100010110011;
    rom[12715] = 25'b1111111110111100011000010;
    rom[12716] = 25'b1111111110111100011010001;
    rom[12717] = 25'b1111111110111100011100001;
    rom[12718] = 25'b1111111110111100011110000;
    rom[12719] = 25'b1111111110111100100000000;
    rom[12720] = 25'b1111111110111100100001111;
    rom[12721] = 25'b1111111110111100100011111;
    rom[12722] = 25'b1111111110111100100101111;
    rom[12723] = 25'b1111111110111100100111111;
    rom[12724] = 25'b1111111110111100101001111;
    rom[12725] = 25'b1111111110111100101011110;
    rom[12726] = 25'b1111111110111100101101111;
    rom[12727] = 25'b1111111110111100101111111;
    rom[12728] = 25'b1111111110111100110001111;
    rom[12729] = 25'b1111111110111100110011111;
    rom[12730] = 25'b1111111110111100110101111;
    rom[12731] = 25'b1111111110111100111000000;
    rom[12732] = 25'b1111111110111100111010000;
    rom[12733] = 25'b1111111110111100111100000;
    rom[12734] = 25'b1111111110111100111110001;
    rom[12735] = 25'b1111111110111101000000001;
    rom[12736] = 25'b1111111110111101000010010;
    rom[12737] = 25'b1111111110111101000100011;
    rom[12738] = 25'b1111111110111101000110011;
    rom[12739] = 25'b1111111110111101001000100;
    rom[12740] = 25'b1111111110111101001010101;
    rom[12741] = 25'b1111111110111101001100110;
    rom[12742] = 25'b1111111110111101001110111;
    rom[12743] = 25'b1111111110111101010001000;
    rom[12744] = 25'b1111111110111101010011001;
    rom[12745] = 25'b1111111110111101010101010;
    rom[12746] = 25'b1111111110111101010111011;
    rom[12747] = 25'b1111111110111101011001101;
    rom[12748] = 25'b1111111110111101011011110;
    rom[12749] = 25'b1111111110111101011101111;
    rom[12750] = 25'b1111111110111101100000001;
    rom[12751] = 25'b1111111110111101100010010;
    rom[12752] = 25'b1111111110111101100100100;
    rom[12753] = 25'b1111111110111101100110101;
    rom[12754] = 25'b1111111110111101101000111;
    rom[12755] = 25'b1111111110111101101011001;
    rom[12756] = 25'b1111111110111101101101010;
    rom[12757] = 25'b1111111110111101101111100;
    rom[12758] = 25'b1111111110111101110001110;
    rom[12759] = 25'b1111111110111101110100000;
    rom[12760] = 25'b1111111110111101110110010;
    rom[12761] = 25'b1111111110111101111000101;
    rom[12762] = 25'b1111111110111101111010111;
    rom[12763] = 25'b1111111110111101111101000;
    rom[12764] = 25'b1111111110111101111111011;
    rom[12765] = 25'b1111111110111110000001101;
    rom[12766] = 25'b1111111110111110000100000;
    rom[12767] = 25'b1111111110111110000110010;
    rom[12768] = 25'b1111111110111110001000100;
    rom[12769] = 25'b1111111110111110001010111;
    rom[12770] = 25'b1111111110111110001101010;
    rom[12771] = 25'b1111111110111110001111100;
    rom[12772] = 25'b1111111110111110010001111;
    rom[12773] = 25'b1111111110111110010100010;
    rom[12774] = 25'b1111111110111110010110100;
    rom[12775] = 25'b1111111110111110011001000;
    rom[12776] = 25'b1111111110111110011011010;
    rom[12777] = 25'b1111111110111110011101101;
    rom[12778] = 25'b1111111110111110100000001;
    rom[12779] = 25'b1111111110111110100010100;
    rom[12780] = 25'b1111111110111110100100111;
    rom[12781] = 25'b1111111110111110100111010;
    rom[12782] = 25'b1111111110111110101001110;
    rom[12783] = 25'b1111111110111110101100001;
    rom[12784] = 25'b1111111110111110101110100;
    rom[12785] = 25'b1111111110111110110001000;
    rom[12786] = 25'b1111111110111110110011011;
    rom[12787] = 25'b1111111110111110110101111;
    rom[12788] = 25'b1111111110111110111000011;
    rom[12789] = 25'b1111111110111110111010110;
    rom[12790] = 25'b1111111110111110111101010;
    rom[12791] = 25'b1111111110111110111111110;
    rom[12792] = 25'b1111111110111111000010010;
    rom[12793] = 25'b1111111110111111000100110;
    rom[12794] = 25'b1111111110111111000111010;
    rom[12795] = 25'b1111111110111111001001110;
    rom[12796] = 25'b1111111110111111001100010;
    rom[12797] = 25'b1111111110111111001110110;
    rom[12798] = 25'b1111111110111111010001010;
    rom[12799] = 25'b1111111110111111010011111;
    rom[12800] = 25'b1111111110111111010110011;
    rom[12801] = 25'b1111111110111111011001000;
    rom[12802] = 25'b1111111110111111011011100;
    rom[12803] = 25'b1111111110111111011110001;
    rom[12804] = 25'b1111111110111111100000110;
    rom[12805] = 25'b1111111110111111100011011;
    rom[12806] = 25'b1111111110111111100101111;
    rom[12807] = 25'b1111111110111111101000100;
    rom[12808] = 25'b1111111110111111101011001;
    rom[12809] = 25'b1111111110111111101101101;
    rom[12810] = 25'b1111111110111111110000010;
    rom[12811] = 25'b1111111110111111110010111;
    rom[12812] = 25'b1111111110111111110101101;
    rom[12813] = 25'b1111111110111111111000010;
    rom[12814] = 25'b1111111110111111111010111;
    rom[12815] = 25'b1111111110111111111101100;
    rom[12816] = 25'b1111111111000000000000001;
    rom[12817] = 25'b1111111111000000000010111;
    rom[12818] = 25'b1111111111000000000101101;
    rom[12819] = 25'b1111111111000000001000010;
    rom[12820] = 25'b1111111111000000001010111;
    rom[12821] = 25'b1111111111000000001101101;
    rom[12822] = 25'b1111111111000000010000011;
    rom[12823] = 25'b1111111111000000010011001;
    rom[12824] = 25'b1111111111000000010101111;
    rom[12825] = 25'b1111111111000000011000100;
    rom[12826] = 25'b1111111111000000011011010;
    rom[12827] = 25'b1111111111000000011110000;
    rom[12828] = 25'b1111111111000000100000110;
    rom[12829] = 25'b1111111111000000100011101;
    rom[12830] = 25'b1111111111000000100110011;
    rom[12831] = 25'b1111111111000000101001001;
    rom[12832] = 25'b1111111111000000101011111;
    rom[12833] = 25'b1111111111000000101110101;
    rom[12834] = 25'b1111111111000000110001100;
    rom[12835] = 25'b1111111111000000110100010;
    rom[12836] = 25'b1111111111000000110111001;
    rom[12837] = 25'b1111111111000000111010000;
    rom[12838] = 25'b1111111111000000111100110;
    rom[12839] = 25'b1111111111000000111111101;
    rom[12840] = 25'b1111111111000001000010100;
    rom[12841] = 25'b1111111111000001000101010;
    rom[12842] = 25'b1111111111000001001000001;
    rom[12843] = 25'b1111111111000001001011001;
    rom[12844] = 25'b1111111111000001001110000;
    rom[12845] = 25'b1111111111000001010000110;
    rom[12846] = 25'b1111111111000001010011101;
    rom[12847] = 25'b1111111111000001010110100;
    rom[12848] = 25'b1111111111000001011001100;
    rom[12849] = 25'b1111111111000001011100011;
    rom[12850] = 25'b1111111111000001011111011;
    rom[12851] = 25'b1111111111000001100010010;
    rom[12852] = 25'b1111111111000001100101010;
    rom[12853] = 25'b1111111111000001101000001;
    rom[12854] = 25'b1111111111000001101011001;
    rom[12855] = 25'b1111111111000001101110001;
    rom[12856] = 25'b1111111111000001110001000;
    rom[12857] = 25'b1111111111000001110100000;
    rom[12858] = 25'b1111111111000001110111000;
    rom[12859] = 25'b1111111111000001111010000;
    rom[12860] = 25'b1111111111000001111100111;
    rom[12861] = 25'b1111111111000001111111111;
    rom[12862] = 25'b1111111111000010000010111;
    rom[12863] = 25'b1111111111000010000110000;
    rom[12864] = 25'b1111111111000010001001000;
    rom[12865] = 25'b1111111111000010001100001;
    rom[12866] = 25'b1111111111000010001111000;
    rom[12867] = 25'b1111111111000010010010001;
    rom[12868] = 25'b1111111111000010010101010;
    rom[12869] = 25'b1111111111000010011000010;
    rom[12870] = 25'b1111111111000010011011010;
    rom[12871] = 25'b1111111111000010011110011;
    rom[12872] = 25'b1111111111000010100001100;
    rom[12873] = 25'b1111111111000010100100100;
    rom[12874] = 25'b1111111111000010100111110;
    rom[12875] = 25'b1111111111000010101010110;
    rom[12876] = 25'b1111111111000010101101111;
    rom[12877] = 25'b1111111111000010110001000;
    rom[12878] = 25'b1111111111000010110100001;
    rom[12879] = 25'b1111111111000010110111010;
    rom[12880] = 25'b1111111111000010111010011;
    rom[12881] = 25'b1111111111000010111101100;
    rom[12882] = 25'b1111111111000011000000110;
    rom[12883] = 25'b1111111111000011000011111;
    rom[12884] = 25'b1111111111000011000111001;
    rom[12885] = 25'b1111111111000011001010010;
    rom[12886] = 25'b1111111111000011001101011;
    rom[12887] = 25'b1111111111000011010000101;
    rom[12888] = 25'b1111111111000011010011111;
    rom[12889] = 25'b1111111111000011010111000;
    rom[12890] = 25'b1111111111000011011010010;
    rom[12891] = 25'b1111111111000011011101100;
    rom[12892] = 25'b1111111111000011100000110;
    rom[12893] = 25'b1111111111000011100100000;
    rom[12894] = 25'b1111111111000011100111010;
    rom[12895] = 25'b1111111111000011101010100;
    rom[12896] = 25'b1111111111000011101101110;
    rom[12897] = 25'b1111111111000011110001000;
    rom[12898] = 25'b1111111111000011110100010;
    rom[12899] = 25'b1111111111000011110111100;
    rom[12900] = 25'b1111111111000011111010111;
    rom[12901] = 25'b1111111111000011111110001;
    rom[12902] = 25'b1111111111000100000001100;
    rom[12903] = 25'b1111111111000100000100111;
    rom[12904] = 25'b1111111111000100001000001;
    rom[12905] = 25'b1111111111000100001011100;
    rom[12906] = 25'b1111111111000100001110110;
    rom[12907] = 25'b1111111111000100010010001;
    rom[12908] = 25'b1111111111000100010101100;
    rom[12909] = 25'b1111111111000100011000111;
    rom[12910] = 25'b1111111111000100011100010;
    rom[12911] = 25'b1111111111000100011111101;
    rom[12912] = 25'b1111111111000100100011000;
    rom[12913] = 25'b1111111111000100100110011;
    rom[12914] = 25'b1111111111000100101001110;
    rom[12915] = 25'b1111111111000100101101001;
    rom[12916] = 25'b1111111111000100110000101;
    rom[12917] = 25'b1111111111000100110100000;
    rom[12918] = 25'b1111111111000100110111011;
    rom[12919] = 25'b1111111111000100111010111;
    rom[12920] = 25'b1111111111000100111110011;
    rom[12921] = 25'b1111111111000101000001110;
    rom[12922] = 25'b1111111111000101000101010;
    rom[12923] = 25'b1111111111000101001000110;
    rom[12924] = 25'b1111111111000101001100001;
    rom[12925] = 25'b1111111111000101001111101;
    rom[12926] = 25'b1111111111000101010011001;
    rom[12927] = 25'b1111111111000101010110101;
    rom[12928] = 25'b1111111111000101011010001;
    rom[12929] = 25'b1111111111000101011101101;
    rom[12930] = 25'b1111111111000101100001001;
    rom[12931] = 25'b1111111111000101100100101;
    rom[12932] = 25'b1111111111000101101000001;
    rom[12933] = 25'b1111111111000101101011110;
    rom[12934] = 25'b1111111111000101101111010;
    rom[12935] = 25'b1111111111000101110010111;
    rom[12936] = 25'b1111111111000101110110011;
    rom[12937] = 25'b1111111111000101111010000;
    rom[12938] = 25'b1111111111000101111101100;
    rom[12939] = 25'b1111111111000110000001001;
    rom[12940] = 25'b1111111111000110000100110;
    rom[12941] = 25'b1111111111000110001000010;
    rom[12942] = 25'b1111111111000110001100000;
    rom[12943] = 25'b1111111111000110001111101;
    rom[12944] = 25'b1111111111000110010011001;
    rom[12945] = 25'b1111111111000110010110110;
    rom[12946] = 25'b1111111111000110011010011;
    rom[12947] = 25'b1111111111000110011110000;
    rom[12948] = 25'b1111111111000110100001110;
    rom[12949] = 25'b1111111111000110100101100;
    rom[12950] = 25'b1111111111000110101001001;
    rom[12951] = 25'b1111111111000110101100110;
    rom[12952] = 25'b1111111111000110110000100;
    rom[12953] = 25'b1111111111000110110100001;
    rom[12954] = 25'b1111111111000110110111111;
    rom[12955] = 25'b1111111111000110111011100;
    rom[12956] = 25'b1111111111000110111111010;
    rom[12957] = 25'b1111111111000111000011000;
    rom[12958] = 25'b1111111111000111000110101;
    rom[12959] = 25'b1111111111000111001010011;
    rom[12960] = 25'b1111111111000111001110001;
    rom[12961] = 25'b1111111111000111010001111;
    rom[12962] = 25'b1111111111000111010101101;
    rom[12963] = 25'b1111111111000111011001011;
    rom[12964] = 25'b1111111111000111011101010;
    rom[12965] = 25'b1111111111000111100000111;
    rom[12966] = 25'b1111111111000111100100110;
    rom[12967] = 25'b1111111111000111101000100;
    rom[12968] = 25'b1111111111000111101100011;
    rom[12969] = 25'b1111111111000111110000001;
    rom[12970] = 25'b1111111111000111110100000;
    rom[12971] = 25'b1111111111000111110111110;
    rom[12972] = 25'b1111111111000111111011101;
    rom[12973] = 25'b1111111111000111111111100;
    rom[12974] = 25'b1111111111001000000011010;
    rom[12975] = 25'b1111111111001000000111001;
    rom[12976] = 25'b1111111111001000001011000;
    rom[12977] = 25'b1111111111001000001110111;
    rom[12978] = 25'b1111111111001000010010110;
    rom[12979] = 25'b1111111111001000010110101;
    rom[12980] = 25'b1111111111001000011010100;
    rom[12981] = 25'b1111111111001000011110011;
    rom[12982] = 25'b1111111111001000100010010;
    rom[12983] = 25'b1111111111001000100110010;
    rom[12984] = 25'b1111111111001000101010001;
    rom[12985] = 25'b1111111111001000101110001;
    rom[12986] = 25'b1111111111001000110010000;
    rom[12987] = 25'b1111111111001000110101111;
    rom[12988] = 25'b1111111111001000111001111;
    rom[12989] = 25'b1111111111001000111101111;
    rom[12990] = 25'b1111111111001001000001110;
    rom[12991] = 25'b1111111111001001000101110;
    rom[12992] = 25'b1111111111001001001001110;
    rom[12993] = 25'b1111111111001001001101110;
    rom[12994] = 25'b1111111111001001010001110;
    rom[12995] = 25'b1111111111001001010101110;
    rom[12996] = 25'b1111111111001001011001110;
    rom[12997] = 25'b1111111111001001011101110;
    rom[12998] = 25'b1111111111001001100001110;
    rom[12999] = 25'b1111111111001001100101111;
    rom[13000] = 25'b1111111111001001101001111;
    rom[13001] = 25'b1111111111001001101101111;
    rom[13002] = 25'b1111111111001001110010000;
    rom[13003] = 25'b1111111111001001110110000;
    rom[13004] = 25'b1111111111001001111010001;
    rom[13005] = 25'b1111111111001001111110001;
    rom[13006] = 25'b1111111111001010000010010;
    rom[13007] = 25'b1111111111001010000110011;
    rom[13008] = 25'b1111111111001010001010011;
    rom[13009] = 25'b1111111111001010001110100;
    rom[13010] = 25'b1111111111001010010010101;
    rom[13011] = 25'b1111111111001010010110110;
    rom[13012] = 25'b1111111111001010011010111;
    rom[13013] = 25'b1111111111001010011111000;
    rom[13014] = 25'b1111111111001010100011001;
    rom[13015] = 25'b1111111111001010100111010;
    rom[13016] = 25'b1111111111001010101011011;
    rom[13017] = 25'b1111111111001010101111101;
    rom[13018] = 25'b1111111111001010110011110;
    rom[13019] = 25'b1111111111001010110111111;
    rom[13020] = 25'b1111111111001010111100001;
    rom[13021] = 25'b1111111111001011000000010;
    rom[13022] = 25'b1111111111001011000100100;
    rom[13023] = 25'b1111111111001011001000110;
    rom[13024] = 25'b1111111111001011001100111;
    rom[13025] = 25'b1111111111001011010001001;
    rom[13026] = 25'b1111111111001011010101011;
    rom[13027] = 25'b1111111111001011011001101;
    rom[13028] = 25'b1111111111001011011101111;
    rom[13029] = 25'b1111111111001011100010001;
    rom[13030] = 25'b1111111111001011100110011;
    rom[13031] = 25'b1111111111001011101010101;
    rom[13032] = 25'b1111111111001011101110111;
    rom[13033] = 25'b1111111111001011110011010;
    rom[13034] = 25'b1111111111001011110111100;
    rom[13035] = 25'b1111111111001011111011110;
    rom[13036] = 25'b1111111111001100000000001;
    rom[13037] = 25'b1111111111001100000100011;
    rom[13038] = 25'b1111111111001100001000101;
    rom[13039] = 25'b1111111111001100001101000;
    rom[13040] = 25'b1111111111001100010001011;
    rom[13041] = 25'b1111111111001100010101101;
    rom[13042] = 25'b1111111111001100011010000;
    rom[13043] = 25'b1111111111001100011110011;
    rom[13044] = 25'b1111111111001100100010110;
    rom[13045] = 25'b1111111111001100100111001;
    rom[13046] = 25'b1111111111001100101011100;
    rom[13047] = 25'b1111111111001100101111110;
    rom[13048] = 25'b1111111111001100110100010;
    rom[13049] = 25'b1111111111001100111000101;
    rom[13050] = 25'b1111111111001100111101001;
    rom[13051] = 25'b1111111111001101000001100;
    rom[13052] = 25'b1111111111001101000101111;
    rom[13053] = 25'b1111111111001101001010011;
    rom[13054] = 25'b1111111111001101001110110;
    rom[13055] = 25'b1111111111001101010011010;
    rom[13056] = 25'b1111111111001101010111101;
    rom[13057] = 25'b1111111111001101011100001;
    rom[13058] = 25'b1111111111001101100000100;
    rom[13059] = 25'b1111111111001101100101000;
    rom[13060] = 25'b1111111111001101101001100;
    rom[13061] = 25'b1111111111001101101110000;
    rom[13062] = 25'b1111111111001101110010100;
    rom[13063] = 25'b1111111111001101110111000;
    rom[13064] = 25'b1111111111001101111011100;
    rom[13065] = 25'b1111111111001110000000000;
    rom[13066] = 25'b1111111111001110000100100;
    rom[13067] = 25'b1111111111001110001001000;
    rom[13068] = 25'b1111111111001110001101101;
    rom[13069] = 25'b1111111111001110010010001;
    rom[13070] = 25'b1111111111001110010110101;
    rom[13071] = 25'b1111111111001110011011010;
    rom[13072] = 25'b1111111111001110011111110;
    rom[13073] = 25'b1111111111001110100100011;
    rom[13074] = 25'b1111111111001110101000111;
    rom[13075] = 25'b1111111111001110101101100;
    rom[13076] = 25'b1111111111001110110010001;
    rom[13077] = 25'b1111111111001110110110101;
    rom[13078] = 25'b1111111111001110111011011;
    rom[13079] = 25'b1111111111001110111111111;
    rom[13080] = 25'b1111111111001111000100101;
    rom[13081] = 25'b1111111111001111001001001;
    rom[13082] = 25'b1111111111001111001101111;
    rom[13083] = 25'b1111111111001111010010100;
    rom[13084] = 25'b1111111111001111010111001;
    rom[13085] = 25'b1111111111001111011011110;
    rom[13086] = 25'b1111111111001111100000011;
    rom[13087] = 25'b1111111111001111100101001;
    rom[13088] = 25'b1111111111001111101001110;
    rom[13089] = 25'b1111111111001111101110100;
    rom[13090] = 25'b1111111111001111110011001;
    rom[13091] = 25'b1111111111001111110111111;
    rom[13092] = 25'b1111111111001111111100101;
    rom[13093] = 25'b1111111111010000000001010;
    rom[13094] = 25'b1111111111010000000110000;
    rom[13095] = 25'b1111111111010000001010110;
    rom[13096] = 25'b1111111111010000001111100;
    rom[13097] = 25'b1111111111010000010100010;
    rom[13098] = 25'b1111111111010000011001000;
    rom[13099] = 25'b1111111111010000011101110;
    rom[13100] = 25'b1111111111010000100010100;
    rom[13101] = 25'b1111111111010000100111010;
    rom[13102] = 25'b1111111111010000101100000;
    rom[13103] = 25'b1111111111010000110000111;
    rom[13104] = 25'b1111111111010000110101101;
    rom[13105] = 25'b1111111111010000111010011;
    rom[13106] = 25'b1111111111010000111111010;
    rom[13107] = 25'b1111111111010001000100000;
    rom[13108] = 25'b1111111111010001001000111;
    rom[13109] = 25'b1111111111010001001101110;
    rom[13110] = 25'b1111111111010001010010101;
    rom[13111] = 25'b1111111111010001010111011;
    rom[13112] = 25'b1111111111010001011100010;
    rom[13113] = 25'b1111111111010001100001001;
    rom[13114] = 25'b1111111111010001100110000;
    rom[13115] = 25'b1111111111010001101010111;
    rom[13116] = 25'b1111111111010001101111110;
    rom[13117] = 25'b1111111111010001110100101;
    rom[13118] = 25'b1111111111010001111001100;
    rom[13119] = 25'b1111111111010001111110011;
    rom[13120] = 25'b1111111111010010000011011;
    rom[13121] = 25'b1111111111010010001000010;
    rom[13122] = 25'b1111111111010010001101001;
    rom[13123] = 25'b1111111111010010010010001;
    rom[13124] = 25'b1111111111010010010111001;
    rom[13125] = 25'b1111111111010010011100000;
    rom[13126] = 25'b1111111111010010100001000;
    rom[13127] = 25'b1111111111010010100101111;
    rom[13128] = 25'b1111111111010010101010111;
    rom[13129] = 25'b1111111111010010101111111;
    rom[13130] = 25'b1111111111010010110100111;
    rom[13131] = 25'b1111111111010010111001110;
    rom[13132] = 25'b1111111111010010111110111;
    rom[13133] = 25'b1111111111010011000011110;
    rom[13134] = 25'b1111111111010011001000111;
    rom[13135] = 25'b1111111111010011001101111;
    rom[13136] = 25'b1111111111010011010010111;
    rom[13137] = 25'b1111111111010011010111111;
    rom[13138] = 25'b1111111111010011011100111;
    rom[13139] = 25'b1111111111010011100010000;
    rom[13140] = 25'b1111111111010011100111000;
    rom[13141] = 25'b1111111111010011101100000;
    rom[13142] = 25'b1111111111010011110001010;
    rom[13143] = 25'b1111111111010011110110010;
    rom[13144] = 25'b1111111111010011111011010;
    rom[13145] = 25'b1111111111010100000000011;
    rom[13146] = 25'b1111111111010100000101100;
    rom[13147] = 25'b1111111111010100001010101;
    rom[13148] = 25'b1111111111010100001111110;
    rom[13149] = 25'b1111111111010100010100111;
    rom[13150] = 25'b1111111111010100011001111;
    rom[13151] = 25'b1111111111010100011111000;
    rom[13152] = 25'b1111111111010100100100001;
    rom[13153] = 25'b1111111111010100101001011;
    rom[13154] = 25'b1111111111010100101110100;
    rom[13155] = 25'b1111111111010100110011101;
    rom[13156] = 25'b1111111111010100111000111;
    rom[13157] = 25'b1111111111010100111110000;
    rom[13158] = 25'b1111111111010101000011001;
    rom[13159] = 25'b1111111111010101001000011;
    rom[13160] = 25'b1111111111010101001101100;
    rom[13161] = 25'b1111111111010101010010110;
    rom[13162] = 25'b1111111111010101011000000;
    rom[13163] = 25'b1111111111010101011101001;
    rom[13164] = 25'b1111111111010101100010011;
    rom[13165] = 25'b1111111111010101100111101;
    rom[13166] = 25'b1111111111010101101100111;
    rom[13167] = 25'b1111111111010101110010001;
    rom[13168] = 25'b1111111111010101110111011;
    rom[13169] = 25'b1111111111010101111100101;
    rom[13170] = 25'b1111111111010110000001111;
    rom[13171] = 25'b1111111111010110000111001;
    rom[13172] = 25'b1111111111010110001100011;
    rom[13173] = 25'b1111111111010110010001110;
    rom[13174] = 25'b1111111111010110010111000;
    rom[13175] = 25'b1111111111010110011100010;
    rom[13176] = 25'b1111111111010110100001101;
    rom[13177] = 25'b1111111111010110100110111;
    rom[13178] = 25'b1111111111010110101100010;
    rom[13179] = 25'b1111111111010110110001101;
    rom[13180] = 25'b1111111111010110110110111;
    rom[13181] = 25'b1111111111010110111100010;
    rom[13182] = 25'b1111111111010111000001100;
    rom[13183] = 25'b1111111111010111000111000;
    rom[13184] = 25'b1111111111010111001100010;
    rom[13185] = 25'b1111111111010111010001110;
    rom[13186] = 25'b1111111111010111010111000;
    rom[13187] = 25'b1111111111010111011100011;
    rom[13188] = 25'b1111111111010111100001111;
    rom[13189] = 25'b1111111111010111100111001;
    rom[13190] = 25'b1111111111010111101100101;
    rom[13191] = 25'b1111111111010111110010000;
    rom[13192] = 25'b1111111111010111110111011;
    rom[13193] = 25'b1111111111010111111100111;
    rom[13194] = 25'b1111111111011000000010010;
    rom[13195] = 25'b1111111111011000000111110;
    rom[13196] = 25'b1111111111011000001101001;
    rom[13197] = 25'b1111111111011000010010101;
    rom[13198] = 25'b1111111111011000011000001;
    rom[13199] = 25'b1111111111011000011101100;
    rom[13200] = 25'b1111111111011000100011000;
    rom[13201] = 25'b1111111111011000101000100;
    rom[13202] = 25'b1111111111011000101110000;
    rom[13203] = 25'b1111111111011000110011100;
    rom[13204] = 25'b1111111111011000111001000;
    rom[13205] = 25'b1111111111011000111110100;
    rom[13206] = 25'b1111111111011001000100000;
    rom[13207] = 25'b1111111111011001001001100;
    rom[13208] = 25'b1111111111011001001111000;
    rom[13209] = 25'b1111111111011001010100100;
    rom[13210] = 25'b1111111111011001011010001;
    rom[13211] = 25'b1111111111011001011111101;
    rom[13212] = 25'b1111111111011001100101001;
    rom[13213] = 25'b1111111111011001101010110;
    rom[13214] = 25'b1111111111011001110000011;
    rom[13215] = 25'b1111111111011001110101111;
    rom[13216] = 25'b1111111111011001111011100;
    rom[13217] = 25'b1111111111011010000001001;
    rom[13218] = 25'b1111111111011010000110101;
    rom[13219] = 25'b1111111111011010001100010;
    rom[13220] = 25'b1111111111011010010001111;
    rom[13221] = 25'b1111111111011010010111100;
    rom[13222] = 25'b1111111111011010011101001;
    rom[13223] = 25'b1111111111011010100010110;
    rom[13224] = 25'b1111111111011010101000011;
    rom[13225] = 25'b1111111111011010101110000;
    rom[13226] = 25'b1111111111011010110011110;
    rom[13227] = 25'b1111111111011010111001010;
    rom[13228] = 25'b1111111111011010111111000;
    rom[13229] = 25'b1111111111011011000100101;
    rom[13230] = 25'b1111111111011011001010010;
    rom[13231] = 25'b1111111111011011010000000;
    rom[13232] = 25'b1111111111011011010101101;
    rom[13233] = 25'b1111111111011011011011011;
    rom[13234] = 25'b1111111111011011100001001;
    rom[13235] = 25'b1111111111011011100110110;
    rom[13236] = 25'b1111111111011011101100100;
    rom[13237] = 25'b1111111111011011110010010;
    rom[13238] = 25'b1111111111011011111000000;
    rom[13239] = 25'b1111111111011011111101110;
    rom[13240] = 25'b1111111111011100000011100;
    rom[13241] = 25'b1111111111011100001001010;
    rom[13242] = 25'b1111111111011100001110111;
    rom[13243] = 25'b1111111111011100010100110;
    rom[13244] = 25'b1111111111011100011010100;
    rom[13245] = 25'b1111111111011100100000010;
    rom[13246] = 25'b1111111111011100100110001;
    rom[13247] = 25'b1111111111011100101011111;
    rom[13248] = 25'b1111111111011100110001101;
    rom[13249] = 25'b1111111111011100110111100;
    rom[13250] = 25'b1111111111011100111101010;
    rom[13251] = 25'b1111111111011101000011000;
    rom[13252] = 25'b1111111111011101001000111;
    rom[13253] = 25'b1111111111011101001110110;
    rom[13254] = 25'b1111111111011101010100101;
    rom[13255] = 25'b1111111111011101011010011;
    rom[13256] = 25'b1111111111011101100000010;
    rom[13257] = 25'b1111111111011101100110001;
    rom[13258] = 25'b1111111111011101101100000;
    rom[13259] = 25'b1111111111011101110001111;
    rom[13260] = 25'b1111111111011101110111110;
    rom[13261] = 25'b1111111111011101111101101;
    rom[13262] = 25'b1111111111011110000011100;
    rom[13263] = 25'b1111111111011110001001011;
    rom[13264] = 25'b1111111111011110001111011;
    rom[13265] = 25'b1111111111011110010101010;
    rom[13266] = 25'b1111111111011110011011001;
    rom[13267] = 25'b1111111111011110100001001;
    rom[13268] = 25'b1111111111011110100111000;
    rom[13269] = 25'b1111111111011110101101000;
    rom[13270] = 25'b1111111111011110110010111;
    rom[13271] = 25'b1111111111011110111000110;
    rom[13272] = 25'b1111111111011110111110110;
    rom[13273] = 25'b1111111111011111000100110;
    rom[13274] = 25'b1111111111011111001010110;
    rom[13275] = 25'b1111111111011111010000110;
    rom[13276] = 25'b1111111111011111010110101;
    rom[13277] = 25'b1111111111011111011100101;
    rom[13278] = 25'b1111111111011111100010101;
    rom[13279] = 25'b1111111111011111101000101;
    rom[13280] = 25'b1111111111011111101110101;
    rom[13281] = 25'b1111111111011111110100101;
    rom[13282] = 25'b1111111111011111111010101;
    rom[13283] = 25'b1111111111100000000000110;
    rom[13284] = 25'b1111111111100000000110110;
    rom[13285] = 25'b1111111111100000001100110;
    rom[13286] = 25'b1111111111100000010010111;
    rom[13287] = 25'b1111111111100000011000111;
    rom[13288] = 25'b1111111111100000011111000;
    rom[13289] = 25'b1111111111100000100101000;
    rom[13290] = 25'b1111111111100000101011001;
    rom[13291] = 25'b1111111111100000110001001;
    rom[13292] = 25'b1111111111100000110111010;
    rom[13293] = 25'b1111111111100000111101011;
    rom[13294] = 25'b1111111111100001000011100;
    rom[13295] = 25'b1111111111100001001001100;
    rom[13296] = 25'b1111111111100001001111110;
    rom[13297] = 25'b1111111111100001010101110;
    rom[13298] = 25'b1111111111100001011100000;
    rom[13299] = 25'b1111111111100001100010000;
    rom[13300] = 25'b1111111111100001101000001;
    rom[13301] = 25'b1111111111100001101110011;
    rom[13302] = 25'b1111111111100001110100100;
    rom[13303] = 25'b1111111111100001111010101;
    rom[13304] = 25'b1111111111100010000000111;
    rom[13305] = 25'b1111111111100010000111000;
    rom[13306] = 25'b1111111111100010001101001;
    rom[13307] = 25'b1111111111100010010011011;
    rom[13308] = 25'b1111111111100010011001100;
    rom[13309] = 25'b1111111111100010011111110;
    rom[13310] = 25'b1111111111100010100101111;
    rom[13311] = 25'b1111111111100010101100001;
    rom[13312] = 25'b1111111111100010110010011;
    rom[13313] = 25'b1111111111100010111000101;
    rom[13314] = 25'b1111111111100010111110111;
    rom[13315] = 25'b1111111111100011000101000;
    rom[13316] = 25'b1111111111100011001011010;
    rom[13317] = 25'b1111111111100011010001100;
    rom[13318] = 25'b1111111111100011010111110;
    rom[13319] = 25'b1111111111100011011110000;
    rom[13320] = 25'b1111111111100011100100010;
    rom[13321] = 25'b1111111111100011101010100;
    rom[13322] = 25'b1111111111100011110000111;
    rom[13323] = 25'b1111111111100011110111001;
    rom[13324] = 25'b1111111111100011111101011;
    rom[13325] = 25'b1111111111100100000011110;
    rom[13326] = 25'b1111111111100100001010000;
    rom[13327] = 25'b1111111111100100010000011;
    rom[13328] = 25'b1111111111100100010110101;
    rom[13329] = 25'b1111111111100100011101000;
    rom[13330] = 25'b1111111111100100100011011;
    rom[13331] = 25'b1111111111100100101001101;
    rom[13332] = 25'b1111111111100100110000000;
    rom[13333] = 25'b1111111111100100110110011;
    rom[13334] = 25'b1111111111100100111100110;
    rom[13335] = 25'b1111111111100101000011001;
    rom[13336] = 25'b1111111111100101001001011;
    rom[13337] = 25'b1111111111100101001111110;
    rom[13338] = 25'b1111111111100101010110010;
    rom[13339] = 25'b1111111111100101011100101;
    rom[13340] = 25'b1111111111100101100010111;
    rom[13341] = 25'b1111111111100101101001011;
    rom[13342] = 25'b1111111111100101101111110;
    rom[13343] = 25'b1111111111100101110110001;
    rom[13344] = 25'b1111111111100101111100101;
    rom[13345] = 25'b1111111111100110000011000;
    rom[13346] = 25'b1111111111100110001001100;
    rom[13347] = 25'b1111111111100110001111111;
    rom[13348] = 25'b1111111111100110010110010;
    rom[13349] = 25'b1111111111100110011100110;
    rom[13350] = 25'b1111111111100110100011010;
    rom[13351] = 25'b1111111111100110101001110;
    rom[13352] = 25'b1111111111100110110000001;
    rom[13353] = 25'b1111111111100110110110101;
    rom[13354] = 25'b1111111111100110111101001;
    rom[13355] = 25'b1111111111100111000011101;
    rom[13356] = 25'b1111111111100111001010001;
    rom[13357] = 25'b1111111111100111010000100;
    rom[13358] = 25'b1111111111100111010111001;
    rom[13359] = 25'b1111111111100111011101101;
    rom[13360] = 25'b1111111111100111100100001;
    rom[13361] = 25'b1111111111100111101010101;
    rom[13362] = 25'b1111111111100111110001001;
    rom[13363] = 25'b1111111111100111110111110;
    rom[13364] = 25'b1111111111100111111110010;
    rom[13365] = 25'b1111111111101000000100110;
    rom[13366] = 25'b1111111111101000001011010;
    rom[13367] = 25'b1111111111101000010001111;
    rom[13368] = 25'b1111111111101000011000100;
    rom[13369] = 25'b1111111111101000011111000;
    rom[13370] = 25'b1111111111101000100101101;
    rom[13371] = 25'b1111111111101000101100001;
    rom[13372] = 25'b1111111111101000110010110;
    rom[13373] = 25'b1111111111101000111001011;
    rom[13374] = 25'b1111111111101001000000000;
    rom[13375] = 25'b1111111111101001000110101;
    rom[13376] = 25'b1111111111101001001101010;
    rom[13377] = 25'b1111111111101001010011111;
    rom[13378] = 25'b1111111111101001011010100;
    rom[13379] = 25'b1111111111101001100001001;
    rom[13380] = 25'b1111111111101001100111110;
    rom[13381] = 25'b1111111111101001101110011;
    rom[13382] = 25'b1111111111101001110101000;
    rom[13383] = 25'b1111111111101001111011101;
    rom[13384] = 25'b1111111111101010000010011;
    rom[13385] = 25'b1111111111101010001001000;
    rom[13386] = 25'b1111111111101010001111101;
    rom[13387] = 25'b1111111111101010010110011;
    rom[13388] = 25'b1111111111101010011101001;
    rom[13389] = 25'b1111111111101010100011110;
    rom[13390] = 25'b1111111111101010101010011;
    rom[13391] = 25'b1111111111101010110001001;
    rom[13392] = 25'b1111111111101010110111111;
    rom[13393] = 25'b1111111111101010111110100;
    rom[13394] = 25'b1111111111101011000101010;
    rom[13395] = 25'b1111111111101011001100000;
    rom[13396] = 25'b1111111111101011010010110;
    rom[13397] = 25'b1111111111101011011001100;
    rom[13398] = 25'b1111111111101011100000010;
    rom[13399] = 25'b1111111111101011100111000;
    rom[13400] = 25'b1111111111101011101101110;
    rom[13401] = 25'b1111111111101011110100100;
    rom[13402] = 25'b1111111111101011111011010;
    rom[13403] = 25'b1111111111101100000010000;
    rom[13404] = 25'b1111111111101100001000111;
    rom[13405] = 25'b1111111111101100001111101;
    rom[13406] = 25'b1111111111101100010110011;
    rom[13407] = 25'b1111111111101100011101010;
    rom[13408] = 25'b1111111111101100100100000;
    rom[13409] = 25'b1111111111101100101010111;
    rom[13410] = 25'b1111111111101100110001101;
    rom[13411] = 25'b1111111111101100111000100;
    rom[13412] = 25'b1111111111101100111111010;
    rom[13413] = 25'b1111111111101101000110001;
    rom[13414] = 25'b1111111111101101001100111;
    rom[13415] = 25'b1111111111101101010011110;
    rom[13416] = 25'b1111111111101101011010101;
    rom[13417] = 25'b1111111111101101100001100;
    rom[13418] = 25'b1111111111101101101000011;
    rom[13419] = 25'b1111111111101101101111010;
    rom[13420] = 25'b1111111111101101110110001;
    rom[13421] = 25'b1111111111101101111100111;
    rom[13422] = 25'b1111111111101110000011111;
    rom[13423] = 25'b1111111111101110001010110;
    rom[13424] = 25'b1111111111101110010001101;
    rom[13425] = 25'b1111111111101110011000101;
    rom[13426] = 25'b1111111111101110011111100;
    rom[13427] = 25'b1111111111101110100110011;
    rom[13428] = 25'b1111111111101110101101010;
    rom[13429] = 25'b1111111111101110110100010;
    rom[13430] = 25'b1111111111101110111011001;
    rom[13431] = 25'b1111111111101111000010000;
    rom[13432] = 25'b1111111111101111001001000;
    rom[13433] = 25'b1111111111101111010000000;
    rom[13434] = 25'b1111111111101111010111000;
    rom[13435] = 25'b1111111111101111011101111;
    rom[13436] = 25'b1111111111101111100100111;
    rom[13437] = 25'b1111111111101111101011110;
    rom[13438] = 25'b1111111111101111110010110;
    rom[13439] = 25'b1111111111101111111001110;
    rom[13440] = 25'b1111111111110000000000110;
    rom[13441] = 25'b1111111111110000000111110;
    rom[13442] = 25'b1111111111110000001110110;
    rom[13443] = 25'b1111111111110000010101110;
    rom[13444] = 25'b1111111111110000011100110;
    rom[13445] = 25'b1111111111110000100011110;
    rom[13446] = 25'b1111111111110000101010111;
    rom[13447] = 25'b1111111111110000110001111;
    rom[13448] = 25'b1111111111110000111000111;
    rom[13449] = 25'b1111111111110000111111111;
    rom[13450] = 25'b1111111111110001000110111;
    rom[13451] = 25'b1111111111110001001110000;
    rom[13452] = 25'b1111111111110001010101000;
    rom[13453] = 25'b1111111111110001011100001;
    rom[13454] = 25'b1111111111110001100011010;
    rom[13455] = 25'b1111111111110001101010010;
    rom[13456] = 25'b1111111111110001110001011;
    rom[13457] = 25'b1111111111110001111000011;
    rom[13458] = 25'b1111111111110001111111100;
    rom[13459] = 25'b1111111111110010000110101;
    rom[13460] = 25'b1111111111110010001101110;
    rom[13461] = 25'b1111111111110010010100110;
    rom[13462] = 25'b1111111111110010011011111;
    rom[13463] = 25'b1111111111110010100011000;
    rom[13464] = 25'b1111111111110010101010001;
    rom[13465] = 25'b1111111111110010110001010;
    rom[13466] = 25'b1111111111110010111000011;
    rom[13467] = 25'b1111111111110010111111101;
    rom[13468] = 25'b1111111111110011000110101;
    rom[13469] = 25'b1111111111110011001101111;
    rom[13470] = 25'b1111111111110011010101000;
    rom[13471] = 25'b1111111111110011011100001;
    rom[13472] = 25'b1111111111110011100011011;
    rom[13473] = 25'b1111111111110011101010100;
    rom[13474] = 25'b1111111111110011110001101;
    rom[13475] = 25'b1111111111110011111000111;
    rom[13476] = 25'b1111111111110100000000000;
    rom[13477] = 25'b1111111111110100000111010;
    rom[13478] = 25'b1111111111110100001110011;
    rom[13479] = 25'b1111111111110100010101101;
    rom[13480] = 25'b1111111111110100011100110;
    rom[13481] = 25'b1111111111110100100100001;
    rom[13482] = 25'b1111111111110100101011010;
    rom[13483] = 25'b1111111111110100110010100;
    rom[13484] = 25'b1111111111110100111001110;
    rom[13485] = 25'b1111111111110101000000111;
    rom[13486] = 25'b1111111111110101001000010;
    rom[13487] = 25'b1111111111110101001111011;
    rom[13488] = 25'b1111111111110101010110101;
    rom[13489] = 25'b1111111111110101011110000;
    rom[13490] = 25'b1111111111110101100101001;
    rom[13491] = 25'b1111111111110101101100100;
    rom[13492] = 25'b1111111111110101110011110;
    rom[13493] = 25'b1111111111110101111011000;
    rom[13494] = 25'b1111111111110110000010010;
    rom[13495] = 25'b1111111111110110001001101;
    rom[13496] = 25'b1111111111110110010000111;
    rom[13497] = 25'b1111111111110110011000001;
    rom[13498] = 25'b1111111111110110011111011;
    rom[13499] = 25'b1111111111110110100110110;
    rom[13500] = 25'b1111111111110110101110001;
    rom[13501] = 25'b1111111111110110110101011;
    rom[13502] = 25'b1111111111110110111100110;
    rom[13503] = 25'b1111111111110111000100000;
    rom[13504] = 25'b1111111111110111001011011;
    rom[13505] = 25'b1111111111110111010010110;
    rom[13506] = 25'b1111111111110111011010001;
    rom[13507] = 25'b1111111111110111100001100;
    rom[13508] = 25'b1111111111110111101000110;
    rom[13509] = 25'b1111111111110111110000001;
    rom[13510] = 25'b1111111111110111110111100;
    rom[13511] = 25'b1111111111110111111110111;
    rom[13512] = 25'b1111111111111000000110010;
    rom[13513] = 25'b1111111111111000001101101;
    rom[13514] = 25'b1111111111111000010101000;
    rom[13515] = 25'b1111111111111000011100011;
    rom[13516] = 25'b1111111111111000100011110;
    rom[13517] = 25'b1111111111111000101011010;
    rom[13518] = 25'b1111111111111000110010101;
    rom[13519] = 25'b1111111111111000111010000;
    rom[13520] = 25'b1111111111111001000001100;
    rom[13521] = 25'b1111111111111001001000111;
    rom[13522] = 25'b1111111111111001010000010;
    rom[13523] = 25'b1111111111111001010111101;
    rom[13524] = 25'b1111111111111001011111001;
    rom[13525] = 25'b1111111111111001100110101;
    rom[13526] = 25'b1111111111111001101110000;
    rom[13527] = 25'b1111111111111001110101100;
    rom[13528] = 25'b1111111111111001111101000;
    rom[13529] = 25'b1111111111111010000100011;
    rom[13530] = 25'b1111111111111010001011111;
    rom[13531] = 25'b1111111111111010010011011;
    rom[13532] = 25'b1111111111111010011010111;
    rom[13533] = 25'b1111111111111010100010010;
    rom[13534] = 25'b1111111111111010101001110;
    rom[13535] = 25'b1111111111111010110001010;
    rom[13536] = 25'b1111111111111010111000110;
    rom[13537] = 25'b1111111111111011000000010;
    rom[13538] = 25'b1111111111111011000111110;
    rom[13539] = 25'b1111111111111011001111010;
    rom[13540] = 25'b1111111111111011010110110;
    rom[13541] = 25'b1111111111111011011110011;
    rom[13542] = 25'b1111111111111011100101111;
    rom[13543] = 25'b1111111111111011101101011;
    rom[13544] = 25'b1111111111111011110101000;
    rom[13545] = 25'b1111111111111011111100011;
    rom[13546] = 25'b1111111111111100000100000;
    rom[13547] = 25'b1111111111111100001011100;
    rom[13548] = 25'b1111111111111100010011001;
    rom[13549] = 25'b1111111111111100011010101;
    rom[13550] = 25'b1111111111111100100010010;
    rom[13551] = 25'b1111111111111100101001110;
    rom[13552] = 25'b1111111111111100110001011;
    rom[13553] = 25'b1111111111111100111000111;
    rom[13554] = 25'b1111111111111101000000100;
    rom[13555] = 25'b1111111111111101001000001;
    rom[13556] = 25'b1111111111111101001111110;
    rom[13557] = 25'b1111111111111101010111010;
    rom[13558] = 25'b1111111111111101011111000;
    rom[13559] = 25'b1111111111111101100110100;
    rom[13560] = 25'b1111111111111101101110001;
    rom[13561] = 25'b1111111111111101110101110;
    rom[13562] = 25'b1111111111111101111101011;
    rom[13563] = 25'b1111111111111110000101000;
    rom[13564] = 25'b1111111111111110001100101;
    rom[13565] = 25'b1111111111111110010100010;
    rom[13566] = 25'b1111111111111110011011111;
    rom[13567] = 25'b1111111111111110100011101;
    rom[13568] = 25'b1111111111111110101011010;
    rom[13569] = 25'b1111111111111110110010111;
    rom[13570] = 25'b1111111111111110111010100;
    rom[13571] = 25'b1111111111111111000010010;
    rom[13572] = 25'b1111111111111111001001111;
    rom[13573] = 25'b1111111111111111010001100;
    rom[13574] = 25'b1111111111111111011001001;
    rom[13575] = 25'b1111111111111111100000111;
    rom[13576] = 25'b1111111111111111101000101;
    rom[13577] = 25'b1111111111111111110000010;
    rom[13578] = 25'b1111111111111111111000000;
    rom[13579] = 25'b1111111111111111111111101;
    rom[13580] = 25'b0000000000000000000111011;
    rom[13581] = 25'b0000000000000000001111000;
    rom[13582] = 25'b0000000000000000010110110;
    rom[13583] = 25'b0000000000000000011110100;
    rom[13584] = 25'b0000000000000000100110001;
    rom[13585] = 25'b0000000000000000101101111;
    rom[13586] = 25'b0000000000000000110101101;
    rom[13587] = 25'b0000000000000000111101011;
    rom[13588] = 25'b0000000000000001000101001;
    rom[13589] = 25'b0000000000000001001100111;
    rom[13590] = 25'b0000000000000001010100101;
    rom[13591] = 25'b0000000000000001011100011;
    rom[13592] = 25'b0000000000000001100100001;
    rom[13593] = 25'b0000000000000001101011111;
    rom[13594] = 25'b0000000000000001110011101;
    rom[13595] = 25'b0000000000000001111011011;
    rom[13596] = 25'b0000000000000010000011010;
    rom[13597] = 25'b0000000000000010001011000;
    rom[13598] = 25'b0000000000000010010010110;
    rom[13599] = 25'b0000000000000010011010101;
    rom[13600] = 25'b0000000000000010100010011;
    rom[13601] = 25'b0000000000000010101010001;
    rom[13602] = 25'b0000000000000010110001111;
    rom[13603] = 25'b0000000000000010111001110;
    rom[13604] = 25'b0000000000000011000001101;
    rom[13605] = 25'b0000000000000011001001011;
    rom[13606] = 25'b0000000000000011010001010;
    rom[13607] = 25'b0000000000000011011001000;
    rom[13608] = 25'b0000000000000011100000111;
    rom[13609] = 25'b0000000000000011101000110;
    rom[13610] = 25'b0000000000000011110000101;
    rom[13611] = 25'b0000000000000011111000100;
    rom[13612] = 25'b0000000000000100000000010;
    rom[13613] = 25'b0000000000000100001000001;
    rom[13614] = 25'b0000000000000100010000000;
    rom[13615] = 25'b0000000000000100010111111;
    rom[13616] = 25'b0000000000000100011111101;
    rom[13617] = 25'b0000000000000100100111101;
    rom[13618] = 25'b0000000000000100101111100;
    rom[13619] = 25'b0000000000000100110111010;
    rom[13620] = 25'b0000000000000100111111010;
    rom[13621] = 25'b0000000000000101000111001;
    rom[13622] = 25'b0000000000000101001111000;
    rom[13623] = 25'b0000000000000101010110111;
    rom[13624] = 25'b0000000000000101011110110;
    rom[13625] = 25'b0000000000000101100110110;
    rom[13626] = 25'b0000000000000101101110101;
    rom[13627] = 25'b0000000000000101110110100;
    rom[13628] = 25'b0000000000000101111110100;
    rom[13629] = 25'b0000000000000110000110011;
    rom[13630] = 25'b0000000000000110001110010;
    rom[13631] = 25'b0000000000000110010110001;
    rom[13632] = 25'b0000000000000110011110001;
    rom[13633] = 25'b0000000000000110100110000;
    rom[13634] = 25'b0000000000000110101110000;
    rom[13635] = 25'b0000000000000110110101111;
    rom[13636] = 25'b0000000000000110111110000;
    rom[13637] = 25'b0000000000000111000101111;
    rom[13638] = 25'b0000000000000111001101111;
    rom[13639] = 25'b0000000000000111010101110;
    rom[13640] = 25'b0000000000000111011101110;
    rom[13641] = 25'b0000000000000111100101110;
    rom[13642] = 25'b0000000000000111101101101;
    rom[13643] = 25'b0000000000000111110101110;
    rom[13644] = 25'b0000000000000111111101101;
    rom[13645] = 25'b0000000000001000000101101;
    rom[13646] = 25'b0000000000001000001101101;
    rom[13647] = 25'b0000000000001000010101101;
    rom[13648] = 25'b0000000000001000011101101;
    rom[13649] = 25'b0000000000001000100101101;
    rom[13650] = 25'b0000000000001000101101101;
    rom[13651] = 25'b0000000000001000110101101;
    rom[13652] = 25'b0000000000001000111101101;
    rom[13653] = 25'b0000000000001001000101101;
    rom[13654] = 25'b0000000000001001001101101;
    rom[13655] = 25'b0000000000001001010101110;
    rom[13656] = 25'b0000000000001001011101110;
    rom[13657] = 25'b0000000000001001100101110;
    rom[13658] = 25'b0000000000001001101101110;
    rom[13659] = 25'b0000000000001001110101111;
    rom[13660] = 25'b0000000000001001111110000;
    rom[13661] = 25'b0000000000001010000110000;
    rom[13662] = 25'b0000000000001010001110000;
    rom[13663] = 25'b0000000000001010010110000;
    rom[13664] = 25'b0000000000001010011110001;
    rom[13665] = 25'b0000000000001010100110010;
    rom[13666] = 25'b0000000000001010101110010;
    rom[13667] = 25'b0000000000001010110110011;
    rom[13668] = 25'b0000000000001010111110011;
    rom[13669] = 25'b0000000000001011000110100;
    rom[13670] = 25'b0000000000001011001110100;
    rom[13671] = 25'b0000000000001011010110101;
    rom[13672] = 25'b0000000000001011011110110;
    rom[13673] = 25'b0000000000001011100110111;
    rom[13674] = 25'b0000000000001011101111000;
    rom[13675] = 25'b0000000000001011110111001;
    rom[13676] = 25'b0000000000001011111111010;
    rom[13677] = 25'b0000000000001100000111010;
    rom[13678] = 25'b0000000000001100001111011;
    rom[13679] = 25'b0000000000001100010111100;
    rom[13680] = 25'b0000000000001100011111101;
    rom[13681] = 25'b0000000000001100100111110;
    rom[13682] = 25'b0000000000001100101111111;
    rom[13683] = 25'b0000000000001100111000000;
    rom[13684] = 25'b0000000000001101000000010;
    rom[13685] = 25'b0000000000001101001000011;
    rom[13686] = 25'b0000000000001101010000100;
    rom[13687] = 25'b0000000000001101011000101;
    rom[13688] = 25'b0000000000001101100000110;
    rom[13689] = 25'b0000000000001101101000111;
    rom[13690] = 25'b0000000000001101110001000;
    rom[13691] = 25'b0000000000001101111001001;
    rom[13692] = 25'b0000000000001110000001011;
    rom[13693] = 25'b0000000000001110001001100;
    rom[13694] = 25'b0000000000001110010001110;
    rom[13695] = 25'b0000000000001110011001111;
    rom[13696] = 25'b0000000000001110100010001;
    rom[13697] = 25'b0000000000001110101010010;
    rom[13698] = 25'b0000000000001110110010011;
    rom[13699] = 25'b0000000000001110111010101;
    rom[13700] = 25'b0000000000001111000010111;
    rom[13701] = 25'b0000000000001111001011001;
    rom[13702] = 25'b0000000000001111010011010;
    rom[13703] = 25'b0000000000001111011011011;
    rom[13704] = 25'b0000000000001111100011101;
    rom[13705] = 25'b0000000000001111101011111;
    rom[13706] = 25'b0000000000001111110100001;
    rom[13707] = 25'b0000000000001111111100010;
    rom[13708] = 25'b0000000000010000000100100;
    rom[13709] = 25'b0000000000010000001100110;
    rom[13710] = 25'b0000000000010000010101000;
    rom[13711] = 25'b0000000000010000011101001;
    rom[13712] = 25'b0000000000010000100101100;
    rom[13713] = 25'b0000000000010000101101101;
    rom[13714] = 25'b0000000000010000110101111;
    rom[13715] = 25'b0000000000010000111110001;
    rom[13716] = 25'b0000000000010001000110011;
    rom[13717] = 25'b0000000000010001001110101;
    rom[13718] = 25'b0000000000010001010110111;
    rom[13719] = 25'b0000000000010001011111001;
    rom[13720] = 25'b0000000000010001100111011;
    rom[13721] = 25'b0000000000010001101111110;
    rom[13722] = 25'b0000000000010001110111111;
    rom[13723] = 25'b0000000000010010000000010;
    rom[13724] = 25'b0000000000010010001000100;
    rom[13725] = 25'b0000000000010010010000110;
    rom[13726] = 25'b0000000000010010011001001;
    rom[13727] = 25'b0000000000010010100001011;
    rom[13728] = 25'b0000000000010010101001101;
    rom[13729] = 25'b0000000000010010110001111;
    rom[13730] = 25'b0000000000010010111010010;
    rom[13731] = 25'b0000000000010011000010100;
    rom[13732] = 25'b0000000000010011001010111;
    rom[13733] = 25'b0000000000010011010011001;
    rom[13734] = 25'b0000000000010011011011100;
    rom[13735] = 25'b0000000000010011100011110;
    rom[13736] = 25'b0000000000010011101100001;
    rom[13737] = 25'b0000000000010011110100011;
    rom[13738] = 25'b0000000000010011111100110;
    rom[13739] = 25'b0000000000010100000101000;
    rom[13740] = 25'b0000000000010100001101011;
    rom[13741] = 25'b0000000000010100010101101;
    rom[13742] = 25'b0000000000010100011110001;
    rom[13743] = 25'b0000000000010100100110011;
    rom[13744] = 25'b0000000000010100101110101;
    rom[13745] = 25'b0000000000010100110111000;
    rom[13746] = 25'b0000000000010100111111011;
    rom[13747] = 25'b0000000000010101000111110;
    rom[13748] = 25'b0000000000010101010000001;
    rom[13749] = 25'b0000000000010101011000011;
    rom[13750] = 25'b0000000000010101100000111;
    rom[13751] = 25'b0000000000010101101001001;
    rom[13752] = 25'b0000000000010101110001100;
    rom[13753] = 25'b0000000000010101111001111;
    rom[13754] = 25'b0000000000010110000010010;
    rom[13755] = 25'b0000000000010110001010101;
    rom[13756] = 25'b0000000000010110010011000;
    rom[13757] = 25'b0000000000010110011011011;
    rom[13758] = 25'b0000000000010110100011110;
    rom[13759] = 25'b0000000000010110101100001;
    rom[13760] = 25'b0000000000010110110100100;
    rom[13761] = 25'b0000000000010110111100111;
    rom[13762] = 25'b0000000000010111000101011;
    rom[13763] = 25'b0000000000010111001101110;
    rom[13764] = 25'b0000000000010111010110001;
    rom[13765] = 25'b0000000000010111011110100;
    rom[13766] = 25'b0000000000010111100111000;
    rom[13767] = 25'b0000000000010111101111011;
    rom[13768] = 25'b0000000000010111110111110;
    rom[13769] = 25'b0000000000011000000000001;
    rom[13770] = 25'b0000000000011000001000100;
    rom[13771] = 25'b0000000000011000010001000;
    rom[13772] = 25'b0000000000011000011001011;
    rom[13773] = 25'b0000000000011000100001111;
    rom[13774] = 25'b0000000000011000101010010;
    rom[13775] = 25'b0000000000011000110010101;
    rom[13776] = 25'b0000000000011000111011001;
    rom[13777] = 25'b0000000000011001000011101;
    rom[13778] = 25'b0000000000011001001100000;
    rom[13779] = 25'b0000000000011001010100011;
    rom[13780] = 25'b0000000000011001011100111;
    rom[13781] = 25'b0000000000011001100101010;
    rom[13782] = 25'b0000000000011001101101110;
    rom[13783] = 25'b0000000000011001110110010;
    rom[13784] = 25'b0000000000011001111110110;
    rom[13785] = 25'b0000000000011010000111001;
    rom[13786] = 25'b0000000000011010001111101;
    rom[13787] = 25'b0000000000011010011000001;
    rom[13788] = 25'b0000000000011010100000100;
    rom[13789] = 25'b0000000000011010101001000;
    rom[13790] = 25'b0000000000011010110001100;
    rom[13791] = 25'b0000000000011010111001111;
    rom[13792] = 25'b0000000000011011000010011;
    rom[13793] = 25'b0000000000011011001010111;
    rom[13794] = 25'b0000000000011011010011011;
    rom[13795] = 25'b0000000000011011011011110;
    rom[13796] = 25'b0000000000011011100100010;
    rom[13797] = 25'b0000000000011011101100110;
    rom[13798] = 25'b0000000000011011110101010;
    rom[13799] = 25'b0000000000011011111101110;
    rom[13800] = 25'b0000000000011100000110010;
    rom[13801] = 25'b0000000000011100001110110;
    rom[13802] = 25'b0000000000011100010111010;
    rom[13803] = 25'b0000000000011100011111110;
    rom[13804] = 25'b0000000000011100101000010;
    rom[13805] = 25'b0000000000011100110000110;
    rom[13806] = 25'b0000000000011100111001010;
    rom[13807] = 25'b0000000000011101000001111;
    rom[13808] = 25'b0000000000011101001010011;
    rom[13809] = 25'b0000000000011101010010111;
    rom[13810] = 25'b0000000000011101011011011;
    rom[13811] = 25'b0000000000011101100011111;
    rom[13812] = 25'b0000000000011101101100100;
    rom[13813] = 25'b0000000000011101110101000;
    rom[13814] = 25'b0000000000011101111101100;
    rom[13815] = 25'b0000000000011110000110000;
    rom[13816] = 25'b0000000000011110001110100;
    rom[13817] = 25'b0000000000011110010111000;
    rom[13818] = 25'b0000000000011110011111101;
    rom[13819] = 25'b0000000000011110101000001;
    rom[13820] = 25'b0000000000011110110000110;
    rom[13821] = 25'b0000000000011110111001010;
    rom[13822] = 25'b0000000000011111000001110;
    rom[13823] = 25'b0000000000011111001010010;
    rom[13824] = 25'b0000000000011111010010111;
    rom[13825] = 25'b0000000000011111011011100;
    rom[13826] = 25'b0000000000011111100100000;
    rom[13827] = 25'b0000000000011111101100101;
    rom[13828] = 25'b0000000000011111110101001;
    rom[13829] = 25'b0000000000011111111101101;
    rom[13830] = 25'b0000000000100000000110010;
    rom[13831] = 25'b0000000000100000001110111;
    rom[13832] = 25'b0000000000100000010111011;
    rom[13833] = 25'b0000000000100000100000000;
    rom[13834] = 25'b0000000000100000101000100;
    rom[13835] = 25'b0000000000100000110001001;
    rom[13836] = 25'b0000000000100000111001110;
    rom[13837] = 25'b0000000000100001000010011;
    rom[13838] = 25'b0000000000100001001010110;
    rom[13839] = 25'b0000000000100001010011011;
    rom[13840] = 25'b0000000000100001011100000;
    rom[13841] = 25'b0000000000100001100100101;
    rom[13842] = 25'b0000000000100001101101001;
    rom[13843] = 25'b0000000000100001110101110;
    rom[13844] = 25'b0000000000100001111110011;
    rom[13845] = 25'b0000000000100010000111000;
    rom[13846] = 25'b0000000000100010001111100;
    rom[13847] = 25'b0000000000100010011000010;
    rom[13848] = 25'b0000000000100010100000111;
    rom[13849] = 25'b0000000000100010101001011;
    rom[13850] = 25'b0000000000100010110010000;
    rom[13851] = 25'b0000000000100010111010101;
    rom[13852] = 25'b0000000000100011000011001;
    rom[13853] = 25'b0000000000100011001011111;
    rom[13854] = 25'b0000000000100011010100100;
    rom[13855] = 25'b0000000000100011011101000;
    rom[13856] = 25'b0000000000100011100101101;
    rom[13857] = 25'b0000000000100011101110011;
    rom[13858] = 25'b0000000000100011110110111;
    rom[13859] = 25'b0000000000100011111111100;
    rom[13860] = 25'b0000000000100100001000010;
    rom[13861] = 25'b0000000000100100010000110;
    rom[13862] = 25'b0000000000100100011001100;
    rom[13863] = 25'b0000000000100100100010001;
    rom[13864] = 25'b0000000000100100101010101;
    rom[13865] = 25'b0000000000100100110011011;
    rom[13866] = 25'b0000000000100100111011111;
    rom[13867] = 25'b0000000000100101000100101;
    rom[13868] = 25'b0000000000100101001101010;
    rom[13869] = 25'b0000000000100101010101111;
    rom[13870] = 25'b0000000000100101011110100;
    rom[13871] = 25'b0000000000100101100111001;
    rom[13872] = 25'b0000000000100101101111111;
    rom[13873] = 25'b0000000000100101111000100;
    rom[13874] = 25'b0000000000100110000001001;
    rom[13875] = 25'b0000000000100110001001110;
    rom[13876] = 25'b0000000000100110010010011;
    rom[13877] = 25'b0000000000100110011011001;
    rom[13878] = 25'b0000000000100110100011110;
    rom[13879] = 25'b0000000000100110101100011;
    rom[13880] = 25'b0000000000100110110101000;
    rom[13881] = 25'b0000000000100110111101110;
    rom[13882] = 25'b0000000000100111000110011;
    rom[13883] = 25'b0000000000100111001111000;
    rom[13884] = 25'b0000000000100111010111110;
    rom[13885] = 25'b0000000000100111100000011;
    rom[13886] = 25'b0000000000100111101001001;
    rom[13887] = 25'b0000000000100111110001110;
    rom[13888] = 25'b0000000000100111111010011;
    rom[13889] = 25'b0000000000101000000011000;
    rom[13890] = 25'b0000000000101000001011110;
    rom[13891] = 25'b0000000000101000010100011;
    rom[13892] = 25'b0000000000101000011101001;
    rom[13893] = 25'b0000000000101000100101110;
    rom[13894] = 25'b0000000000101000101110100;
    rom[13895] = 25'b0000000000101000110111001;
    rom[13896] = 25'b0000000000101000111111111;
    rom[13897] = 25'b0000000000101001001000100;
    rom[13898] = 25'b0000000000101001010001010;
    rom[13899] = 25'b0000000000101001011001111;
    rom[13900] = 25'b0000000000101001100010101;
    rom[13901] = 25'b0000000000101001101011010;
    rom[13902] = 25'b0000000000101001110100000;
    rom[13903] = 25'b0000000000101001111100101;
    rom[13904] = 25'b0000000000101010000101011;
    rom[13905] = 25'b0000000000101010001110001;
    rom[13906] = 25'b0000000000101010010110110;
    rom[13907] = 25'b0000000000101010011111100;
    rom[13908] = 25'b0000000000101010101000001;
    rom[13909] = 25'b0000000000101010110000111;
    rom[13910] = 25'b0000000000101010111001100;
    rom[13911] = 25'b0000000000101011000010010;
    rom[13912] = 25'b0000000000101011001011000;
    rom[13913] = 25'b0000000000101011010011101;
    rom[13914] = 25'b0000000000101011011100011;
    rom[13915] = 25'b0000000000101011100101001;
    rom[13916] = 25'b0000000000101011101101111;
    rom[13917] = 25'b0000000000101011110110100;
    rom[13918] = 25'b0000000000101011111111001;
    rom[13919] = 25'b0000000000101100001000000;
    rom[13920] = 25'b0000000000101100010000101;
    rom[13921] = 25'b0000000000101100011001011;
    rom[13922] = 25'b0000000000101100100010001;
    rom[13923] = 25'b0000000000101100101010110;
    rom[13924] = 25'b0000000000101100110011100;
    rom[13925] = 25'b0000000000101100111100010;
    rom[13926] = 25'b0000000000101101000101000;
    rom[13927] = 25'b0000000000101101001101110;
    rom[13928] = 25'b0000000000101101010110011;
    rom[13929] = 25'b0000000000101101011111001;
    rom[13930] = 25'b0000000000101101100111111;
    rom[13931] = 25'b0000000000101101110000100;
    rom[13932] = 25'b0000000000101101111001011;
    rom[13933] = 25'b0000000000101110000010000;
    rom[13934] = 25'b0000000000101110001010110;
    rom[13935] = 25'b0000000000101110010011100;
    rom[13936] = 25'b0000000000101110011100010;
    rom[13937] = 25'b0000000000101110100101000;
    rom[13938] = 25'b0000000000101110101101110;
    rom[13939] = 25'b0000000000101110110110011;
    rom[13940] = 25'b0000000000101110111111001;
    rom[13941] = 25'b0000000000101111001000000;
    rom[13942] = 25'b0000000000101111010000101;
    rom[13943] = 25'b0000000000101111011001011;
    rom[13944] = 25'b0000000000101111100010001;
    rom[13945] = 25'b0000000000101111101010111;
    rom[13946] = 25'b0000000000101111110011101;
    rom[13947] = 25'b0000000000101111111100011;
    rom[13948] = 25'b0000000000110000000101001;
    rom[13949] = 25'b0000000000110000001101111;
    rom[13950] = 25'b0000000000110000010110101;
    rom[13951] = 25'b0000000000110000011111011;
    rom[13952] = 25'b0000000000110000101000000;
    rom[13953] = 25'b0000000000110000110000111;
    rom[13954] = 25'b0000000000110000111001101;
    rom[13955] = 25'b0000000000110001000010010;
    rom[13956] = 25'b0000000000110001001011001;
    rom[13957] = 25'b0000000000110001010011111;
    rom[13958] = 25'b0000000000110001011100100;
    rom[13959] = 25'b0000000000110001100101011;
    rom[13960] = 25'b0000000000110001101110001;
    rom[13961] = 25'b0000000000110001110110110;
    rom[13962] = 25'b0000000000110001111111101;
    rom[13963] = 25'b0000000000110010001000011;
    rom[13964] = 25'b0000000000110010010001001;
    rom[13965] = 25'b0000000000110010011001110;
    rom[13966] = 25'b0000000000110010100010101;
    rom[13967] = 25'b0000000000110010101011011;
    rom[13968] = 25'b0000000000110010110100001;
    rom[13969] = 25'b0000000000110010111100111;
    rom[13970] = 25'b0000000000110011000101101;
    rom[13971] = 25'b0000000000110011001110011;
    rom[13972] = 25'b0000000000110011010111001;
    rom[13973] = 25'b0000000000110011100000000;
    rom[13974] = 25'b0000000000110011101000101;
    rom[13975] = 25'b0000000000110011110001011;
    rom[13976] = 25'b0000000000110011111010001;
    rom[13977] = 25'b0000000000110100000011000;
    rom[13978] = 25'b0000000000110100001011110;
    rom[13979] = 25'b0000000000110100010100100;
    rom[13980] = 25'b0000000000110100011101010;
    rom[13981] = 25'b0000000000110100100110000;
    rom[13982] = 25'b0000000000110100101110110;
    rom[13983] = 25'b0000000000110100110111100;
    rom[13984] = 25'b0000000000110101000000011;
    rom[13985] = 25'b0000000000110101001001001;
    rom[13986] = 25'b0000000000110101010001110;
    rom[13987] = 25'b0000000000110101011010100;
    rom[13988] = 25'b0000000000110101100011011;
    rom[13989] = 25'b0000000000110101101100001;
    rom[13990] = 25'b0000000000110101110100111;
    rom[13991] = 25'b0000000000110101111101101;
    rom[13992] = 25'b0000000000110110000110100;
    rom[13993] = 25'b0000000000110110001111010;
    rom[13994] = 25'b0000000000110110010111111;
    rom[13995] = 25'b0000000000110110100000110;
    rom[13996] = 25'b0000000000110110101001100;
    rom[13997] = 25'b0000000000110110110010010;
    rom[13998] = 25'b0000000000110110111011000;
    rom[13999] = 25'b0000000000110111000011110;
    rom[14000] = 25'b0000000000110111001100101;
    rom[14001] = 25'b0000000000110111010101011;
    rom[14002] = 25'b0000000000110111011110001;
    rom[14003] = 25'b0000000000110111100110111;
    rom[14004] = 25'b0000000000110111101111101;
    rom[14005] = 25'b0000000000110111111000011;
    rom[14006] = 25'b0000000000111000000001001;
    rom[14007] = 25'b0000000000111000001001111;
    rom[14008] = 25'b0000000000111000010010110;
    rom[14009] = 25'b0000000000111000011011100;
    rom[14010] = 25'b0000000000111000100100010;
    rom[14011] = 25'b0000000000111000101101000;
    rom[14012] = 25'b0000000000111000110101111;
    rom[14013] = 25'b0000000000111000111110101;
    rom[14014] = 25'b0000000000111001000111010;
    rom[14015] = 25'b0000000000111001010000001;
    rom[14016] = 25'b0000000000111001011000111;
    rom[14017] = 25'b0000000000111001100001101;
    rom[14018] = 25'b0000000000111001101010011;
    rom[14019] = 25'b0000000000111001110011001;
    rom[14020] = 25'b0000000000111001111100000;
    rom[14021] = 25'b0000000000111010000100110;
    rom[14022] = 25'b0000000000111010001101100;
    rom[14023] = 25'b0000000000111010010110010;
    rom[14024] = 25'b0000000000111010011111001;
    rom[14025] = 25'b0000000000111010100111110;
    rom[14026] = 25'b0000000000111010110000100;
    rom[14027] = 25'b0000000000111010111001011;
    rom[14028] = 25'b0000000000111011000010001;
    rom[14029] = 25'b0000000000111011001010111;
    rom[14030] = 25'b0000000000111011010011101;
    rom[14031] = 25'b0000000000111011011100011;
    rom[14032] = 25'b0000000000111011100101010;
    rom[14033] = 25'b0000000000111011101110000;
    rom[14034] = 25'b0000000000111011110110110;
    rom[14035] = 25'b0000000000111011111111100;
    rom[14036] = 25'b0000000000111100001000010;
    rom[14037] = 25'b0000000000111100010001000;
    rom[14038] = 25'b0000000000111100011001110;
    rom[14039] = 25'b0000000000111100100010101;
    rom[14040] = 25'b0000000000111100101011011;
    rom[14041] = 25'b0000000000111100110100001;
    rom[14042] = 25'b0000000000111100111100111;
    rom[14043] = 25'b0000000000111101000101101;
    rom[14044] = 25'b0000000000111101001110011;
    rom[14045] = 25'b0000000000111101010111001;
    rom[14046] = 25'b0000000000111101011111111;
    rom[14047] = 25'b0000000000111101101000110;
    rom[14048] = 25'b0000000000111101110001100;
    rom[14049] = 25'b0000000000111101111010001;
    rom[14050] = 25'b0000000000111110000011000;
    rom[14051] = 25'b0000000000111110001011110;
    rom[14052] = 25'b0000000000111110010100100;
    rom[14053] = 25'b0000000000111110011101010;
    rom[14054] = 25'b0000000000111110100110000;
    rom[14055] = 25'b0000000000111110101110110;
    rom[14056] = 25'b0000000000111110110111100;
    rom[14057] = 25'b0000000000111111000000010;
    rom[14058] = 25'b0000000000111111001001001;
    rom[14059] = 25'b0000000000111111010001110;
    rom[14060] = 25'b0000000000111111011010100;
    rom[14061] = 25'b0000000000111111100011011;
    rom[14062] = 25'b0000000000111111101100001;
    rom[14063] = 25'b0000000000111111110100111;
    rom[14064] = 25'b0000000000111111111101100;
    rom[14065] = 25'b0000000001000000000110011;
    rom[14066] = 25'b0000000001000000001111001;
    rom[14067] = 25'b0000000001000000010111110;
    rom[14068] = 25'b0000000001000000100000101;
    rom[14069] = 25'b0000000001000000101001011;
    rom[14070] = 25'b0000000001000000110010001;
    rom[14071] = 25'b0000000001000000111010111;
    rom[14072] = 25'b0000000001000001000011101;
    rom[14073] = 25'b0000000001000001001100011;
    rom[14074] = 25'b0000000001000001010101000;
    rom[14075] = 25'b0000000001000001011101111;
    rom[14076] = 25'b0000000001000001100110101;
    rom[14077] = 25'b0000000001000001101111010;
    rom[14078] = 25'b0000000001000001111000001;
    rom[14079] = 25'b0000000001000010000000111;
    rom[14080] = 25'b0000000001000010001001100;
    rom[14081] = 25'b0000000001000010010010011;
    rom[14082] = 25'b0000000001000010011011000;
    rom[14083] = 25'b0000000001000010100011110;
    rom[14084] = 25'b0000000001000010101100101;
    rom[14085] = 25'b0000000001000010110101010;
    rom[14086] = 25'b0000000001000010111110000;
    rom[14087] = 25'b0000000001000011000110110;
    rom[14088] = 25'b0000000001000011001111100;
    rom[14089] = 25'b0000000001000011011000001;
    rom[14090] = 25'b0000000001000011100001000;
    rom[14091] = 25'b0000000001000011101001101;
    rom[14092] = 25'b0000000001000011110010011;
    rom[14093] = 25'b0000000001000011111011001;
    rom[14094] = 25'b0000000001000100000011111;
    rom[14095] = 25'b0000000001000100001100101;
    rom[14096] = 25'b0000000001000100010101011;
    rom[14097] = 25'b0000000001000100011110000;
    rom[14098] = 25'b0000000001000100100110110;
    rom[14099] = 25'b0000000001000100101111100;
    rom[14100] = 25'b0000000001000100111000010;
    rom[14101] = 25'b0000000001000101000001000;
    rom[14102] = 25'b0000000001000101001001101;
    rom[14103] = 25'b0000000001000101010010011;
    rom[14104] = 25'b0000000001000101011011001;
    rom[14105] = 25'b0000000001000101100011110;
    rom[14106] = 25'b0000000001000101101100101;
    rom[14107] = 25'b0000000001000101110101010;
    rom[14108] = 25'b0000000001000101111110000;
    rom[14109] = 25'b0000000001000110000110110;
    rom[14110] = 25'b0000000001000110001111011;
    rom[14111] = 25'b0000000001000110011000001;
    rom[14112] = 25'b0000000001000110100000111;
    rom[14113] = 25'b0000000001000110101001100;
    rom[14114] = 25'b0000000001000110110010010;
    rom[14115] = 25'b0000000001000110111010111;
    rom[14116] = 25'b0000000001000111000011101;
    rom[14117] = 25'b0000000001000111001100011;
    rom[14118] = 25'b0000000001000111010101001;
    rom[14119] = 25'b0000000001000111011101110;
    rom[14120] = 25'b0000000001000111100110100;
    rom[14121] = 25'b0000000001000111101111001;
    rom[14122] = 25'b0000000001000111110111110;
    rom[14123] = 25'b0000000001001000000000101;
    rom[14124] = 25'b0000000001001000001001010;
    rom[14125] = 25'b0000000001001000010010000;
    rom[14126] = 25'b0000000001001000011010101;
    rom[14127] = 25'b0000000001001000100011011;
    rom[14128] = 25'b0000000001001000101100000;
    rom[14129] = 25'b0000000001001000110100110;
    rom[14130] = 25'b0000000001001000111101011;
    rom[14131] = 25'b0000000001001001000110001;
    rom[14132] = 25'b0000000001001001001110110;
    rom[14133] = 25'b0000000001001001010111011;
    rom[14134] = 25'b0000000001001001100000001;
    rom[14135] = 25'b0000000001001001101000110;
    rom[14136] = 25'b0000000001001001110001011;
    rom[14137] = 25'b0000000001001001111010001;
    rom[14138] = 25'b0000000001001010000010110;
    rom[14139] = 25'b0000000001001010001011100;
    rom[14140] = 25'b0000000001001010010100001;
    rom[14141] = 25'b0000000001001010011100111;
    rom[14142] = 25'b0000000001001010100101100;
    rom[14143] = 25'b0000000001001010101110001;
    rom[14144] = 25'b0000000001001010110110110;
    rom[14145] = 25'b0000000001001010111111100;
    rom[14146] = 25'b0000000001001011001000001;
    rom[14147] = 25'b0000000001001011010000110;
    rom[14148] = 25'b0000000001001011011001011;
    rom[14149] = 25'b0000000001001011100010001;
    rom[14150] = 25'b0000000001001011101010110;
    rom[14151] = 25'b0000000001001011110011011;
    rom[14152] = 25'b0000000001001011111100001;
    rom[14153] = 25'b0000000001001100000100101;
    rom[14154] = 25'b0000000001001100001101011;
    rom[14155] = 25'b0000000001001100010110000;
    rom[14156] = 25'b0000000001001100011110101;
    rom[14157] = 25'b0000000001001100100111010;
    rom[14158] = 25'b0000000001001100101111111;
    rom[14159] = 25'b0000000001001100111000100;
    rom[14160] = 25'b0000000001001101000001001;
    rom[14161] = 25'b0000000001001101001001110;
    rom[14162] = 25'b0000000001001101010010100;
    rom[14163] = 25'b0000000001001101011011000;
    rom[14164] = 25'b0000000001001101100011101;
    rom[14165] = 25'b0000000001001101101100011;
    rom[14166] = 25'b0000000001001101110100111;
    rom[14167] = 25'b0000000001001101111101100;
    rom[14168] = 25'b0000000001001110000110010;
    rom[14169] = 25'b0000000001001110001110110;
    rom[14170] = 25'b0000000001001110010111011;
    rom[14171] = 25'b0000000001001110100000000;
    rom[14172] = 25'b0000000001001110101000101;
    rom[14173] = 25'b0000000001001110110001010;
    rom[14174] = 25'b0000000001001110111001111;
    rom[14175] = 25'b0000000001001111000010011;
    rom[14176] = 25'b0000000001001111001011000;
    rom[14177] = 25'b0000000001001111010011101;
    rom[14178] = 25'b0000000001001111011100010;
    rom[14179] = 25'b0000000001001111100100110;
    rom[14180] = 25'b0000000001001111101101011;
    rom[14181] = 25'b0000000001001111110110000;
    rom[14182] = 25'b0000000001001111111110101;
    rom[14183] = 25'b0000000001010000000111001;
    rom[14184] = 25'b0000000001010000001111110;
    rom[14185] = 25'b0000000001010000011000011;
    rom[14186] = 25'b0000000001010000100001000;
    rom[14187] = 25'b0000000001010000101001100;
    rom[14188] = 25'b0000000001010000110010001;
    rom[14189] = 25'b0000000001010000111010110;
    rom[14190] = 25'b0000000001010001000011010;
    rom[14191] = 25'b0000000001010001001011110;
    rom[14192] = 25'b0000000001010001010100011;
    rom[14193] = 25'b0000000001010001011101000;
    rom[14194] = 25'b0000000001010001100101100;
    rom[14195] = 25'b0000000001010001101110001;
    rom[14196] = 25'b0000000001010001110110101;
    rom[14197] = 25'b0000000001010001111111001;
    rom[14198] = 25'b0000000001010010000111110;
    rom[14199] = 25'b0000000001010010010000010;
    rom[14200] = 25'b0000000001010010011000111;
    rom[14201] = 25'b0000000001010010100001011;
    rom[14202] = 25'b0000000001010010101010000;
    rom[14203] = 25'b0000000001010010110010011;
    rom[14204] = 25'b0000000001010010111011000;
    rom[14205] = 25'b0000000001010011000011100;
    rom[14206] = 25'b0000000001010011001100000;
    rom[14207] = 25'b0000000001010011010100101;
    rom[14208] = 25'b0000000001010011011101001;
    rom[14209] = 25'b0000000001010011100101101;
    rom[14210] = 25'b0000000001010011101110010;
    rom[14211] = 25'b0000000001010011110110110;
    rom[14212] = 25'b0000000001010011111111010;
    rom[14213] = 25'b0000000001010100000111110;
    rom[14214] = 25'b0000000001010100010000010;
    rom[14215] = 25'b0000000001010100011000110;
    rom[14216] = 25'b0000000001010100100001010;
    rom[14217] = 25'b0000000001010100101001110;
    rom[14218] = 25'b0000000001010100110010010;
    rom[14219] = 25'b0000000001010100111010110;
    rom[14220] = 25'b0000000001010101000011010;
    rom[14221] = 25'b0000000001010101001011110;
    rom[14222] = 25'b0000000001010101010100010;
    rom[14223] = 25'b0000000001010101011100110;
    rom[14224] = 25'b0000000001010101100101001;
    rom[14225] = 25'b0000000001010101101101101;
    rom[14226] = 25'b0000000001010101110110001;
    rom[14227] = 25'b0000000001010101111110101;
    rom[14228] = 25'b0000000001010110000111001;
    rom[14229] = 25'b0000000001010110001111101;
    rom[14230] = 25'b0000000001010110011000001;
    rom[14231] = 25'b0000000001010110100000101;
    rom[14232] = 25'b0000000001010110101001000;
    rom[14233] = 25'b0000000001010110110001100;
    rom[14234] = 25'b0000000001010110111001111;
    rom[14235] = 25'b0000000001010111000010011;
    rom[14236] = 25'b0000000001010111001010110;
    rom[14237] = 25'b0000000001010111010011010;
    rom[14238] = 25'b0000000001010111011011110;
    rom[14239] = 25'b0000000001010111100100001;
    rom[14240] = 25'b0000000001010111101100101;
    rom[14241] = 25'b0000000001010111110101000;
    rom[14242] = 25'b0000000001010111111101100;
    rom[14243] = 25'b0000000001011000000101111;
    rom[14244] = 25'b0000000001011000001110010;
    rom[14245] = 25'b0000000001011000010110110;
    rom[14246] = 25'b0000000001011000011111010;
    rom[14247] = 25'b0000000001011000100111101;
    rom[14248] = 25'b0000000001011000110000000;
    rom[14249] = 25'b0000000001011000111000011;
    rom[14250] = 25'b0000000001011001000000111;
    rom[14251] = 25'b0000000001011001001001010;
    rom[14252] = 25'b0000000001011001010001101;
    rom[14253] = 25'b0000000001011001011010000;
    rom[14254] = 25'b0000000001011001100010100;
    rom[14255] = 25'b0000000001011001101010111;
    rom[14256] = 25'b0000000001011001110011010;
    rom[14257] = 25'b0000000001011001111011101;
    rom[14258] = 25'b0000000001011010000100000;
    rom[14259] = 25'b0000000001011010001100011;
    rom[14260] = 25'b0000000001011010010100110;
    rom[14261] = 25'b0000000001011010011101001;
    rom[14262] = 25'b0000000001011010100101100;
    rom[14263] = 25'b0000000001011010101101111;
    rom[14264] = 25'b0000000001011010110110010;
    rom[14265] = 25'b0000000001011010111110101;
    rom[14266] = 25'b0000000001011011000110111;
    rom[14267] = 25'b0000000001011011001111011;
    rom[14268] = 25'b0000000001011011010111101;
    rom[14269] = 25'b0000000001011011100000000;
    rom[14270] = 25'b0000000001011011101000011;
    rom[14271] = 25'b0000000001011011110000101;
    rom[14272] = 25'b0000000001011011111001000;
    rom[14273] = 25'b0000000001011100000001011;
    rom[14274] = 25'b0000000001011100001001110;
    rom[14275] = 25'b0000000001011100010010000;
    rom[14276] = 25'b0000000001011100011010011;
    rom[14277] = 25'b0000000001011100100010101;
    rom[14278] = 25'b0000000001011100101011000;
    rom[14279] = 25'b0000000001011100110011010;
    rom[14280] = 25'b0000000001011100111011101;
    rom[14281] = 25'b0000000001011101000011111;
    rom[14282] = 25'b0000000001011101001100010;
    rom[14283] = 25'b0000000001011101010100100;
    rom[14284] = 25'b0000000001011101011100111;
    rom[14285] = 25'b0000000001011101100101001;
    rom[14286] = 25'b0000000001011101101101011;
    rom[14287] = 25'b0000000001011101110101101;
    rom[14288] = 25'b0000000001011101111110000;
    rom[14289] = 25'b0000000001011110000110001;
    rom[14290] = 25'b0000000001011110001110100;
    rom[14291] = 25'b0000000001011110010110110;
    rom[14292] = 25'b0000000001011110011111000;
    rom[14293] = 25'b0000000001011110100111011;
    rom[14294] = 25'b0000000001011110101111100;
    rom[14295] = 25'b0000000001011110110111110;
    rom[14296] = 25'b0000000001011111000000001;
    rom[14297] = 25'b0000000001011111001000010;
    rom[14298] = 25'b0000000001011111010000100;
    rom[14299] = 25'b0000000001011111011000111;
    rom[14300] = 25'b0000000001011111100001000;
    rom[14301] = 25'b0000000001011111101001010;
    rom[14302] = 25'b0000000001011111110001100;
    rom[14303] = 25'b0000000001011111111001110;
    rom[14304] = 25'b0000000001100000000001111;
    rom[14305] = 25'b0000000001100000001010001;
    rom[14306] = 25'b0000000001100000010010011;
    rom[14307] = 25'b0000000001100000011010101;
    rom[14308] = 25'b0000000001100000100010110;
    rom[14309] = 25'b0000000001100000101011000;
    rom[14310] = 25'b0000000001100000110011001;
    rom[14311] = 25'b0000000001100000111011011;
    rom[14312] = 25'b0000000001100001000011101;
    rom[14313] = 25'b0000000001100001001011110;
    rom[14314] = 25'b0000000001100001010011111;
    rom[14315] = 25'b0000000001100001011100001;
    rom[14316] = 25'b0000000001100001100100010;
    rom[14317] = 25'b0000000001100001101100100;
    rom[14318] = 25'b0000000001100001110100101;
    rom[14319] = 25'b0000000001100001111100111;
    rom[14320] = 25'b0000000001100010000101000;
    rom[14321] = 25'b0000000001100010001101001;
    rom[14322] = 25'b0000000001100010010101010;
    rom[14323] = 25'b0000000001100010011101011;
    rom[14324] = 25'b0000000001100010100101100;
    rom[14325] = 25'b0000000001100010101101101;
    rom[14326] = 25'b0000000001100010110101110;
    rom[14327] = 25'b0000000001100010111101111;
    rom[14328] = 25'b0000000001100011000110000;
    rom[14329] = 25'b0000000001100011001110001;
    rom[14330] = 25'b0000000001100011010110010;
    rom[14331] = 25'b0000000001100011011110011;
    rom[14332] = 25'b0000000001100011100110100;
    rom[14333] = 25'b0000000001100011101110101;
    rom[14334] = 25'b0000000001100011110110110;
    rom[14335] = 25'b0000000001100011111110111;
    rom[14336] = 25'b0000000001100100000110111;
    rom[14337] = 25'b0000000001100100001111000;
    rom[14338] = 25'b0000000001100100010111001;
    rom[14339] = 25'b0000000001100100011111001;
    rom[14340] = 25'b0000000001100100100111001;
    rom[14341] = 25'b0000000001100100101111010;
    rom[14342] = 25'b0000000001100100110111011;
    rom[14343] = 25'b0000000001100100111111100;
    rom[14344] = 25'b0000000001100101000111100;
    rom[14345] = 25'b0000000001100101001111100;
    rom[14346] = 25'b0000000001100101010111100;
    rom[14347] = 25'b0000000001100101011111101;
    rom[14348] = 25'b0000000001100101100111101;
    rom[14349] = 25'b0000000001100101101111101;
    rom[14350] = 25'b0000000001100101110111101;
    rom[14351] = 25'b0000000001100101111111110;
    rom[14352] = 25'b0000000001100110000111110;
    rom[14353] = 25'b0000000001100110001111110;
    rom[14354] = 25'b0000000001100110010111110;
    rom[14355] = 25'b0000000001100110011111110;
    rom[14356] = 25'b0000000001100110100111110;
    rom[14357] = 25'b0000000001100110101111110;
    rom[14358] = 25'b0000000001100110110111110;
    rom[14359] = 25'b0000000001100110111111110;
    rom[14360] = 25'b0000000001100111000111110;
    rom[14361] = 25'b0000000001100111001111110;
    rom[14362] = 25'b0000000001100111010111101;
    rom[14363] = 25'b0000000001100111011111101;
    rom[14364] = 25'b0000000001100111100111101;
    rom[14365] = 25'b0000000001100111101111101;
    rom[14366] = 25'b0000000001100111110111100;
    rom[14367] = 25'b0000000001100111111111100;
    rom[14368] = 25'b0000000001101000000111011;
    rom[14369] = 25'b0000000001101000001111011;
    rom[14370] = 25'b0000000001101000010111010;
    rom[14371] = 25'b0000000001101000011111010;
    rom[14372] = 25'b0000000001101000100111001;
    rom[14373] = 25'b0000000001101000101111001;
    rom[14374] = 25'b0000000001101000110111000;
    rom[14375] = 25'b0000000001101000111110111;
    rom[14376] = 25'b0000000001101001000110110;
    rom[14377] = 25'b0000000001101001001110110;
    rom[14378] = 25'b0000000001101001010110101;
    rom[14379] = 25'b0000000001101001011110100;
    rom[14380] = 25'b0000000001101001100110011;
    rom[14381] = 25'b0000000001101001101110010;
    rom[14382] = 25'b0000000001101001110110001;
    rom[14383] = 25'b0000000001101001111110000;
    rom[14384] = 25'b0000000001101010000101111;
    rom[14385] = 25'b0000000001101010001101110;
    rom[14386] = 25'b0000000001101010010101101;
    rom[14387] = 25'b0000000001101010011101100;
    rom[14388] = 25'b0000000001101010100101010;
    rom[14389] = 25'b0000000001101010101101001;
    rom[14390] = 25'b0000000001101010110101000;
    rom[14391] = 25'b0000000001101010111100111;
    rom[14392] = 25'b0000000001101011000100101;
    rom[14393] = 25'b0000000001101011001100011;
    rom[14394] = 25'b0000000001101011010100010;
    rom[14395] = 25'b0000000001101011011100001;
    rom[14396] = 25'b0000000001101011100011111;
    rom[14397] = 25'b0000000001101011101011110;
    rom[14398] = 25'b0000000001101011110011100;
    rom[14399] = 25'b0000000001101011111011010;
    rom[14400] = 25'b0000000001101100000011000;
    rom[14401] = 25'b0000000001101100001010110;
    rom[14402] = 25'b0000000001101100010010101;
    rom[14403] = 25'b0000000001101100011010011;
    rom[14404] = 25'b0000000001101100100010001;
    rom[14405] = 25'b0000000001101100101001111;
    rom[14406] = 25'b0000000001101100110001101;
    rom[14407] = 25'b0000000001101100111001011;
    rom[14408] = 25'b0000000001101101000001001;
    rom[14409] = 25'b0000000001101101001000111;
    rom[14410] = 25'b0000000001101101010000101;
    rom[14411] = 25'b0000000001101101011000011;
    rom[14412] = 25'b0000000001101101100000001;
    rom[14413] = 25'b0000000001101101100111111;
    rom[14414] = 25'b0000000001101101101111100;
    rom[14415] = 25'b0000000001101101110111010;
    rom[14416] = 25'b0000000001101101111110111;
    rom[14417] = 25'b0000000001101110000110101;
    rom[14418] = 25'b0000000001101110001110010;
    rom[14419] = 25'b0000000001101110010110000;
    rom[14420] = 25'b0000000001101110011101101;
    rom[14421] = 25'b0000000001101110100101011;
    rom[14422] = 25'b0000000001101110101101000;
    rom[14423] = 25'b0000000001101110110100101;
    rom[14424] = 25'b0000000001101110111100011;
    rom[14425] = 25'b0000000001101111000100000;
    rom[14426] = 25'b0000000001101111001011100;
    rom[14427] = 25'b0000000001101111010011010;
    rom[14428] = 25'b0000000001101111011010111;
    rom[14429] = 25'b0000000001101111100010100;
    rom[14430] = 25'b0000000001101111101010001;
    rom[14431] = 25'b0000000001101111110001110;
    rom[14432] = 25'b0000000001101111111001011;
    rom[14433] = 25'b0000000001110000000001000;
    rom[14434] = 25'b0000000001110000001000100;
    rom[14435] = 25'b0000000001110000010000010;
    rom[14436] = 25'b0000000001110000010111110;
    rom[14437] = 25'b0000000001110000011111011;
    rom[14438] = 25'b0000000001110000100110111;
    rom[14439] = 25'b0000000001110000101110100;
    rom[14440] = 25'b0000000001110000110110000;
    rom[14441] = 25'b0000000001110000111101101;
    rom[14442] = 25'b0000000001110001000101001;
    rom[14443] = 25'b0000000001110001001100110;
    rom[14444] = 25'b0000000001110001010100010;
    rom[14445] = 25'b0000000001110001011011110;
    rom[14446] = 25'b0000000001110001100011011;
    rom[14447] = 25'b0000000001110001101010111;
    rom[14448] = 25'b0000000001110001110010011;
    rom[14449] = 25'b0000000001110001111001111;
    rom[14450] = 25'b0000000001110010000001011;
    rom[14451] = 25'b0000000001110010001000111;
    rom[14452] = 25'b0000000001110010010000011;
    rom[14453] = 25'b0000000001110010010111111;
    rom[14454] = 25'b0000000001110010011111011;
    rom[14455] = 25'b0000000001110010100110111;
    rom[14456] = 25'b0000000001110010101110010;
    rom[14457] = 25'b0000000001110010110101110;
    rom[14458] = 25'b0000000001110010111101010;
    rom[14459] = 25'b0000000001110011000100110;
    rom[14460] = 25'b0000000001110011001100001;
    rom[14461] = 25'b0000000001110011010011101;
    rom[14462] = 25'b0000000001110011011011000;
    rom[14463] = 25'b0000000001110011100010011;
    rom[14464] = 25'b0000000001110011101001111;
    rom[14465] = 25'b0000000001110011110001010;
    rom[14466] = 25'b0000000001110011111000101;
    rom[14467] = 25'b0000000001110100000000001;
    rom[14468] = 25'b0000000001110100000111100;
    rom[14469] = 25'b0000000001110100001110111;
    rom[14470] = 25'b0000000001110100010110010;
    rom[14471] = 25'b0000000001110100011101101;
    rom[14472] = 25'b0000000001110100100101000;
    rom[14473] = 25'b0000000001110100101100011;
    rom[14474] = 25'b0000000001110100110011110;
    rom[14475] = 25'b0000000001110100111011001;
    rom[14476] = 25'b0000000001110101000010011;
    rom[14477] = 25'b0000000001110101001001110;
    rom[14478] = 25'b0000000001110101010001001;
    rom[14479] = 25'b0000000001110101011000100;
    rom[14480] = 25'b0000000001110101011111110;
    rom[14481] = 25'b0000000001110101100111001;
    rom[14482] = 25'b0000000001110101101110011;
    rom[14483] = 25'b0000000001110101110101101;
    rom[14484] = 25'b0000000001110101111101000;
    rom[14485] = 25'b0000000001110110000100010;
    rom[14486] = 25'b0000000001110110001011100;
    rom[14487] = 25'b0000000001110110010010111;
    rom[14488] = 25'b0000000001110110011010001;
    rom[14489] = 25'b0000000001110110100001011;
    rom[14490] = 25'b0000000001110110101000101;
    rom[14491] = 25'b0000000001110110101111111;
    rom[14492] = 25'b0000000001110110110111001;
    rom[14493] = 25'b0000000001110110111110011;
    rom[14494] = 25'b0000000001110111000101101;
    rom[14495] = 25'b0000000001110111001100111;
    rom[14496] = 25'b0000000001110111010100001;
    rom[14497] = 25'b0000000001110111011011010;
    rom[14498] = 25'b0000000001110111100010100;
    rom[14499] = 25'b0000000001110111101001101;
    rom[14500] = 25'b0000000001110111110000111;
    rom[14501] = 25'b0000000001110111111000000;
    rom[14502] = 25'b0000000001110111111111010;
    rom[14503] = 25'b0000000001111000000110011;
    rom[14504] = 25'b0000000001111000001101101;
    rom[14505] = 25'b0000000001111000010100110;
    rom[14506] = 25'b0000000001111000011011111;
    rom[14507] = 25'b0000000001111000100011001;
    rom[14508] = 25'b0000000001111000101010010;
    rom[14509] = 25'b0000000001111000110001010;
    rom[14510] = 25'b0000000001111000111000100;
    rom[14511] = 25'b0000000001111000111111101;
    rom[14512] = 25'b0000000001111001000110101;
    rom[14513] = 25'b0000000001111001001101110;
    rom[14514] = 25'b0000000001111001010100111;
    rom[14515] = 25'b0000000001111001011100000;
    rom[14516] = 25'b0000000001111001100011001;
    rom[14517] = 25'b0000000001111001101010001;
    rom[14518] = 25'b0000000001111001110001010;
    rom[14519] = 25'b0000000001111001111000010;
    rom[14520] = 25'b0000000001111001111111011;
    rom[14521] = 25'b0000000001111010000110011;
    rom[14522] = 25'b0000000001111010001101100;
    rom[14523] = 25'b0000000001111010010100100;
    rom[14524] = 25'b0000000001111010011011100;
    rom[14525] = 25'b0000000001111010100010101;
    rom[14526] = 25'b0000000001111010101001101;
    rom[14527] = 25'b0000000001111010110000101;
    rom[14528] = 25'b0000000001111010110111101;
    rom[14529] = 25'b0000000001111010111110101;
    rom[14530] = 25'b0000000001111011000101101;
    rom[14531] = 25'b0000000001111011001100100;
    rom[14532] = 25'b0000000001111011010011100;
    rom[14533] = 25'b0000000001111011011010100;
    rom[14534] = 25'b0000000001111011100001011;
    rom[14535] = 25'b0000000001111011101000011;
    rom[14536] = 25'b0000000001111011101111011;
    rom[14537] = 25'b0000000001111011110110010;
    rom[14538] = 25'b0000000001111011111101010;
    rom[14539] = 25'b0000000001111100000100001;
    rom[14540] = 25'b0000000001111100001011001;
    rom[14541] = 25'b0000000001111100010010000;
    rom[14542] = 25'b0000000001111100011000111;
    rom[14543] = 25'b0000000001111100011111110;
    rom[14544] = 25'b0000000001111100100110101;
    rom[14545] = 25'b0000000001111100101101100;
    rom[14546] = 25'b0000000001111100110100100;
    rom[14547] = 25'b0000000001111100111011010;
    rom[14548] = 25'b0000000001111101000010001;
    rom[14549] = 25'b0000000001111101001001000;
    rom[14550] = 25'b0000000001111101001111110;
    rom[14551] = 25'b0000000001111101010110110;
    rom[14552] = 25'b0000000001111101011101100;
    rom[14553] = 25'b0000000001111101100100011;
    rom[14554] = 25'b0000000001111101101011001;
    rom[14555] = 25'b0000000001111101110010000;
    rom[14556] = 25'b0000000001111101111000110;
    rom[14557] = 25'b0000000001111101111111100;
    rom[14558] = 25'b0000000001111110000110011;
    rom[14559] = 25'b0000000001111110001101001;
    rom[14560] = 25'b0000000001111110010011111;
    rom[14561] = 25'b0000000001111110011010101;
    rom[14562] = 25'b0000000001111110100001011;
    rom[14563] = 25'b0000000001111110101000001;
    rom[14564] = 25'b0000000001111110101110111;
    rom[14565] = 25'b0000000001111110110101101;
    rom[14566] = 25'b0000000001111110111100011;
    rom[14567] = 25'b0000000001111111000011000;
    rom[14568] = 25'b0000000001111111001001110;
    rom[14569] = 25'b0000000001111111010000100;
    rom[14570] = 25'b0000000001111111010111010;
    rom[14571] = 25'b0000000001111111011101111;
    rom[14572] = 25'b0000000001111111100100101;
    rom[14573] = 25'b0000000001111111101011010;
    rom[14574] = 25'b0000000001111111110001111;
    rom[14575] = 25'b0000000001111111111000101;
    rom[14576] = 25'b0000000001111111111111010;
    rom[14577] = 25'b0000000010000000000101111;
    rom[14578] = 25'b0000000010000000001100100;
    rom[14579] = 25'b0000000010000000010011001;
    rom[14580] = 25'b0000000010000000011001110;
    rom[14581] = 25'b0000000010000000100000011;
    rom[14582] = 25'b0000000010000000100111000;
    rom[14583] = 25'b0000000010000000101101100;
    rom[14584] = 25'b0000000010000000110100001;
    rom[14585] = 25'b0000000010000000111010101;
    rom[14586] = 25'b0000000010000001000001010;
    rom[14587] = 25'b0000000010000001000111111;
    rom[14588] = 25'b0000000010000001001110011;
    rom[14589] = 25'b0000000010000001010100111;
    rom[14590] = 25'b0000000010000001011011100;
    rom[14591] = 25'b0000000010000001100010000;
    rom[14592] = 25'b0000000010000001101000100;
    rom[14593] = 25'b0000000010000001101111001;
    rom[14594] = 25'b0000000010000001110101101;
    rom[14595] = 25'b0000000010000001111100000;
    rom[14596] = 25'b0000000010000010000010101;
    rom[14597] = 25'b0000000010000010001001000;
    rom[14598] = 25'b0000000010000010001111101;
    rom[14599] = 25'b0000000010000010010110000;
    rom[14600] = 25'b0000000010000010011100100;
    rom[14601] = 25'b0000000010000010100010111;
    rom[14602] = 25'b0000000010000010101001011;
    rom[14603] = 25'b0000000010000010101111110;
    rom[14604] = 25'b0000000010000010110110010;
    rom[14605] = 25'b0000000010000010111100101;
    rom[14606] = 25'b0000000010000011000011001;
    rom[14607] = 25'b0000000010000011001001100;
    rom[14608] = 25'b0000000010000011001111111;
    rom[14609] = 25'b0000000010000011010110010;
    rom[14610] = 25'b0000000010000011011100101;
    rom[14611] = 25'b0000000010000011100011000;
    rom[14612] = 25'b0000000010000011101001011;
    rom[14613] = 25'b0000000010000011101111110;
    rom[14614] = 25'b0000000010000011110110001;
    rom[14615] = 25'b0000000010000011111100100;
    rom[14616] = 25'b0000000010000100000010110;
    rom[14617] = 25'b0000000010000100001001001;
    rom[14618] = 25'b0000000010000100001111011;
    rom[14619] = 25'b0000000010000100010101101;
    rom[14620] = 25'b0000000010000100011100000;
    rom[14621] = 25'b0000000010000100100010010;
    rom[14622] = 25'b0000000010000100101000101;
    rom[14623] = 25'b0000000010000100101110111;
    rom[14624] = 25'b0000000010000100110101001;
    rom[14625] = 25'b0000000010000100111011011;
    rom[14626] = 25'b0000000010000101000001101;
    rom[14627] = 25'b0000000010000101000111111;
    rom[14628] = 25'b0000000010000101001110001;
    rom[14629] = 25'b0000000010000101010100011;
    rom[14630] = 25'b0000000010000101011010100;
    rom[14631] = 25'b0000000010000101100000110;
    rom[14632] = 25'b0000000010000101100110111;
    rom[14633] = 25'b0000000010000101101101001;
    rom[14634] = 25'b0000000010000101110011011;
    rom[14635] = 25'b0000000010000101111001100;
    rom[14636] = 25'b0000000010000101111111101;
    rom[14637] = 25'b0000000010000110000101111;
    rom[14638] = 25'b0000000010000110001100000;
    rom[14639] = 25'b0000000010000110010010001;
    rom[14640] = 25'b0000000010000110011000010;
    rom[14641] = 25'b0000000010000110011110011;
    rom[14642] = 25'b0000000010000110100100100;
    rom[14643] = 25'b0000000010000110101010100;
    rom[14644] = 25'b0000000010000110110000110;
    rom[14645] = 25'b0000000010000110110110110;
    rom[14646] = 25'b0000000010000110111100111;
    rom[14647] = 25'b0000000010000111000010111;
    rom[14648] = 25'b0000000010000111001001000;
    rom[14649] = 25'b0000000010000111001111000;
    rom[14650] = 25'b0000000010000111010101000;
    rom[14651] = 25'b0000000010000111011011001;
    rom[14652] = 25'b0000000010000111100001001;
    rom[14653] = 25'b0000000010000111100111001;
    rom[14654] = 25'b0000000010000111101101001;
    rom[14655] = 25'b0000000010000111110011001;
    rom[14656] = 25'b0000000010000111111001001;
    rom[14657] = 25'b0000000010000111111111001;
    rom[14658] = 25'b0000000010001000000101001;
    rom[14659] = 25'b0000000010001000001011001;
    rom[14660] = 25'b0000000010001000010001001;
    rom[14661] = 25'b0000000010001000010111000;
    rom[14662] = 25'b0000000010001000011100111;
    rom[14663] = 25'b0000000010001000100010111;
    rom[14664] = 25'b0000000010001000101000110;
    rom[14665] = 25'b0000000010001000101110101;
    rom[14666] = 25'b0000000010001000110100100;
    rom[14667] = 25'b0000000010001000111010100;
    rom[14668] = 25'b0000000010001001000000011;
    rom[14669] = 25'b0000000010001001000110010;
    rom[14670] = 25'b0000000010001001001100001;
    rom[14671] = 25'b0000000010001001010010000;
    rom[14672] = 25'b0000000010001001010111111;
    rom[14673] = 25'b0000000010001001011101101;
    rom[14674] = 25'b0000000010001001100011100;
    rom[14675] = 25'b0000000010001001101001011;
    rom[14676] = 25'b0000000010001001101111001;
    rom[14677] = 25'b0000000010001001110100111;
    rom[14678] = 25'b0000000010001001111010110;
    rom[14679] = 25'b0000000010001010000000100;
    rom[14680] = 25'b0000000010001010000110010;
    rom[14681] = 25'b0000000010001010001100000;
    rom[14682] = 25'b0000000010001010010001111;
    rom[14683] = 25'b0000000010001010010111100;
    rom[14684] = 25'b0000000010001010011101011;
    rom[14685] = 25'b0000000010001010100011000;
    rom[14686] = 25'b0000000010001010101000110;
    rom[14687] = 25'b0000000010001010101110011;
    rom[14688] = 25'b0000000010001010110100010;
    rom[14689] = 25'b0000000010001010111001111;
    rom[14690] = 25'b0000000010001010111111100;
    rom[14691] = 25'b0000000010001011000101010;
    rom[14692] = 25'b0000000010001011001010111;
    rom[14693] = 25'b0000000010001011010000100;
    rom[14694] = 25'b0000000010001011010110010;
    rom[14695] = 25'b0000000010001011011011111;
    rom[14696] = 25'b0000000010001011100001100;
    rom[14697] = 25'b0000000010001011100111001;
    rom[14698] = 25'b0000000010001011101100110;
    rom[14699] = 25'b0000000010001011110010011;
    rom[14700] = 25'b0000000010001011110111111;
    rom[14701] = 25'b0000000010001011111101100;
    rom[14702] = 25'b0000000010001100000011000;
    rom[14703] = 25'b0000000010001100001000101;
    rom[14704] = 25'b0000000010001100001110001;
    rom[14705] = 25'b0000000010001100010011110;
    rom[14706] = 25'b0000000010001100011001010;
    rom[14707] = 25'b0000000010001100011110110;
    rom[14708] = 25'b0000000010001100100100010;
    rom[14709] = 25'b0000000010001100101001110;
    rom[14710] = 25'b0000000010001100101111010;
    rom[14711] = 25'b0000000010001100110100110;
    rom[14712] = 25'b0000000010001100111010010;
    rom[14713] = 25'b0000000010001100111111110;
    rom[14714] = 25'b0000000010001101000101010;
    rom[14715] = 25'b0000000010001101001010101;
    rom[14716] = 25'b0000000010001101010000001;
    rom[14717] = 25'b0000000010001101010101100;
    rom[14718] = 25'b0000000010001101011010111;
    rom[14719] = 25'b0000000010001101100000011;
    rom[14720] = 25'b0000000010001101100101110;
    rom[14721] = 25'b0000000010001101101011001;
    rom[14722] = 25'b0000000010001101110000101;
    rom[14723] = 25'b0000000010001101110101111;
    rom[14724] = 25'b0000000010001101111011011;
    rom[14725] = 25'b0000000010001110000000101;
    rom[14726] = 25'b0000000010001110000110000;
    rom[14727] = 25'b0000000010001110001011010;
    rom[14728] = 25'b0000000010001110010000101;
    rom[14729] = 25'b0000000010001110010101111;
    rom[14730] = 25'b0000000010001110011011010;
    rom[14731] = 25'b0000000010001110100000101;
    rom[14732] = 25'b0000000010001110100101110;
    rom[14733] = 25'b0000000010001110101011001;
    rom[14734] = 25'b0000000010001110110000011;
    rom[14735] = 25'b0000000010001110110101101;
    rom[14736] = 25'b0000000010001110111010111;
    rom[14737] = 25'b0000000010001111000000001;
    rom[14738] = 25'b0000000010001111000101011;
    rom[14739] = 25'b0000000010001111001010101;
    rom[14740] = 25'b0000000010001111001111110;
    rom[14741] = 25'b0000000010001111010101000;
    rom[14742] = 25'b0000000010001111011010010;
    rom[14743] = 25'b0000000010001111011111011;
    rom[14744] = 25'b0000000010001111100100100;
    rom[14745] = 25'b0000000010001111101001110;
    rom[14746] = 25'b0000000010001111101110111;
    rom[14747] = 25'b0000000010001111110100000;
    rom[14748] = 25'b0000000010001111111001001;
    rom[14749] = 25'b0000000010001111111110001;
    rom[14750] = 25'b0000000010010000000011010;
    rom[14751] = 25'b0000000010010000001000011;
    rom[14752] = 25'b0000000010010000001101100;
    rom[14753] = 25'b0000000010010000010010101;
    rom[14754] = 25'b0000000010010000010111101;
    rom[14755] = 25'b0000000010010000011100110;
    rom[14756] = 25'b0000000010010000100001110;
    rom[14757] = 25'b0000000010010000100110110;
    rom[14758] = 25'b0000000010010000101011111;
    rom[14759] = 25'b0000000010010000110000110;
    rom[14760] = 25'b0000000010010000110101111;
    rom[14761] = 25'b0000000010010000111010111;
    rom[14762] = 25'b0000000010010000111111110;
    rom[14763] = 25'b0000000010010001000100110;
    rom[14764] = 25'b0000000010010001001001110;
    rom[14765] = 25'b0000000010010001001110110;
    rom[14766] = 25'b0000000010010001010011101;
    rom[14767] = 25'b0000000010010001011000100;
    rom[14768] = 25'b0000000010010001011101100;
    rom[14769] = 25'b0000000010010001100010100;
    rom[14770] = 25'b0000000010010001100111010;
    rom[14771] = 25'b0000000010010001101100010;
    rom[14772] = 25'b0000000010010001110001001;
    rom[14773] = 25'b0000000010010001110110000;
    rom[14774] = 25'b0000000010010001111010111;
    rom[14775] = 25'b0000000010010001111111101;
    rom[14776] = 25'b0000000010010010000100100;
    rom[14777] = 25'b0000000010010010001001011;
    rom[14778] = 25'b0000000010010010001110001;
    rom[14779] = 25'b0000000010010010010011000;
    rom[14780] = 25'b0000000010010010010111110;
    rom[14781] = 25'b0000000010010010011100101;
    rom[14782] = 25'b0000000010010010100001011;
    rom[14783] = 25'b0000000010010010100110001;
    rom[14784] = 25'b0000000010010010101010111;
    rom[14785] = 25'b0000000010010010101111101;
    rom[14786] = 25'b0000000010010010110100011;
    rom[14787] = 25'b0000000010010010111001001;
    rom[14788] = 25'b0000000010010010111101111;
    rom[14789] = 25'b0000000010010011000010100;
    rom[14790] = 25'b0000000010010011000111010;
    rom[14791] = 25'b0000000010010011001011111;
    rom[14792] = 25'b0000000010010011010000100;
    rom[14793] = 25'b0000000010010011010101010;
    rom[14794] = 25'b0000000010010011011001111;
    rom[14795] = 25'b0000000010010011011110101;
    rom[14796] = 25'b0000000010010011100011010;
    rom[14797] = 25'b0000000010010011100111110;
    rom[14798] = 25'b0000000010010011101100011;
    rom[14799] = 25'b0000000010010011110001000;
    rom[14800] = 25'b0000000010010011110101101;
    rom[14801] = 25'b0000000010010011111010010;
    rom[14802] = 25'b0000000010010011111110110;
    rom[14803] = 25'b0000000010010100000011011;
    rom[14804] = 25'b0000000010010100000111111;
    rom[14805] = 25'b0000000010010100001100011;
    rom[14806] = 25'b0000000010010100010000111;
    rom[14807] = 25'b0000000010010100010101100;
    rom[14808] = 25'b0000000010010100011010000;
    rom[14809] = 25'b0000000010010100011110100;
    rom[14810] = 25'b0000000010010100100010111;
    rom[14811] = 25'b0000000010010100100111011;
    rom[14812] = 25'b0000000010010100101011111;
    rom[14813] = 25'b0000000010010100110000010;
    rom[14814] = 25'b0000000010010100110100110;
    rom[14815] = 25'b0000000010010100111001001;
    rom[14816] = 25'b0000000010010100111101101;
    rom[14817] = 25'b0000000010010101000010000;
    rom[14818] = 25'b0000000010010101000110011;
    rom[14819] = 25'b0000000010010101001010110;
    rom[14820] = 25'b0000000010010101001111010;
    rom[14821] = 25'b0000000010010101010011101;
    rom[14822] = 25'b0000000010010101010111111;
    rom[14823] = 25'b0000000010010101011100010;
    rom[14824] = 25'b0000000010010101100000100;
    rom[14825] = 25'b0000000010010101100100111;
    rom[14826] = 25'b0000000010010101101001001;
    rom[14827] = 25'b0000000010010101101101100;
    rom[14828] = 25'b0000000010010101110001110;
    rom[14829] = 25'b0000000010010101110110000;
    rom[14830] = 25'b0000000010010101111010011;
    rom[14831] = 25'b0000000010010101111110100;
    rom[14832] = 25'b0000000010010110000010111;
    rom[14833] = 25'b0000000010010110000111000;
    rom[14834] = 25'b0000000010010110001011010;
    rom[14835] = 25'b0000000010010110001111100;
    rom[14836] = 25'b0000000010010110010011101;
    rom[14837] = 25'b0000000010010110010111111;
    rom[14838] = 25'b0000000010010110011100000;
    rom[14839] = 25'b0000000010010110100000001;
    rom[14840] = 25'b0000000010010110100100011;
    rom[14841] = 25'b0000000010010110101000100;
    rom[14842] = 25'b0000000010010110101100101;
    rom[14843] = 25'b0000000010010110110000110;
    rom[14844] = 25'b0000000010010110110100111;
    rom[14845] = 25'b0000000010010110111001000;
    rom[14846] = 25'b0000000010010110111101000;
    rom[14847] = 25'b0000000010010111000001001;
    rom[14848] = 25'b0000000010010111000101001;
    rom[14849] = 25'b0000000010010111001001010;
    rom[14850] = 25'b0000000010010111001101010;
    rom[14851] = 25'b0000000010010111010001010;
    rom[14852] = 25'b0000000010010111010101010;
    rom[14853] = 25'b0000000010010111011001010;
    rom[14854] = 25'b0000000010010111011101011;
    rom[14855] = 25'b0000000010010111100001011;
    rom[14856] = 25'b0000000010010111100101010;
    rom[14857] = 25'b0000000010010111101001010;
    rom[14858] = 25'b0000000010010111101101010;
    rom[14859] = 25'b0000000010010111110001001;
    rom[14860] = 25'b0000000010010111110101000;
    rom[14861] = 25'b0000000010010111111001000;
    rom[14862] = 25'b0000000010010111111100111;
    rom[14863] = 25'b0000000010011000000000110;
    rom[14864] = 25'b0000000010011000000100101;
    rom[14865] = 25'b0000000010011000001000100;
    rom[14866] = 25'b0000000010011000001100011;
    rom[14867] = 25'b0000000010011000010000010;
    rom[14868] = 25'b0000000010011000010100000;
    rom[14869] = 25'b0000000010011000010111111;
    rom[14870] = 25'b0000000010011000011011110;
    rom[14871] = 25'b0000000010011000011111100;
    rom[14872] = 25'b0000000010011000100011010;
    rom[14873] = 25'b0000000010011000100111001;
    rom[14874] = 25'b0000000010011000101010111;
    rom[14875] = 25'b0000000010011000101110101;
    rom[14876] = 25'b0000000010011000110010011;
    rom[14877] = 25'b0000000010011000110110001;
    rom[14878] = 25'b0000000010011000111001110;
    rom[14879] = 25'b0000000010011000111101100;
    rom[14880] = 25'b0000000010011001000001010;
    rom[14881] = 25'b0000000010011001000100111;
    rom[14882] = 25'b0000000010011001001000101;
    rom[14883] = 25'b0000000010011001001100010;
    rom[14884] = 25'b0000000010011001001111111;
    rom[14885] = 25'b0000000010011001010011100;
    rom[14886] = 25'b0000000010011001010111010;
    rom[14887] = 25'b0000000010011001011010110;
    rom[14888] = 25'b0000000010011001011110011;
    rom[14889] = 25'b0000000010011001100001111;
    rom[14890] = 25'b0000000010011001100101101;
    rom[14891] = 25'b0000000010011001101001001;
    rom[14892] = 25'b0000000010011001101100101;
    rom[14893] = 25'b0000000010011001110000010;
    rom[14894] = 25'b0000000010011001110011110;
    rom[14895] = 25'b0000000010011001110111011;
    rom[14896] = 25'b0000000010011001111010110;
    rom[14897] = 25'b0000000010011001111110011;
    rom[14898] = 25'b0000000010011010000001110;
    rom[14899] = 25'b0000000010011010000101010;
    rom[14900] = 25'b0000000010011010001000110;
    rom[14901] = 25'b0000000010011010001100001;
    rom[14902] = 25'b0000000010011010001111101;
    rom[14903] = 25'b0000000010011010010011000;
    rom[14904] = 25'b0000000010011010010110011;
    rom[14905] = 25'b0000000010011010011001111;
    rom[14906] = 25'b0000000010011010011101010;
    rom[14907] = 25'b0000000010011010100000101;
    rom[14908] = 25'b0000000010011010100100000;
    rom[14909] = 25'b0000000010011010100111011;
    rom[14910] = 25'b0000000010011010101010101;
    rom[14911] = 25'b0000000010011010101110000;
    rom[14912] = 25'b0000000010011010110001010;
    rom[14913] = 25'b0000000010011010110100101;
    rom[14914] = 25'b0000000010011010111000000;
    rom[14915] = 25'b0000000010011010111011010;
    rom[14916] = 25'b0000000010011010111110100;
    rom[14917] = 25'b0000000010011011000001110;
    rom[14918] = 25'b0000000010011011000101000;
    rom[14919] = 25'b0000000010011011001000010;
    rom[14920] = 25'b0000000010011011001011100;
    rom[14921] = 25'b0000000010011011001110101;
    rom[14922] = 25'b0000000010011011010001111;
    rom[14923] = 25'b0000000010011011010101001;
    rom[14924] = 25'b0000000010011011011000010;
    rom[14925] = 25'b0000000010011011011011011;
    rom[14926] = 25'b0000000010011011011110100;
    rom[14927] = 25'b0000000010011011100001101;
    rom[14928] = 25'b0000000010011011100100110;
    rom[14929] = 25'b0000000010011011101000000;
    rom[14930] = 25'b0000000010011011101011000;
    rom[14931] = 25'b0000000010011011101110001;
    rom[14932] = 25'b0000000010011011110001010;
    rom[14933] = 25'b0000000010011011110100010;
    rom[14934] = 25'b0000000010011011110111010;
    rom[14935] = 25'b0000000010011011111010011;
    rom[14936] = 25'b0000000010011011111101011;
    rom[14937] = 25'b0000000010011100000000011;
    rom[14938] = 25'b0000000010011100000011011;
    rom[14939] = 25'b0000000010011100000110011;
    rom[14940] = 25'b0000000010011100001001011;
    rom[14941] = 25'b0000000010011100001100010;
    rom[14942] = 25'b0000000010011100001111010;
    rom[14943] = 25'b0000000010011100010010010;
    rom[14944] = 25'b0000000010011100010101001;
    rom[14945] = 25'b0000000010011100011000000;
    rom[14946] = 25'b0000000010011100011010111;
    rom[14947] = 25'b0000000010011100011101111;
    rom[14948] = 25'b0000000010011100100000110;
    rom[14949] = 25'b0000000010011100100011101;
    rom[14950] = 25'b0000000010011100100110011;
    rom[14951] = 25'b0000000010011100101001011;
    rom[14952] = 25'b0000000010011100101100001;
    rom[14953] = 25'b0000000010011100101110111;
    rom[14954] = 25'b0000000010011100110001110;
    rom[14955] = 25'b0000000010011100110100100;
    rom[14956] = 25'b0000000010011100110111011;
    rom[14957] = 25'b0000000010011100111010001;
    rom[14958] = 25'b0000000010011100111100111;
    rom[14959] = 25'b0000000010011100111111100;
    rom[14960] = 25'b0000000010011101000010011;
    rom[14961] = 25'b0000000010011101000101000;
    rom[14962] = 25'b0000000010011101000111110;
    rom[14963] = 25'b0000000010011101001010100;
    rom[14964] = 25'b0000000010011101001101001;
    rom[14965] = 25'b0000000010011101001111110;
    rom[14966] = 25'b0000000010011101010010011;
    rom[14967] = 25'b0000000010011101010101000;
    rom[14968] = 25'b0000000010011101010111110;
    rom[14969] = 25'b0000000010011101011010011;
    rom[14970] = 25'b0000000010011101011100111;
    rom[14971] = 25'b0000000010011101011111100;
    rom[14972] = 25'b0000000010011101100010001;
    rom[14973] = 25'b0000000010011101100100101;
    rom[14974] = 25'b0000000010011101100111010;
    rom[14975] = 25'b0000000010011101101001110;
    rom[14976] = 25'b0000000010011101101100010;
    rom[14977] = 25'b0000000010011101101110110;
    rom[14978] = 25'b0000000010011101110001011;
    rom[14979] = 25'b0000000010011101110011110;
    rom[14980] = 25'b0000000010011101110110010;
    rom[14981] = 25'b0000000010011101111000110;
    rom[14982] = 25'b0000000010011101111011001;
    rom[14983] = 25'b0000000010011101111101100;
    rom[14984] = 25'b0000000010011110000000000;
    rom[14985] = 25'b0000000010011110000010011;
    rom[14986] = 25'b0000000010011110000100111;
    rom[14987] = 25'b0000000010011110000111010;
    rom[14988] = 25'b0000000010011110001001101;
    rom[14989] = 25'b0000000010011110001011111;
    rom[14990] = 25'b0000000010011110001110010;
    rom[14991] = 25'b0000000010011110010000101;
    rom[14992] = 25'b0000000010011110010010111;
    rom[14993] = 25'b0000000010011110010101010;
    rom[14994] = 25'b0000000010011110010111101;
    rom[14995] = 25'b0000000010011110011001111;
    rom[14996] = 25'b0000000010011110011100001;
    rom[14997] = 25'b0000000010011110011110011;
    rom[14998] = 25'b0000000010011110100000101;
    rom[14999] = 25'b0000000010011110100010110;
    rom[15000] = 25'b0000000010011110100101000;
    rom[15001] = 25'b0000000010011110100111010;
    rom[15002] = 25'b0000000010011110101001100;
    rom[15003] = 25'b0000000010011110101011101;
    rom[15004] = 25'b0000000010011110101101111;
    rom[15005] = 25'b0000000010011110110000000;
    rom[15006] = 25'b0000000010011110110010001;
    rom[15007] = 25'b0000000010011110110100010;
    rom[15008] = 25'b0000000010011110110110011;
    rom[15009] = 25'b0000000010011110111000100;
    rom[15010] = 25'b0000000010011110111010100;
    rom[15011] = 25'b0000000010011110111100101;
    rom[15012] = 25'b0000000010011110111110101;
    rom[15013] = 25'b0000000010011111000000110;
    rom[15014] = 25'b0000000010011111000010110;
    rom[15015] = 25'b0000000010011111000100110;
    rom[15016] = 25'b0000000010011111000110110;
    rom[15017] = 25'b0000000010011111001000111;
    rom[15018] = 25'b0000000010011111001010110;
    rom[15019] = 25'b0000000010011111001100110;
    rom[15020] = 25'b0000000010011111001110110;
    rom[15021] = 25'b0000000010011111010000101;
    rom[15022] = 25'b0000000010011111010010100;
    rom[15023] = 25'b0000000010011111010100100;
    rom[15024] = 25'b0000000010011111010110011;
    rom[15025] = 25'b0000000010011111011000011;
    rom[15026] = 25'b0000000010011111011010010;
    rom[15027] = 25'b0000000010011111011100000;
    rom[15028] = 25'b0000000010011111011101111;
    rom[15029] = 25'b0000000010011111011111110;
    rom[15030] = 25'b0000000010011111100001101;
    rom[15031] = 25'b0000000010011111100011011;
    rom[15032] = 25'b0000000010011111100101001;
    rom[15033] = 25'b0000000010011111100110111;
    rom[15034] = 25'b0000000010011111101000101;
    rom[15035] = 25'b0000000010011111101010100;
    rom[15036] = 25'b0000000010011111101100010;
    rom[15037] = 25'b0000000010011111101101111;
    rom[15038] = 25'b0000000010011111101111101;
    rom[15039] = 25'b0000000010011111110001011;
    rom[15040] = 25'b0000000010011111110011000;
    rom[15041] = 25'b0000000010011111110100110;
    rom[15042] = 25'b0000000010011111110110011;
    rom[15043] = 25'b0000000010011111111000001;
    rom[15044] = 25'b0000000010011111111001101;
    rom[15045] = 25'b0000000010011111111011011;
    rom[15046] = 25'b0000000010011111111100111;
    rom[15047] = 25'b0000000010011111111110100;
    rom[15048] = 25'b0000000010100000000000001;
    rom[15049] = 25'b0000000010100000000001110;
    rom[15050] = 25'b0000000010100000000011001;
    rom[15051] = 25'b0000000010100000000100110;
    rom[15052] = 25'b0000000010100000000110010;
    rom[15053] = 25'b0000000010100000000111110;
    rom[15054] = 25'b0000000010100000001001011;
    rom[15055] = 25'b0000000010100000001010110;
    rom[15056] = 25'b0000000010100000001100010;
    rom[15057] = 25'b0000000010100000001101110;
    rom[15058] = 25'b0000000010100000001111001;
    rom[15059] = 25'b0000000010100000010000101;
    rom[15060] = 25'b0000000010100000010010000;
    rom[15061] = 25'b0000000010100000010011011;
    rom[15062] = 25'b0000000010100000010100111;
    rom[15063] = 25'b0000000010100000010110010;
    rom[15064] = 25'b0000000010100000010111100;
    rom[15065] = 25'b0000000010100000011001000;
    rom[15066] = 25'b0000000010100000011010010;
    rom[15067] = 25'b0000000010100000011011100;
    rom[15068] = 25'b0000000010100000011100111;
    rom[15069] = 25'b0000000010100000011110001;
    rom[15070] = 25'b0000000010100000011111100;
    rom[15071] = 25'b0000000010100000100000110;
    rom[15072] = 25'b0000000010100000100010000;
    rom[15073] = 25'b0000000010100000100011010;
    rom[15074] = 25'b0000000010100000100100100;
    rom[15075] = 25'b0000000010100000100101110;
    rom[15076] = 25'b0000000010100000100111000;
    rom[15077] = 25'b0000000010100000101000001;
    rom[15078] = 25'b0000000010100000101001010;
    rom[15079] = 25'b0000000010100000101010011;
    rom[15080] = 25'b0000000010100000101011101;
    rom[15081] = 25'b0000000010100000101100110;
    rom[15082] = 25'b0000000010100000101101111;
    rom[15083] = 25'b0000000010100000101111000;
    rom[15084] = 25'b0000000010100000110000000;
    rom[15085] = 25'b0000000010100000110001001;
    rom[15086] = 25'b0000000010100000110010001;
    rom[15087] = 25'b0000000010100000110011001;
    rom[15088] = 25'b0000000010100000110100010;
    rom[15089] = 25'b0000000010100000110101011;
    rom[15090] = 25'b0000000010100000110110010;
    rom[15091] = 25'b0000000010100000110111010;
    rom[15092] = 25'b0000000010100000111000011;
    rom[15093] = 25'b0000000010100000111001010;
    rom[15094] = 25'b0000000010100000111010010;
    rom[15095] = 25'b0000000010100000111011001;
    rom[15096] = 25'b0000000010100000111100000;
    rom[15097] = 25'b0000000010100000111101000;
    rom[15098] = 25'b0000000010100000111101111;
    rom[15099] = 25'b0000000010100000111110110;
    rom[15100] = 25'b0000000010100000111111101;
    rom[15101] = 25'b0000000010100001000000100;
    rom[15102] = 25'b0000000010100001000001010;
    rom[15103] = 25'b0000000010100001000010001;
    rom[15104] = 25'b0000000010100001000011000;
    rom[15105] = 25'b0000000010100001000011110;
    rom[15106] = 25'b0000000010100001000100100;
    rom[15107] = 25'b0000000010100001000101010;
    rom[15108] = 25'b0000000010100001000110000;
    rom[15109] = 25'b0000000010100001000110110;
    rom[15110] = 25'b0000000010100001000111100;
    rom[15111] = 25'b0000000010100001001000010;
    rom[15112] = 25'b0000000010100001001001000;
    rom[15113] = 25'b0000000010100001001001110;
    rom[15114] = 25'b0000000010100001001010011;
    rom[15115] = 25'b0000000010100001001011000;
    rom[15116] = 25'b0000000010100001001011101;
    rom[15117] = 25'b0000000010100001001100010;
    rom[15118] = 25'b0000000010100001001100111;
    rom[15119] = 25'b0000000010100001001101100;
    rom[15120] = 25'b0000000010100001001110001;
    rom[15121] = 25'b0000000010100001001110101;
    rom[15122] = 25'b0000000010100001001111010;
    rom[15123] = 25'b0000000010100001001111110;
    rom[15124] = 25'b0000000010100001010000011;
    rom[15125] = 25'b0000000010100001010000110;
    rom[15126] = 25'b0000000010100001010001011;
    rom[15127] = 25'b0000000010100001010001111;
    rom[15128] = 25'b0000000010100001010010010;
    rom[15129] = 25'b0000000010100001010010110;
    rom[15130] = 25'b0000000010100001010011010;
    rom[15131] = 25'b0000000010100001010011101;
    rom[15132] = 25'b0000000010100001010100000;
    rom[15133] = 25'b0000000010100001010100011;
    rom[15134] = 25'b0000000010100001010100110;
    rom[15135] = 25'b0000000010100001010101001;
    rom[15136] = 25'b0000000010100001010101100;
    rom[15137] = 25'b0000000010100001010101111;
    rom[15138] = 25'b0000000010100001010110010;
    rom[15139] = 25'b0000000010100001010110101;
    rom[15140] = 25'b0000000010100001010110111;
    rom[15141] = 25'b0000000010100001010111001;
    rom[15142] = 25'b0000000010100001010111011;
    rom[15143] = 25'b0000000010100001010111110;
    rom[15144] = 25'b0000000010100001011000000;
    rom[15145] = 25'b0000000010100001011000001;
    rom[15146] = 25'b0000000010100001011000011;
    rom[15147] = 25'b0000000010100001011000101;
    rom[15148] = 25'b0000000010100001011000111;
    rom[15149] = 25'b0000000010100001011000111;
    rom[15150] = 25'b0000000010100001011001001;
    rom[15151] = 25'b0000000010100001011001010;
    rom[15152] = 25'b0000000010100001011001011;
    rom[15153] = 25'b0000000010100001011001100;
    rom[15154] = 25'b0000000010100001011001101;
    rom[15155] = 25'b0000000010100001011001101;
    rom[15156] = 25'b0000000010100001011001110;
    rom[15157] = 25'b0000000010100001011001111;
    rom[15158] = 25'b0000000010100001011001111;
    rom[15159] = 25'b0000000010100001011010000;
    rom[15160] = 25'b0000000010100001011010000;
    rom[15161] = 25'b0000000010100001011010000;
    rom[15162] = 25'b0000000010100001011010000;
    rom[15163] = 25'b0000000010100001011001111;
    rom[15164] = 25'b0000000010100001011001111;
    rom[15165] = 25'b0000000010100001011001110;
    rom[15166] = 25'b0000000010100001011001110;
    rom[15167] = 25'b0000000010100001011001101;
    rom[15168] = 25'b0000000010100001011001101;
    rom[15169] = 25'b0000000010100001011001011;
    rom[15170] = 25'b0000000010100001011001010;
    rom[15171] = 25'b0000000010100001011001010;
    rom[15172] = 25'b0000000010100001011001000;
    rom[15173] = 25'b0000000010100001011000111;
    rom[15174] = 25'b0000000010100001011000101;
    rom[15175] = 25'b0000000010100001011000100;
    rom[15176] = 25'b0000000010100001011000010;
    rom[15177] = 25'b0000000010100001011000000;
    rom[15178] = 25'b0000000010100001010111110;
    rom[15179] = 25'b0000000010100001010111100;
    rom[15180] = 25'b0000000010100001010111010;
    rom[15181] = 25'b0000000010100001010111000;
    rom[15182] = 25'b0000000010100001010110101;
    rom[15183] = 25'b0000000010100001010110010;
    rom[15184] = 25'b0000000010100001010101111;
    rom[15185] = 25'b0000000010100001010101101;
    rom[15186] = 25'b0000000010100001010101010;
    rom[15187] = 25'b0000000010100001010100111;
    rom[15188] = 25'b0000000010100001010100011;
    rom[15189] = 25'b0000000010100001010100000;
    rom[15190] = 25'b0000000010100001010011101;
    rom[15191] = 25'b0000000010100001010011010;
    rom[15192] = 25'b0000000010100001010010110;
    rom[15193] = 25'b0000000010100001010010010;
    rom[15194] = 25'b0000000010100001010001111;
    rom[15195] = 25'b0000000010100001010001011;
    rom[15196] = 25'b0000000010100001010000110;
    rom[15197] = 25'b0000000010100001010000011;
    rom[15198] = 25'b0000000010100001001111110;
    rom[15199] = 25'b0000000010100001001111010;
    rom[15200] = 25'b0000000010100001001110101;
    rom[15201] = 25'b0000000010100001001110000;
    rom[15202] = 25'b0000000010100001001101011;
    rom[15203] = 25'b0000000010100001001100110;
    rom[15204] = 25'b0000000010100001001100010;
    rom[15205] = 25'b0000000010100001001011100;
    rom[15206] = 25'b0000000010100001001010111;
    rom[15207] = 25'b0000000010100001001010010;
    rom[15208] = 25'b0000000010100001001001100;
    rom[15209] = 25'b0000000010100001001000111;
    rom[15210] = 25'b0000000010100001001000001;
    rom[15211] = 25'b0000000010100001000111011;
    rom[15212] = 25'b0000000010100001000110101;
    rom[15213] = 25'b0000000010100001000101111;
    rom[15214] = 25'b0000000010100001000101001;
    rom[15215] = 25'b0000000010100001000100010;
    rom[15216] = 25'b0000000010100001000011100;
    rom[15217] = 25'b0000000010100001000010110;
    rom[15218] = 25'b0000000010100001000001111;
    rom[15219] = 25'b0000000010100001000001000;
    rom[15220] = 25'b0000000010100001000000001;
    rom[15221] = 25'b0000000010100000111111010;
    rom[15222] = 25'b0000000010100000111110010;
    rom[15223] = 25'b0000000010100000111101100;
    rom[15224] = 25'b0000000010100000111100100;
    rom[15225] = 25'b0000000010100000111011101;
    rom[15226] = 25'b0000000010100000111010101;
    rom[15227] = 25'b0000000010100000111001101;
    rom[15228] = 25'b0000000010100000111000101;
    rom[15229] = 25'b0000000010100000110111101;
    rom[15230] = 25'b0000000010100000110110101;
    rom[15231] = 25'b0000000010100000110101101;
    rom[15232] = 25'b0000000010100000110100100;
    rom[15233] = 25'b0000000010100000110011100;
    rom[15234] = 25'b0000000010100000110010100;
    rom[15235] = 25'b0000000010100000110001011;
    rom[15236] = 25'b0000000010100000110000010;
    rom[15237] = 25'b0000000010100000101111001;
    rom[15238] = 25'b0000000010100000101110000;
    rom[15239] = 25'b0000000010100000101100110;
    rom[15240] = 25'b0000000010100000101011101;
    rom[15241] = 25'b0000000010100000101010011;
    rom[15242] = 25'b0000000010100000101001010;
    rom[15243] = 25'b0000000010100000101000001;
    rom[15244] = 25'b0000000010100000100110110;
    rom[15245] = 25'b0000000010100000100101100;
    rom[15246] = 25'b0000000010100000100100011;
    rom[15247] = 25'b0000000010100000100011000;
    rom[15248] = 25'b0000000010100000100001110;
    rom[15249] = 25'b0000000010100000100000011;
    rom[15250] = 25'b0000000010100000011111001;
    rom[15251] = 25'b0000000010100000011101110;
    rom[15252] = 25'b0000000010100000011100011;
    rom[15253] = 25'b0000000010100000011011001;
    rom[15254] = 25'b0000000010100000011001110;
    rom[15255] = 25'b0000000010100000011000010;
    rom[15256] = 25'b0000000010100000010110111;
    rom[15257] = 25'b0000000010100000010101100;
    rom[15258] = 25'b0000000010100000010100000;
    rom[15259] = 25'b0000000010100000010010101;
    rom[15260] = 25'b0000000010100000010001001;
    rom[15261] = 25'b0000000010100000001111101;
    rom[15262] = 25'b0000000010100000001110001;
    rom[15263] = 25'b0000000010100000001100101;
    rom[15264] = 25'b0000000010100000001011000;
    rom[15265] = 25'b0000000010100000001001100;
    rom[15266] = 25'b0000000010100000001000000;
    rom[15267] = 25'b0000000010100000000110011;
    rom[15268] = 25'b0000000010100000000100110;
    rom[15269] = 25'b0000000010100000000011001;
    rom[15270] = 25'b0000000010100000000001101;
    rom[15271] = 25'b0000000010011111111111111;
    rom[15272] = 25'b0000000010011111111110010;
    rom[15273] = 25'b0000000010011111111100101;
    rom[15274] = 25'b0000000010011111111011000;
    rom[15275] = 25'b0000000010011111111001010;
    rom[15276] = 25'b0000000010011111110111100;
    rom[15277] = 25'b0000000010011111110101110;
    rom[15278] = 25'b0000000010011111110100000;
    rom[15279] = 25'b0000000010011111110010010;
    rom[15280] = 25'b0000000010011111110000100;
    rom[15281] = 25'b0000000010011111101110110;
    rom[15282] = 25'b0000000010011111101100111;
    rom[15283] = 25'b0000000010011111101011001;
    rom[15284] = 25'b0000000010011111101001010;
    rom[15285] = 25'b0000000010011111100111011;
    rom[15286] = 25'b0000000010011111100101100;
    rom[15287] = 25'b0000000010011111100011101;
    rom[15288] = 25'b0000000010011111100001110;
    rom[15289] = 25'b0000000010011111011111110;
    rom[15290] = 25'b0000000010011111011101111;
    rom[15291] = 25'b0000000010011111011100000;
    rom[15292] = 25'b0000000010011111011010000;
    rom[15293] = 25'b0000000010011111011000000;
    rom[15294] = 25'b0000000010011111010110000;
    rom[15295] = 25'b0000000010011111010100000;
    rom[15296] = 25'b0000000010011111010010000;
    rom[15297] = 25'b0000000010011111010000000;
    rom[15298] = 25'b0000000010011111001110000;
    rom[15299] = 25'b0000000010011111001011110;
    rom[15300] = 25'b0000000010011111001001110;
    rom[15301] = 25'b0000000010011111000111110;
    rom[15302] = 25'b0000000010011111000101100;
    rom[15303] = 25'b0000000010011111000011011;
    rom[15304] = 25'b0000000010011111000001010;
    rom[15305] = 25'b0000000010011110111111001;
    rom[15306] = 25'b0000000010011110111101000;
    rom[15307] = 25'b0000000010011110111010110;
    rom[15308] = 25'b0000000010011110111000101;
    rom[15309] = 25'b0000000010011110110110011;
    rom[15310] = 25'b0000000010011110110100001;
    rom[15311] = 25'b0000000010011110110001111;
    rom[15312] = 25'b0000000010011110101111100;
    rom[15313] = 25'b0000000010011110101101010;
    rom[15314] = 25'b0000000010011110101010111;
    rom[15315] = 25'b0000000010011110101000110;
    rom[15316] = 25'b0000000010011110100110011;
    rom[15317] = 25'b0000000010011110100011111;
    rom[15318] = 25'b0000000010011110100001101;
    rom[15319] = 25'b0000000010011110011111010;
    rom[15320] = 25'b0000000010011110011100111;
    rom[15321] = 25'b0000000010011110011010011;
    rom[15322] = 25'b0000000010011110011000000;
    rom[15323] = 25'b0000000010011110010101100;
    rom[15324] = 25'b0000000010011110010011001;
    rom[15325] = 25'b0000000010011110010000101;
    rom[15326] = 25'b0000000010011110001110001;
    rom[15327] = 25'b0000000010011110001011101;
    rom[15328] = 25'b0000000010011110001001001;
    rom[15329] = 25'b0000000010011110000110101;
    rom[15330] = 25'b0000000010011110000100001;
    rom[15331] = 25'b0000000010011110000001100;
    rom[15332] = 25'b0000000010011101111110111;
    rom[15333] = 25'b0000000010011101111100011;
    rom[15334] = 25'b0000000010011101111001110;
    rom[15335] = 25'b0000000010011101110111001;
    rom[15336] = 25'b0000000010011101110100011;
    rom[15337] = 25'b0000000010011101110001110;
    rom[15338] = 25'b0000000010011101101111001;
    rom[15339] = 25'b0000000010011101101100011;
    rom[15340] = 25'b0000000010011101101001101;
    rom[15341] = 25'b0000000010011101100111000;
    rom[15342] = 25'b0000000010011101100100010;
    rom[15343] = 25'b0000000010011101100001100;
    rom[15344] = 25'b0000000010011101011110110;
    rom[15345] = 25'b0000000010011101011011111;
    rom[15346] = 25'b0000000010011101011001001;
    rom[15347] = 25'b0000000010011101010110011;
    rom[15348] = 25'b0000000010011101010011011;
    rom[15349] = 25'b0000000010011101010000101;
    rom[15350] = 25'b0000000010011101001101110;
    rom[15351] = 25'b0000000010011101001010111;
    rom[15352] = 25'b0000000010011101001000000;
    rom[15353] = 25'b0000000010011101000101000;
    rom[15354] = 25'b0000000010011101000010001;
    rom[15355] = 25'b0000000010011100111111010;
    rom[15356] = 25'b0000000010011100111100010;
    rom[15357] = 25'b0000000010011100111001010;
    rom[15358] = 25'b0000000010011100110110010;
    rom[15359] = 25'b0000000010011100110011010;
    rom[15360] = 25'b0000000010011100110000011;
    rom[15361] = 25'b0000000010011100101101010;
    rom[15362] = 25'b0000000010011100101010001;
    rom[15363] = 25'b0000000010011100100111001;
    rom[15364] = 25'b0000000010011100100100000;
    rom[15365] = 25'b0000000010011100100000111;
    rom[15366] = 25'b0000000010011100011101111;
    rom[15367] = 25'b0000000010011100011010101;
    rom[15368] = 25'b0000000010011100010111101;
    rom[15369] = 25'b0000000010011100010100011;
    rom[15370] = 25'b0000000010011100010001010;
    rom[15371] = 25'b0000000010011100001110000;
    rom[15372] = 25'b0000000010011100001010110;
    rom[15373] = 25'b0000000010011100000111101;
    rom[15374] = 25'b0000000010011100000100011;
    rom[15375] = 25'b0000000010011100000001001;
    rom[15376] = 25'b0000000010011011111101110;
    rom[15377] = 25'b0000000010011011111010100;
    rom[15378] = 25'b0000000010011011110111001;
    rom[15379] = 25'b0000000010011011110011111;
    rom[15380] = 25'b0000000010011011110000100;
    rom[15381] = 25'b0000000010011011101101001;
    rom[15382] = 25'b0000000010011011101001110;
    rom[15383] = 25'b0000000010011011100110100;
    rom[15384] = 25'b0000000010011011100011001;
    rom[15385] = 25'b0000000010011011011111101;
    rom[15386] = 25'b0000000010011011011100001;
    rom[15387] = 25'b0000000010011011011000110;
    rom[15388] = 25'b0000000010011011010101010;
    rom[15389] = 25'b0000000010011011010001110;
    rom[15390] = 25'b0000000010011011001110011;
    rom[15391] = 25'b0000000010011011001010110;
    rom[15392] = 25'b0000000010011011000111010;
    rom[15393] = 25'b0000000010011011000011110;
    rom[15394] = 25'b0000000010011011000000001;
    rom[15395] = 25'b0000000010011010111100101;
    rom[15396] = 25'b0000000010011010111001000;
    rom[15397] = 25'b0000000010011010110101011;
    rom[15398] = 25'b0000000010011010110001110;
    rom[15399] = 25'b0000000010011010101110001;
    rom[15400] = 25'b0000000010011010101010100;
    rom[15401] = 25'b0000000010011010100110111;
    rom[15402] = 25'b0000000010011010100011001;
    rom[15403] = 25'b0000000010011010011111100;
    rom[15404] = 25'b0000000010011010011011110;
    rom[15405] = 25'b0000000010011010011000000;
    rom[15406] = 25'b0000000010011010010100010;
    rom[15407] = 25'b0000000010011010010000100;
    rom[15408] = 25'b0000000010011010001100110;
    rom[15409] = 25'b0000000010011010001000111;
    rom[15410] = 25'b0000000010011010000101000;
    rom[15411] = 25'b0000000010011010000001010;
    rom[15412] = 25'b0000000010011001111101011;
    rom[15413] = 25'b0000000010011001111001100;
    rom[15414] = 25'b0000000010011001110101101;
    rom[15415] = 25'b0000000010011001110001110;
    rom[15416] = 25'b0000000010011001101101111;
    rom[15417] = 25'b0000000010011001101010000;
    rom[15418] = 25'b0000000010011001100110000;
    rom[15419] = 25'b0000000010011001100010000;
    rom[15420] = 25'b0000000010011001011110001;
    rom[15421] = 25'b0000000010011001011010001;
    rom[15422] = 25'b0000000010011001010110001;
    rom[15423] = 25'b0000000010011001010010000;
    rom[15424] = 25'b0000000010011001001110000;
    rom[15425] = 25'b0000000010011001001001111;
    rom[15426] = 25'b0000000010011001000101111;
    rom[15427] = 25'b0000000010011001000001110;
    rom[15428] = 25'b0000000010011000111101110;
    rom[15429] = 25'b0000000010011000111001101;
    rom[15430] = 25'b0000000010011000110101100;
    rom[15431] = 25'b0000000010011000110001010;
    rom[15432] = 25'b0000000010011000101101001;
    rom[15433] = 25'b0000000010011000101001000;
    rom[15434] = 25'b0000000010011000100100110;
    rom[15435] = 25'b0000000010011000100000100;
    rom[15436] = 25'b0000000010011000011100011;
    rom[15437] = 25'b0000000010011000011000001;
    rom[15438] = 25'b0000000010011000010011110;
    rom[15439] = 25'b0000000010011000001111101;
    rom[15440] = 25'b0000000010011000001011010;
    rom[15441] = 25'b0000000010011000000111000;
    rom[15442] = 25'b0000000010011000000010101;
    rom[15443] = 25'b0000000010010111111110010;
    rom[15444] = 25'b0000000010010111111001111;
    rom[15445] = 25'b0000000010010111110101100;
    rom[15446] = 25'b0000000010010111110001001;
    rom[15447] = 25'b0000000010010111101100110;
    rom[15448] = 25'b0000000010010111101000011;
    rom[15449] = 25'b0000000010010111100011111;
    rom[15450] = 25'b0000000010010111011111011;
    rom[15451] = 25'b0000000010010111011011000;
    rom[15452] = 25'b0000000010010111010110100;
    rom[15453] = 25'b0000000010010111010001111;
    rom[15454] = 25'b0000000010010111001101100;
    rom[15455] = 25'b0000000010010111001000111;
    rom[15456] = 25'b0000000010010111000100011;
    rom[15457] = 25'b0000000010010110111111111;
    rom[15458] = 25'b0000000010010110111011010;
    rom[15459] = 25'b0000000010010110110110101;
    rom[15460] = 25'b0000000010010110110010000;
    rom[15461] = 25'b0000000010010110101101011;
    rom[15462] = 25'b0000000010010110101000110;
    rom[15463] = 25'b0000000010010110100100001;
    rom[15464] = 25'b0000000010010110011111011;
    rom[15465] = 25'b0000000010010110011010101;
    rom[15466] = 25'b0000000010010110010110000;
    rom[15467] = 25'b0000000010010110010001010;
    rom[15468] = 25'b0000000010010110001100100;
    rom[15469] = 25'b0000000010010110000111101;
    rom[15470] = 25'b0000000010010110000010111;
    rom[15471] = 25'b0000000010010101111110001;
    rom[15472] = 25'b0000000010010101111001010;
    rom[15473] = 25'b0000000010010101110100100;
    rom[15474] = 25'b0000000010010101101111101;
    rom[15475] = 25'b0000000010010101101010111;
    rom[15476] = 25'b0000000010010101100110000;
    rom[15477] = 25'b0000000010010101100001000;
    rom[15478] = 25'b0000000010010101011100001;
    rom[15479] = 25'b0000000010010101010111010;
    rom[15480] = 25'b0000000010010101010010010;
    rom[15481] = 25'b0000000010010101001101011;
    rom[15482] = 25'b0000000010010101001000011;
    rom[15483] = 25'b0000000010010101000011011;
    rom[15484] = 25'b0000000010010100111110011;
    rom[15485] = 25'b0000000010010100111001011;
    rom[15486] = 25'b0000000010010100110100010;
    rom[15487] = 25'b0000000010010100101111010;
    rom[15488] = 25'b0000000010010100101010010;
    rom[15489] = 25'b0000000010010100100101001;
    rom[15490] = 25'b0000000010010100100000000;
    rom[15491] = 25'b0000000010010100011010111;
    rom[15492] = 25'b0000000010010100010101110;
    rom[15493] = 25'b0000000010010100010000101;
    rom[15494] = 25'b0000000010010100001011100;
    rom[15495] = 25'b0000000010010100000110010;
    rom[15496] = 25'b0000000010010100000001001;
    rom[15497] = 25'b0000000010010011111011111;
    rom[15498] = 25'b0000000010010011110110101;
    rom[15499] = 25'b0000000010010011110001011;
    rom[15500] = 25'b0000000010010011101100010;
    rom[15501] = 25'b0000000010010011100110111;
    rom[15502] = 25'b0000000010010011100001100;
    rom[15503] = 25'b0000000010010011011100010;
    rom[15504] = 25'b0000000010010011010110111;
    rom[15505] = 25'b0000000010010011010001101;
    rom[15506] = 25'b0000000010010011001100010;
    rom[15507] = 25'b0000000010010011000110111;
    rom[15508] = 25'b0000000010010011000001100;
    rom[15509] = 25'b0000000010010010111100001;
    rom[15510] = 25'b0000000010010010110110101;
    rom[15511] = 25'b0000000010010010110001001;
    rom[15512] = 25'b0000000010010010101011110;
    rom[15513] = 25'b0000000010010010100110010;
    rom[15514] = 25'b0000000010010010100000111;
    rom[15515] = 25'b0000000010010010011011011;
    rom[15516] = 25'b0000000010010010010101111;
    rom[15517] = 25'b0000000010010010010000010;
    rom[15518] = 25'b0000000010010010001010110;
    rom[15519] = 25'b0000000010010010000101001;
    rom[15520] = 25'b0000000010010001111111100;
    rom[15521] = 25'b0000000010010001111001111;
    rom[15522] = 25'b0000000010010001110100010;
    rom[15523] = 25'b0000000010010001101110101;
    rom[15524] = 25'b0000000010010001101001000;
    rom[15525] = 25'b0000000010010001100011011;
    rom[15526] = 25'b0000000010010001011101110;
    rom[15527] = 25'b0000000010010001011000000;
    rom[15528] = 25'b0000000010010001010010010;
    rom[15529] = 25'b0000000010010001001100100;
    rom[15530] = 25'b0000000010010001000110110;
    rom[15531] = 25'b0000000010010001000001000;
    rom[15532] = 25'b0000000010010000111011010;
    rom[15533] = 25'b0000000010010000110101100;
    rom[15534] = 25'b0000000010010000101111101;
    rom[15535] = 25'b0000000010010000101001110;
    rom[15536] = 25'b0000000010010000100100000;
    rom[15537] = 25'b0000000010010000011110001;
    rom[15538] = 25'b0000000010010000011000010;
    rom[15539] = 25'b0000000010010000010010011;
    rom[15540] = 25'b0000000010010000001100100;
    rom[15541] = 25'b0000000010010000000110100;
    rom[15542] = 25'b0000000010010000000000101;
    rom[15543] = 25'b0000000010001111111010101;
    rom[15544] = 25'b0000000010001111110100101;
    rom[15545] = 25'b0000000010001111101110101;
    rom[15546] = 25'b0000000010001111101000101;
    rom[15547] = 25'b0000000010001111100010101;
    rom[15548] = 25'b0000000010001111011100100;
    rom[15549] = 25'b0000000010001111010110100;
    rom[15550] = 25'b0000000010001111010000011;
    rom[15551] = 25'b0000000010001111001010011;
    rom[15552] = 25'b0000000010001111000100010;
    rom[15553] = 25'b0000000010001110111110001;
    rom[15554] = 25'b0000000010001110111000000;
    rom[15555] = 25'b0000000010001110110001111;
    rom[15556] = 25'b0000000010001110101011110;
    rom[15557] = 25'b0000000010001110100101011;
    rom[15558] = 25'b0000000010001110011111010;
    rom[15559] = 25'b0000000010001110011001000;
    rom[15560] = 25'b0000000010001110010010111;
    rom[15561] = 25'b0000000010001110001100101;
    rom[15562] = 25'b0000000010001110000110011;
    rom[15563] = 25'b0000000010001110000000000;
    rom[15564] = 25'b0000000010001101111001110;
    rom[15565] = 25'b0000000010001101110011011;
    rom[15566] = 25'b0000000010001101101101000;
    rom[15567] = 25'b0000000010001101100110101;
    rom[15568] = 25'b0000000010001101100000011;
    rom[15569] = 25'b0000000010001101011010000;
    rom[15570] = 25'b0000000010001101010011101;
    rom[15571] = 25'b0000000010001101001101001;
    rom[15572] = 25'b0000000010001101000110110;
    rom[15573] = 25'b0000000010001101000000010;
    rom[15574] = 25'b0000000010001100111001111;
    rom[15575] = 25'b0000000010001100110011011;
    rom[15576] = 25'b0000000010001100101100111;
    rom[15577] = 25'b0000000010001100100110011;
    rom[15578] = 25'b0000000010001100011111110;
    rom[15579] = 25'b0000000010001100011001010;
    rom[15580] = 25'b0000000010001100010010110;
    rom[15581] = 25'b0000000010001100001100010;
    rom[15582] = 25'b0000000010001100000101100;
    rom[15583] = 25'b0000000010001011111110111;
    rom[15584] = 25'b0000000010001011111000010;
    rom[15585] = 25'b0000000010001011110001101;
    rom[15586] = 25'b0000000010001011101011000;
    rom[15587] = 25'b0000000010001011100100011;
    rom[15588] = 25'b0000000010001011011101101;
    rom[15589] = 25'b0000000010001011010111000;
    rom[15590] = 25'b0000000010001011010000010;
    rom[15591] = 25'b0000000010001011001001100;
    rom[15592] = 25'b0000000010001011000010110;
    rom[15593] = 25'b0000000010001010111100000;
    rom[15594] = 25'b0000000010001010110101010;
    rom[15595] = 25'b0000000010001010101110011;
    rom[15596] = 25'b0000000010001010100111101;
    rom[15597] = 25'b0000000010001010100000110;
    rom[15598] = 25'b0000000010001010011001111;
    rom[15599] = 25'b0000000010001010010011001;
    rom[15600] = 25'b0000000010001010001100001;
    rom[15601] = 25'b0000000010001010000101010;
    rom[15602] = 25'b0000000010001001111110011;
    rom[15603] = 25'b0000000010001001110111011;
    rom[15604] = 25'b0000000010001001110000011;
    rom[15605] = 25'b0000000010001001101001100;
    rom[15606] = 25'b0000000010001001100010100;
    rom[15607] = 25'b0000000010001001011011100;
    rom[15608] = 25'b0000000010001001010100100;
    rom[15609] = 25'b0000000010001001001101100;
    rom[15610] = 25'b0000000010001001000110011;
    rom[15611] = 25'b0000000010001000111111011;
    rom[15612] = 25'b0000000010001000111000010;
    rom[15613] = 25'b0000000010001000110001010;
    rom[15614] = 25'b0000000010001000101010001;
    rom[15615] = 25'b0000000010001000100010111;
    rom[15616] = 25'b0000000010001000011011110;
    rom[15617] = 25'b0000000010001000010100101;
    rom[15618] = 25'b0000000010001000001101011;
    rom[15619] = 25'b0000000010001000000110010;
    rom[15620] = 25'b0000000010000111111111000;
    rom[15621] = 25'b0000000010000111110111111;
    rom[15622] = 25'b0000000010000111110000101;
    rom[15623] = 25'b0000000010000111101001011;
    rom[15624] = 25'b0000000010000111100010001;
    rom[15625] = 25'b0000000010000111011010111;
    rom[15626] = 25'b0000000010000111010011100;
    rom[15627] = 25'b0000000010000111001100001;
    rom[15628] = 25'b0000000010000111000100111;
    rom[15629] = 25'b0000000010000110111101100;
    rom[15630] = 25'b0000000010000110110110001;
    rom[15631] = 25'b0000000010000110101110110;
    rom[15632] = 25'b0000000010000110100111011;
    rom[15633] = 25'b0000000010000110011111111;
    rom[15634] = 25'b0000000010000110011000011;
    rom[15635] = 25'b0000000010000110010001000;
    rom[15636] = 25'b0000000010000110001001101;
    rom[15637] = 25'b0000000010000110000010001;
    rom[15638] = 25'b0000000010000101111010100;
    rom[15639] = 25'b0000000010000101110011000;
    rom[15640] = 25'b0000000010000101101011100;
    rom[15641] = 25'b0000000010000101100011111;
    rom[15642] = 25'b0000000010000101011100011;
    rom[15643] = 25'b0000000010000101010100110;
    rom[15644] = 25'b0000000010000101001101010;
    rom[15645] = 25'b0000000010000101000101101;
    rom[15646] = 25'b0000000010000100111110000;
    rom[15647] = 25'b0000000010000100110110011;
    rom[15648] = 25'b0000000010000100101110110;
    rom[15649] = 25'b0000000010000100100111000;
    rom[15650] = 25'b0000000010000100011111010;
    rom[15651] = 25'b0000000010000100010111101;
    rom[15652] = 25'b0000000010000100001111111;
    rom[15653] = 25'b0000000010000100001000001;
    rom[15654] = 25'b0000000010000100000000011;
    rom[15655] = 25'b0000000010000011111000101;
    rom[15656] = 25'b0000000010000011110000110;
    rom[15657] = 25'b0000000010000011101001000;
    rom[15658] = 25'b0000000010000011100001010;
    rom[15659] = 25'b0000000010000011011001011;
    rom[15660] = 25'b0000000010000011010001100;
    rom[15661] = 25'b0000000010000011001001101;
    rom[15662] = 25'b0000000010000011000001110;
    rom[15663] = 25'b0000000010000010111001111;
    rom[15664] = 25'b0000000010000010110001111;
    rom[15665] = 25'b0000000010000010101010000;
    rom[15666] = 25'b0000000010000010100010000;
    rom[15667] = 25'b0000000010000010011010000;
    rom[15668] = 25'b0000000010000010010010001;
    rom[15669] = 25'b0000000010000010001010000;
    rom[15670] = 25'b0000000010000010000010000;
    rom[15671] = 25'b0000000010000001111010000;
    rom[15672] = 25'b0000000010000001110010000;
    rom[15673] = 25'b0000000010000001101001111;
    rom[15674] = 25'b0000000010000001100001110;
    rom[15675] = 25'b0000000010000001011001110;
    rom[15676] = 25'b0000000010000001010001101;
    rom[15677] = 25'b0000000010000001001001100;
    rom[15678] = 25'b0000000010000001000001010;
    rom[15679] = 25'b0000000010000000111001001;
    rom[15680] = 25'b0000000010000000110001000;
    rom[15681] = 25'b0000000010000000101000111;
    rom[15682] = 25'b0000000010000000100000101;
    rom[15683] = 25'b0000000010000000011000011;
    rom[15684] = 25'b0000000010000000010000010;
    rom[15685] = 25'b0000000010000000000111111;
    rom[15686] = 25'b0000000001111111111111101;
    rom[15687] = 25'b0000000001111111110111011;
    rom[15688] = 25'b0000000001111111101111000;
    rom[15689] = 25'b0000000001111111100110110;
    rom[15690] = 25'b0000000001111111011110011;
    rom[15691] = 25'b0000000001111111010110000;
    rom[15692] = 25'b0000000001111111001101101;
    rom[15693] = 25'b0000000001111111000101010;
    rom[15694] = 25'b0000000001111110111100111;
    rom[15695] = 25'b0000000001111110110100100;
    rom[15696] = 25'b0000000001111110101100000;
    rom[15697] = 25'b0000000001111110100011101;
    rom[15698] = 25'b0000000001111110011011001;
    rom[15699] = 25'b0000000001111110010010101;
    rom[15700] = 25'b0000000001111110001010001;
    rom[15701] = 25'b0000000001111110000001101;
    rom[15702] = 25'b0000000001111101111001001;
    rom[15703] = 25'b0000000001111101110000100;
    rom[15704] = 25'b0000000001111101101000000;
    rom[15705] = 25'b0000000001111101011111011;
    rom[15706] = 25'b0000000001111101010110111;
    rom[15707] = 25'b0000000001111101001110010;
    rom[15708] = 25'b0000000001111101000101100;
    rom[15709] = 25'b0000000001111100111101000;
    rom[15710] = 25'b0000000001111100110100010;
    rom[15711] = 25'b0000000001111100101011101;
    rom[15712] = 25'b0000000001111100100010111;
    rom[15713] = 25'b0000000001111100011010010;
    rom[15714] = 25'b0000000001111100010001011;
    rom[15715] = 25'b0000000001111100001000110;
    rom[15716] = 25'b0000000001111100000000000;
    rom[15717] = 25'b0000000001111011110111010;
    rom[15718] = 25'b0000000001111011101110011;
    rom[15719] = 25'b0000000001111011100101101;
    rom[15720] = 25'b0000000001111011011100110;
    rom[15721] = 25'b0000000001111011010100000;
    rom[15722] = 25'b0000000001111011001011001;
    rom[15723] = 25'b0000000001111011000010010;
    rom[15724] = 25'b0000000001111010111001011;
    rom[15725] = 25'b0000000001111010110000100;
    rom[15726] = 25'b0000000001111010100111100;
    rom[15727] = 25'b0000000001111010011110101;
    rom[15728] = 25'b0000000001111010010101110;
    rom[15729] = 25'b0000000001111010001100110;
    rom[15730] = 25'b0000000001111010000011110;
    rom[15731] = 25'b0000000001111001111010110;
    rom[15732] = 25'b0000000001111001110001110;
    rom[15733] = 25'b0000000001111001101000101;
    rom[15734] = 25'b0000000001111001011111110;
    rom[15735] = 25'b0000000001111001010110101;
    rom[15736] = 25'b0000000001111001001101101;
    rom[15737] = 25'b0000000001111001000100100;
    rom[15738] = 25'b0000000001111000111011011;
    rom[15739] = 25'b0000000001111000110010010;
    rom[15740] = 25'b0000000001111000101001001;
    rom[15741] = 25'b0000000001111000011111111;
    rom[15742] = 25'b0000000001111000010110110;
    rom[15743] = 25'b0000000001111000001101101;
    rom[15744] = 25'b0000000001111000000100011;
    rom[15745] = 25'b0000000001110111111011010;
    rom[15746] = 25'b0000000001110111110010000;
    rom[15747] = 25'b0000000001110111101000110;
    rom[15748] = 25'b0000000001110111011111100;
    rom[15749] = 25'b0000000001110111010110001;
    rom[15750] = 25'b0000000001110111001100111;
    rom[15751] = 25'b0000000001110111000011101;
    rom[15752] = 25'b0000000001110110111010010;
    rom[15753] = 25'b0000000001110110110000111;
    rom[15754] = 25'b0000000001110110100111100;
    rom[15755] = 25'b0000000001110110011110001;
    rom[15756] = 25'b0000000001110110010100110;
    rom[15757] = 25'b0000000001110110001011011;
    rom[15758] = 25'b0000000001110110000001111;
    rom[15759] = 25'b0000000001110101111000100;
    rom[15760] = 25'b0000000001110101101111000;
    rom[15761] = 25'b0000000001110101100101101;
    rom[15762] = 25'b0000000001110101011100001;
    rom[15763] = 25'b0000000001110101010010101;
    rom[15764] = 25'b0000000001110101001001001;
    rom[15765] = 25'b0000000001110100111111100;
    rom[15766] = 25'b0000000001110100110110000;
    rom[15767] = 25'b0000000001110100101100100;
    rom[15768] = 25'b0000000001110100100010111;
    rom[15769] = 25'b0000000001110100011001011;
    rom[15770] = 25'b0000000001110100001111110;
    rom[15771] = 25'b0000000001110100000110001;
    rom[15772] = 25'b0000000001110011111100011;
    rom[15773] = 25'b0000000001110011110010110;
    rom[15774] = 25'b0000000001110011101001000;
    rom[15775] = 25'b0000000001110011011111011;
    rom[15776] = 25'b0000000001110011010101110;
    rom[15777] = 25'b0000000001110011001100000;
    rom[15778] = 25'b0000000001110011000010010;
    rom[15779] = 25'b0000000001110010111000100;
    rom[15780] = 25'b0000000001110010101110101;
    rom[15781] = 25'b0000000001110010100101000;
    rom[15782] = 25'b0000000001110010011011001;
    rom[15783] = 25'b0000000001110010010001011;
    rom[15784] = 25'b0000000001110010000111100;
    rom[15785] = 25'b0000000001110001111101101;
    rom[15786] = 25'b0000000001110001110011110;
    rom[15787] = 25'b0000000001110001101001111;
    rom[15788] = 25'b0000000001110001100000000;
    rom[15789] = 25'b0000000001110001010110000;
    rom[15790] = 25'b0000000001110001001100001;
    rom[15791] = 25'b0000000001110001000010010;
    rom[15792] = 25'b0000000001110000111000010;
    rom[15793] = 25'b0000000001110000101110010;
    rom[15794] = 25'b0000000001110000100100010;
    rom[15795] = 25'b0000000001110000011010010;
    rom[15796] = 25'b0000000001110000010000010;
    rom[15797] = 25'b0000000001110000000110010;
    rom[15798] = 25'b0000000001101111111100010;
    rom[15799] = 25'b0000000001101111110010001;
    rom[15800] = 25'b0000000001101111101000000;
    rom[15801] = 25'b0000000001101111011110000;
    rom[15802] = 25'b0000000001101111010011111;
    rom[15803] = 25'b0000000001101111001001110;
    rom[15804] = 25'b0000000001101110111111101;
    rom[15805] = 25'b0000000001101110110101011;
    rom[15806] = 25'b0000000001101110101011010;
    rom[15807] = 25'b0000000001101110100001001;
    rom[15808] = 25'b0000000001101110010110111;
    rom[15809] = 25'b0000000001101110001100101;
    rom[15810] = 25'b0000000001101110000010100;
    rom[15811] = 25'b0000000001101101111000001;
    rom[15812] = 25'b0000000001101101101101111;
    rom[15813] = 25'b0000000001101101100011101;
    rom[15814] = 25'b0000000001101101011001011;
    rom[15815] = 25'b0000000001101101001111000;
    rom[15816] = 25'b0000000001101101000100110;
    rom[15817] = 25'b0000000001101100111010011;
    rom[15818] = 25'b0000000001101100110000000;
    rom[15819] = 25'b0000000001101100100101101;
    rom[15820] = 25'b0000000001101100011011010;
    rom[15821] = 25'b0000000001101100010000110;
    rom[15822] = 25'b0000000001101100000110011;
    rom[15823] = 25'b0000000001101011111100000;
    rom[15824] = 25'b0000000001101011110001100;
    rom[15825] = 25'b0000000001101011100111000;
    rom[15826] = 25'b0000000001101011011100101;
    rom[15827] = 25'b0000000001101011010010000;
    rom[15828] = 25'b0000000001101011000111101;
    rom[15829] = 25'b0000000001101010111101000;
    rom[15830] = 25'b0000000001101010110010100;
    rom[15831] = 25'b0000000001101010100111111;
    rom[15832] = 25'b0000000001101010011101011;
    rom[15833] = 25'b0000000001101010010010110;
    rom[15834] = 25'b0000000001101010001000001;
    rom[15835] = 25'b0000000001101001111101100;
    rom[15836] = 25'b0000000001101001110010111;
    rom[15837] = 25'b0000000001101001101000010;
    rom[15838] = 25'b0000000001101001011101101;
    rom[15839] = 25'b0000000001101001010010111;
    rom[15840] = 25'b0000000001101001001000010;
    rom[15841] = 25'b0000000001101000111101100;
    rom[15842] = 25'b0000000001101000110010110;
    rom[15843] = 25'b0000000001101000101000000;
    rom[15844] = 25'b0000000001101000011101010;
    rom[15845] = 25'b0000000001101000010010100;
    rom[15846] = 25'b0000000001101000000111101;
    rom[15847] = 25'b0000000001100111111100111;
    rom[15848] = 25'b0000000001100111110010000;
    rom[15849] = 25'b0000000001100111100111001;
    rom[15850] = 25'b0000000001100111011100011;
    rom[15851] = 25'b0000000001100111010001100;
    rom[15852] = 25'b0000000001100111000110101;
    rom[15853] = 25'b0000000001100110111011110;
    rom[15854] = 25'b0000000001100110110000110;
    rom[15855] = 25'b0000000001100110100101111;
    rom[15856] = 25'b0000000001100110011011000;
    rom[15857] = 25'b0000000001100110010000000;
    rom[15858] = 25'b0000000001100110000101000;
    rom[15859] = 25'b0000000001100101111010000;
    rom[15860] = 25'b0000000001100101101111000;
    rom[15861] = 25'b0000000001100101100100000;
    rom[15862] = 25'b0000000001100101011000111;
    rom[15863] = 25'b0000000001100101001101111;
    rom[15864] = 25'b0000000001100101000010110;
    rom[15865] = 25'b0000000001100100110111110;
    rom[15866] = 25'b0000000001100100101100101;
    rom[15867] = 25'b0000000001100100100001100;
    rom[15868] = 25'b0000000001100100010110100;
    rom[15869] = 25'b0000000001100100001011011;
    rom[15870] = 25'b0000000001100100000000001;
    rom[15871] = 25'b0000000001100011110101000;
    rom[15872] = 25'b0000000001100011101001110;
    rom[15873] = 25'b0000000001100011011110101;
    rom[15874] = 25'b0000000001100011010011011;
    rom[15875] = 25'b0000000001100011001000001;
    rom[15876] = 25'b0000000001100010111100111;
    rom[15877] = 25'b0000000001100010110001101;
    rom[15878] = 25'b0000000001100010100110011;
    rom[15879] = 25'b0000000001100010011011001;
    rom[15880] = 25'b0000000001100010001111110;
    rom[15881] = 25'b0000000001100010000100100;
    rom[15882] = 25'b0000000001100001111001001;
    rom[15883] = 25'b0000000001100001101101110;
    rom[15884] = 25'b0000000001100001100010011;
    rom[15885] = 25'b0000000001100001010111000;
    rom[15886] = 25'b0000000001100001001011101;
    rom[15887] = 25'b0000000001100001000000010;
    rom[15888] = 25'b0000000001100000110100111;
    rom[15889] = 25'b0000000001100000101001011;
    rom[15890] = 25'b0000000001100000011101111;
    rom[15891] = 25'b0000000001100000010010100;
    rom[15892] = 25'b0000000001100000000111000;
    rom[15893] = 25'b0000000001011111111011011;
    rom[15894] = 25'b0000000001011111101111111;
    rom[15895] = 25'b0000000001011111100100011;
    rom[15896] = 25'b0000000001011111011000111;
    rom[15897] = 25'b0000000001011111001101010;
    rom[15898] = 25'b0000000001011111000001101;
    rom[15899] = 25'b0000000001011110110110001;
    rom[15900] = 25'b0000000001011110101010100;
    rom[15901] = 25'b0000000001011110011110111;
    rom[15902] = 25'b0000000001011110010011010;
    rom[15903] = 25'b0000000001011110000111101;
    rom[15904] = 25'b0000000001011101111011111;
    rom[15905] = 25'b0000000001011101110000010;
    rom[15906] = 25'b0000000001011101100100101;
    rom[15907] = 25'b0000000001011101011000111;
    rom[15908] = 25'b0000000001011101001101001;
    rom[15909] = 25'b0000000001011101000001011;
    rom[15910] = 25'b0000000001011100110101101;
    rom[15911] = 25'b0000000001011100101001111;
    rom[15912] = 25'b0000000001011100011110000;
    rom[15913] = 25'b0000000001011100010010010;
    rom[15914] = 25'b0000000001011100000110011;
    rom[15915] = 25'b0000000001011011111010101;
    rom[15916] = 25'b0000000001011011101110110;
    rom[15917] = 25'b0000000001011011100011000;
    rom[15918] = 25'b0000000001011011010111001;
    rom[15919] = 25'b0000000001011011001011010;
    rom[15920] = 25'b0000000001011010111111010;
    rom[15921] = 25'b0000000001011010110011011;
    rom[15922] = 25'b0000000001011010100111100;
    rom[15923] = 25'b0000000001011010011011100;
    rom[15924] = 25'b0000000001011010001111100;
    rom[15925] = 25'b0000000001011010000011101;
    rom[15926] = 25'b0000000001011001110111100;
    rom[15927] = 25'b0000000001011001101011101;
    rom[15928] = 25'b0000000001011001011111100;
    rom[15929] = 25'b0000000001011001010011100;
    rom[15930] = 25'b0000000001011001000111100;
    rom[15931] = 25'b0000000001011000111011011;
    rom[15932] = 25'b0000000001011000101111011;
    rom[15933] = 25'b0000000001011000100011010;
    rom[15934] = 25'b0000000001011000010111001;
    rom[15935] = 25'b0000000001011000001011000;
    rom[15936] = 25'b0000000001010111111110111;
    rom[15937] = 25'b0000000001010111110010110;
    rom[15938] = 25'b0000000001010111100110101;
    rom[15939] = 25'b0000000001010111011010011;
    rom[15940] = 25'b0000000001010111001110010;
    rom[15941] = 25'b0000000001010111000010000;
    rom[15942] = 25'b0000000001010110110101110;
    rom[15943] = 25'b0000000001010110101001100;
    rom[15944] = 25'b0000000001010110011101010;
    rom[15945] = 25'b0000000001010110010001001;
    rom[15946] = 25'b0000000001010110000100110;
    rom[15947] = 25'b0000000001010101111000011;
    rom[15948] = 25'b0000000001010101101100001;
    rom[15949] = 25'b0000000001010101011111111;
    rom[15950] = 25'b0000000001010101010011011;
    rom[15951] = 25'b0000000001010101000111001;
    rom[15952] = 25'b0000000001010100111010110;
    rom[15953] = 25'b0000000001010100101110011;
    rom[15954] = 25'b0000000001010100100010000;
    rom[15955] = 25'b0000000001010100010101101;
    rom[15956] = 25'b0000000001010100001001010;
    rom[15957] = 25'b0000000001010011111100101;
    rom[15958] = 25'b0000000001010011110000010;
    rom[15959] = 25'b0000000001010011100011111;
    rom[15960] = 25'b0000000001010011010111011;
    rom[15961] = 25'b0000000001010011001010110;
    rom[15962] = 25'b0000000001010010111110010;
    rom[15963] = 25'b0000000001010010110001110;
    rom[15964] = 25'b0000000001010010100101010;
    rom[15965] = 25'b0000000001010010011000101;
    rom[15966] = 25'b0000000001010010001100001;
    rom[15967] = 25'b0000000001010001111111100;
    rom[15968] = 25'b0000000001010001110010111;
    rom[15969] = 25'b0000000001010001100110011;
    rom[15970] = 25'b0000000001010001011001110;
    rom[15971] = 25'b0000000001010001001101001;
    rom[15972] = 25'b0000000001010001000000011;
    rom[15973] = 25'b0000000001010000110011110;
    rom[15974] = 25'b0000000001010000100111001;
    rom[15975] = 25'b0000000001010000011010011;
    rom[15976] = 25'b0000000001010000001101110;
    rom[15977] = 25'b0000000001010000000000111;
    rom[15978] = 25'b0000000001001111110100010;
    rom[15979] = 25'b0000000001001111100111011;
    rom[15980] = 25'b0000000001001111011010110;
    rom[15981] = 25'b0000000001001111001101111;
    rom[15982] = 25'b0000000001001111000001001;
    rom[15983] = 25'b0000000001001110110100011;
    rom[15984] = 25'b0000000001001110100111100;
    rom[15985] = 25'b0000000001001110011010101;
    rom[15986] = 25'b0000000001001110001101110;
    rom[15987] = 25'b0000000001001110000001000;
    rom[15988] = 25'b0000000001001101110100001;
    rom[15989] = 25'b0000000001001101100111010;
    rom[15990] = 25'b0000000001001101011010010;
    rom[15991] = 25'b0000000001001101001101011;
    rom[15992] = 25'b0000000001001101000000011;
    rom[15993] = 25'b0000000001001100110011100;
    rom[15994] = 25'b0000000001001100100110100;
    rom[15995] = 25'b0000000001001100011001100;
    rom[15996] = 25'b0000000001001100001100100;
    rom[15997] = 25'b0000000001001011111111100;
    rom[15998] = 25'b0000000001001011110010100;
    rom[15999] = 25'b0000000001001011100101100;
    rom[16000] = 25'b0000000001001011011000011;
    rom[16001] = 25'b0000000001001011001011011;
    rom[16002] = 25'b0000000001001010111110010;
    rom[16003] = 25'b0000000001001010110001001;
    rom[16004] = 25'b0000000001001010100100001;
    rom[16005] = 25'b0000000001001010010111000;
    rom[16006] = 25'b0000000001001010001001111;
    rom[16007] = 25'b0000000001001001111100110;
    rom[16008] = 25'b0000000001001001101111100;
    rom[16009] = 25'b0000000001001001100010011;
    rom[16010] = 25'b0000000001001001010101010;
    rom[16011] = 25'b0000000001001001000111111;
    rom[16012] = 25'b0000000001001000111010110;
    rom[16013] = 25'b0000000001001000101101100;
    rom[16014] = 25'b0000000001001000100000011;
    rom[16015] = 25'b0000000001001000010011001;
    rom[16016] = 25'b0000000001001000000101111;
    rom[16017] = 25'b0000000001000111111000100;
    rom[16018] = 25'b0000000001000111101011010;
    rom[16019] = 25'b0000000001000111011101111;
    rom[16020] = 25'b0000000001000111010000101;
    rom[16021] = 25'b0000000001000111000011010;
    rom[16022] = 25'b0000000001000110110101111;
    rom[16023] = 25'b0000000001000110101000100;
    rom[16024] = 25'b0000000001000110011011001;
    rom[16025] = 25'b0000000001000110001101110;
    rom[16026] = 25'b0000000001000110000000011;
    rom[16027] = 25'b0000000001000101110010111;
    rom[16028] = 25'b0000000001000101100101100;
    rom[16029] = 25'b0000000001000101011000000;
    rom[16030] = 25'b0000000001000101001010101;
    rom[16031] = 25'b0000000001000100111101001;
    rom[16032] = 25'b0000000001000100101111101;
    rom[16033] = 25'b0000000001000100100010001;
    rom[16034] = 25'b0000000001000100010100101;
    rom[16035] = 25'b0000000001000100000111000;
    rom[16036] = 25'b0000000001000011111001100;
    rom[16037] = 25'b0000000001000011101100000;
    rom[16038] = 25'b0000000001000011011110011;
    rom[16039] = 25'b0000000001000011010000110;
    rom[16040] = 25'b0000000001000011000011010;
    rom[16041] = 25'b0000000001000010110101101;
    rom[16042] = 25'b0000000001000010101000000;
    rom[16043] = 25'b0000000001000010011010011;
    rom[16044] = 25'b0000000001000010001100110;
    rom[16045] = 25'b0000000001000001111111001;
    rom[16046] = 25'b0000000001000001110001011;
    rom[16047] = 25'b0000000001000001100011110;
    rom[16048] = 25'b0000000001000001010110000;
    rom[16049] = 25'b0000000001000001001000010;
    rom[16050] = 25'b0000000001000000111010100;
    rom[16051] = 25'b0000000001000000101100110;
    rom[16052] = 25'b0000000001000000011111001;
    rom[16053] = 25'b0000000001000000010001010;
    rom[16054] = 25'b0000000001000000000011100;
    rom[16055] = 25'b0000000000111111110101110;
    rom[16056] = 25'b0000000000111111100111111;
    rom[16057] = 25'b0000000000111111011010001;
    rom[16058] = 25'b0000000000111111001100010;
    rom[16059] = 25'b0000000000111110111110011;
    rom[16060] = 25'b0000000000111110110000100;
    rom[16061] = 25'b0000000000111110100010110;
    rom[16062] = 25'b0000000000111110010100110;
    rom[16063] = 25'b0000000000111110000110111;
    rom[16064] = 25'b0000000000111101111001000;
    rom[16065] = 25'b0000000000111101101011000;
    rom[16066] = 25'b0000000000111101011101001;
    rom[16067] = 25'b0000000000111101001111001;
    rom[16068] = 25'b0000000000111101000001010;
    rom[16069] = 25'b0000000000111100110011010;
    rom[16070] = 25'b0000000000111100100101001;
    rom[16071] = 25'b0000000000111100010111001;
    rom[16072] = 25'b0000000000111100001001001;
    rom[16073] = 25'b0000000000111011111011001;
    rom[16074] = 25'b0000000000111011101101000;
    rom[16075] = 25'b0000000000111011011111000;
    rom[16076] = 25'b0000000000111011010001000;
    rom[16077] = 25'b0000000000111011000010111;
    rom[16078] = 25'b0000000000111010110100110;
    rom[16079] = 25'b0000000000111010100110101;
    rom[16080] = 25'b0000000000111010011000100;
    rom[16081] = 25'b0000000000111010001010011;
    rom[16082] = 25'b0000000000111001111100010;
    rom[16083] = 25'b0000000000111001101110001;
    rom[16084] = 25'b0000000000111001100000000;
    rom[16085] = 25'b0000000000111001010001110;
    rom[16086] = 25'b0000000000111001000011100;
    rom[16087] = 25'b0000000000111000110101011;
    rom[16088] = 25'b0000000000111000100111001;
    rom[16089] = 25'b0000000000111000011000111;
    rom[16090] = 25'b0000000000111000001010101;
    rom[16091] = 25'b0000000000110111111100010;
    rom[16092] = 25'b0000000000110111101110000;
    rom[16093] = 25'b0000000000110111011111110;
    rom[16094] = 25'b0000000000110111010001100;
    rom[16095] = 25'b0000000000110111000011001;
    rom[16096] = 25'b0000000000110110110100111;
    rom[16097] = 25'b0000000000110110100110100;
    rom[16098] = 25'b0000000000110110011000001;
    rom[16099] = 25'b0000000000110110001001110;
    rom[16100] = 25'b0000000000110101111011011;
    rom[16101] = 25'b0000000000110101101101000;
    rom[16102] = 25'b0000000000110101011110101;
    rom[16103] = 25'b0000000000110101010000010;
    rom[16104] = 25'b0000000000110101000001110;
    rom[16105] = 25'b0000000000110100110011010;
    rom[16106] = 25'b0000000000110100100100111;
    rom[16107] = 25'b0000000000110100010110011;
    rom[16108] = 25'b0000000000110100000111111;
    rom[16109] = 25'b0000000000110011111001011;
    rom[16110] = 25'b0000000000110011101010111;
    rom[16111] = 25'b0000000000110011011100011;
    rom[16112] = 25'b0000000000110011001101111;
    rom[16113] = 25'b0000000000110010111111010;
    rom[16114] = 25'b0000000000110010110000101;
    rom[16115] = 25'b0000000000110010100010001;
    rom[16116] = 25'b0000000000110010010011100;
    rom[16117] = 25'b0000000000110010000101000;
    rom[16118] = 25'b0000000000110001110110011;
    rom[16119] = 25'b0000000000110001100111110;
    rom[16120] = 25'b0000000000110001011001001;
    rom[16121] = 25'b0000000000110001001010100;
    rom[16122] = 25'b0000000000110000111011111;
    rom[16123] = 25'b0000000000110000101101001;
    rom[16124] = 25'b0000000000110000011110100;
    rom[16125] = 25'b0000000000110000001111110;
    rom[16126] = 25'b0000000000110000000001000;
    rom[16127] = 25'b0000000000101111110010011;
    rom[16128] = 25'b0000000000101111100011101;
    rom[16129] = 25'b0000000000101111010100111;
    rom[16130] = 25'b0000000000101111000110001;
    rom[16131] = 25'b0000000000101110110111011;
    rom[16132] = 25'b0000000000101110101000101;
    rom[16133] = 25'b0000000000101110011001110;
    rom[16134] = 25'b0000000000101110001011000;
    rom[16135] = 25'b0000000000101101111100001;
    rom[16136] = 25'b0000000000101101101101010;
    rom[16137] = 25'b0000000000101101011110100;
    rom[16138] = 25'b0000000000101101001111101;
    rom[16139] = 25'b0000000000101101000000110;
    rom[16140] = 25'b0000000000101100110001111;
    rom[16141] = 25'b0000000000101100100011000;
    rom[16142] = 25'b0000000000101100010100001;
    rom[16143] = 25'b0000000000101100000101001;
    rom[16144] = 25'b0000000000101011110110010;
    rom[16145] = 25'b0000000000101011100111011;
    rom[16146] = 25'b0000000000101011011000011;
    rom[16147] = 25'b0000000000101011001001011;
    rom[16148] = 25'b0000000000101010111010100;
    rom[16149] = 25'b0000000000101010101011011;
    rom[16150] = 25'b0000000000101010011100100;
    rom[16151] = 25'b0000000000101010001101011;
    rom[16152] = 25'b0000000000101001111110011;
    rom[16153] = 25'b0000000000101001101111011;
    rom[16154] = 25'b0000000000101001100000011;
    rom[16155] = 25'b0000000000101001010001010;
    rom[16156] = 25'b0000000000101001000010001;
    rom[16157] = 25'b0000000000101000110011001;
    rom[16158] = 25'b0000000000101000100100000;
    rom[16159] = 25'b0000000000101000010101000;
    rom[16160] = 25'b0000000000101000000101111;
    rom[16161] = 25'b0000000000100111110110110;
    rom[16162] = 25'b0000000000100111100111101;
    rom[16163] = 25'b0000000000100111011000011;
    rom[16164] = 25'b0000000000100111001001010;
    rom[16165] = 25'b0000000000100110111010000;
    rom[16166] = 25'b0000000000100110101010111;
    rom[16167] = 25'b0000000000100110011011101;
    rom[16168] = 25'b0000000000100110001100011;
    rom[16169] = 25'b0000000000100101111101010;
    rom[16170] = 25'b0000000000100101101110000;
    rom[16171] = 25'b0000000000100101011110110;
    rom[16172] = 25'b0000000000100101001111100;
    rom[16173] = 25'b0000000000100101000000010;
    rom[16174] = 25'b0000000000100100110000111;
    rom[16175] = 25'b0000000000100100100001101;
    rom[16176] = 25'b0000000000100100010010010;
    rom[16177] = 25'b0000000000100100000011000;
    rom[16178] = 25'b0000000000100011110011101;
    rom[16179] = 25'b0000000000100011100100011;
    rom[16180] = 25'b0000000000100011010101000;
    rom[16181] = 25'b0000000000100011000101101;
    rom[16182] = 25'b0000000000100010110110010;
    rom[16183] = 25'b0000000000100010100110111;
    rom[16184] = 25'b0000000000100010010111100;
    rom[16185] = 25'b0000000000100010001000001;
    rom[16186] = 25'b0000000000100001111000101;
    rom[16187] = 25'b0000000000100001101001010;
    rom[16188] = 25'b0000000000100001011001110;
    rom[16189] = 25'b0000000000100001001010011;
    rom[16190] = 25'b0000000000100000111010111;
    rom[16191] = 25'b0000000000100000101011011;
    rom[16192] = 25'b0000000000100000011011111;
    rom[16193] = 25'b0000000000100000001100011;
    rom[16194] = 25'b0000000000011111111100111;
    rom[16195] = 25'b0000000000011111101101011;
    rom[16196] = 25'b0000000000011111011101111;
    rom[16197] = 25'b0000000000011111001110010;
    rom[16198] = 25'b0000000000011110111110110;
    rom[16199] = 25'b0000000000011110101111001;
    rom[16200] = 25'b0000000000011110011111100;
    rom[16201] = 25'b0000000000011110010000000;
    rom[16202] = 25'b0000000000011110000000011;
    rom[16203] = 25'b0000000000011101110000110;
    rom[16204] = 25'b0000000000011101100001001;
    rom[16205] = 25'b0000000000011101010001100;
    rom[16206] = 25'b0000000000011101000001111;
    rom[16207] = 25'b0000000000011100110010001;
    rom[16208] = 25'b0000000000011100100010100;
    rom[16209] = 25'b0000000000011100010010110;
    rom[16210] = 25'b0000000000011100000011001;
    rom[16211] = 25'b0000000000011011110011011;
    rom[16212] = 25'b0000000000011011100011110;
    rom[16213] = 25'b0000000000011011010100000;
    rom[16214] = 25'b0000000000011011000100010;
    rom[16215] = 25'b0000000000011010110100100;
    rom[16216] = 25'b0000000000011010100100110;
    rom[16217] = 25'b0000000000011010010101000;
    rom[16218] = 25'b0000000000011010000101010;
    rom[16219] = 25'b0000000000011001110101100;
    rom[16220] = 25'b0000000000011001100101101;
    rom[16221] = 25'b0000000000011001010101110;
    rom[16222] = 25'b0000000000011001000110000;
    rom[16223] = 25'b0000000000011000110110001;
    rom[16224] = 25'b0000000000011000100110011;
    rom[16225] = 25'b0000000000011000010110100;
    rom[16226] = 25'b0000000000011000000110101;
    rom[16227] = 25'b0000000000010111110110110;
    rom[16228] = 25'b0000000000010111100110111;
    rom[16229] = 25'b0000000000010111010111000;
    rom[16230] = 25'b0000000000010111000111000;
    rom[16231] = 25'b0000000000010110110111001;
    rom[16232] = 25'b0000000000010110100111001;
    rom[16233] = 25'b0000000000010110010111001;
    rom[16234] = 25'b0000000000010110000111010;
    rom[16235] = 25'b0000000000010101110111011;
    rom[16236] = 25'b0000000000010101100111011;
    rom[16237] = 25'b0000000000010101010111010;
    rom[16238] = 25'b0000000000010101000111011;
    rom[16239] = 25'b0000000000010100110111011;
    rom[16240] = 25'b0000000000010100100111010;
    rom[16241] = 25'b0000000000010100010111011;
    rom[16242] = 25'b0000000000010100000111010;
    rom[16243] = 25'b0000000000010011110111010;
    rom[16244] = 25'b0000000000010011100111001;
    rom[16245] = 25'b0000000000010011010111001;
    rom[16246] = 25'b0000000000010011000111000;
    rom[16247] = 25'b0000000000010010110111000;
    rom[16248] = 25'b0000000000010010100110110;
    rom[16249] = 25'b0000000000010010010110110;
    rom[16250] = 25'b0000000000010010000110101;
    rom[16251] = 25'b0000000000010001110110011;
    rom[16252] = 25'b0000000000010001100110011;
    rom[16253] = 25'b0000000000010001010110010;
    rom[16254] = 25'b0000000000010001000110000;
    rom[16255] = 25'b0000000000010000110101110;
    rom[16256] = 25'b0000000000010000100101101;
    rom[16257] = 25'b0000000000010000010101100;
    rom[16258] = 25'b0000000000010000000101010;
    rom[16259] = 25'b0000000000001111110101000;
    rom[16260] = 25'b0000000000001111100100111;
    rom[16261] = 25'b0000000000001111010100101;
    rom[16262] = 25'b0000000000001111000100011;
    rom[16263] = 25'b0000000000001110110100001;
    rom[16264] = 25'b0000000000001110100011111;
    rom[16265] = 25'b0000000000001110010011100;
    rom[16266] = 25'b0000000000001110000011010;
    rom[16267] = 25'b0000000000001101110011000;
    rom[16268] = 25'b0000000000001101100010101;
    rom[16269] = 25'b0000000000001101010010011;
    rom[16270] = 25'b0000000000001101000010000;
    rom[16271] = 25'b0000000000001100110001110;
    rom[16272] = 25'b0000000000001100100001010;
    rom[16273] = 25'b0000000000001100010001000;
    rom[16274] = 25'b0000000000001100000000101;
    rom[16275] = 25'b0000000000001011110000010;
    rom[16276] = 25'b0000000000001011011111111;
    rom[16277] = 25'b0000000000001011001111100;
    rom[16278] = 25'b0000000000001010111111000;
    rom[16279] = 25'b0000000000001010101110101;
    rom[16280] = 25'b0000000000001010011110001;
    rom[16281] = 25'b0000000000001010001101110;
    rom[16282] = 25'b0000000000001001111101010;
    rom[16283] = 25'b0000000000001001101100111;
    rom[16284] = 25'b0000000000001001011100011;
    rom[16285] = 25'b0000000000001001001011111;
    rom[16286] = 25'b0000000000001000111011100;
    rom[16287] = 25'b0000000000001000101010111;
    rom[16288] = 25'b0000000000001000011010011;
    rom[16289] = 25'b0000000000001000001010000;
    rom[16290] = 25'b0000000000000111111001100;
    rom[16291] = 25'b0000000000000111101000111;
    rom[16292] = 25'b0000000000000111011000011;
    rom[16293] = 25'b0000000000000111000111110;
    rom[16294] = 25'b0000000000000110110111010;
    rom[16295] = 25'b0000000000000110100110101;
    rom[16296] = 25'b0000000000000110010110001;
    rom[16297] = 25'b0000000000000110000101100;
    rom[16298] = 25'b0000000000000101110100111;
    rom[16299] = 25'b0000000000000101100100010;
    rom[16300] = 25'b0000000000000101010011101;
    rom[16301] = 25'b0000000000000101000011000;
    rom[16302] = 25'b0000000000000100110010011;
    rom[16303] = 25'b0000000000000100100001110;
    rom[16304] = 25'b0000000000000100010001001;
    rom[16305] = 25'b0000000000000100000000011;
    rom[16306] = 25'b0000000000000011101111110;
    rom[16307] = 25'b0000000000000011011111000;
    rom[16308] = 25'b0000000000000011001110011;
    rom[16309] = 25'b0000000000000010111101101;
    rom[16310] = 25'b0000000000000010101100111;
    rom[16311] = 25'b0000000000000010011100001;
    rom[16312] = 25'b0000000000000010001011100;
    rom[16313] = 25'b0000000000000001111010110;
    rom[16314] = 25'b0000000000000001101010000;
    rom[16315] = 25'b0000000000000001011001010;
    rom[16316] = 25'b0000000000000001001000100;
    rom[16317] = 25'b0000000000000000110111110;
    rom[16318] = 25'b0000000000000000100110111;
    rom[16319] = 25'b0000000000000000010110001;
    rom[16320] = 25'b0000000000000000000101010;
    rom[16321] = 25'b1111111111111111110100100;
    rom[16322] = 25'b1111111111111111100011110;
    rom[16323] = 25'b1111111111111111010010111;
    rom[16324] = 25'b1111111111111111000010000;
    rom[16325] = 25'b1111111111111110110001010;
    rom[16326] = 25'b1111111111111110100000010;
    rom[16327] = 25'b1111111111111110001111100;
    rom[16328] = 25'b1111111111111101111110101;
    rom[16329] = 25'b1111111111111101101101110;
    rom[16330] = 25'b1111111111111101011100110;
    rom[16331] = 25'b1111111111111101001011111;
    rom[16332] = 25'b1111111111111100111011000;
    rom[16333] = 25'b1111111111111100101010001;
    rom[16334] = 25'b1111111111111100011001001;
    rom[16335] = 25'b1111111111111100001000001;
    rom[16336] = 25'b1111111111111011110111010;
    rom[16337] = 25'b1111111111111011100110010;
    rom[16338] = 25'b1111111111111011010101010;
    rom[16339] = 25'b1111111111111011000100011;
    rom[16340] = 25'b1111111111111010110011011;
    rom[16341] = 25'b1111111111111010100010011;
    rom[16342] = 25'b1111111111111010010001011;
    rom[16343] = 25'b1111111111111010000000010;
    rom[16344] = 25'b1111111111111001101111010;
    rom[16345] = 25'b1111111111111001011110010;
    rom[16346] = 25'b1111111111111001001101010;
    rom[16347] = 25'b1111111111111000111100010;
    rom[16348] = 25'b1111111111111000101011001;
    rom[16349] = 25'b1111111111111000011010001;
    rom[16350] = 25'b1111111111111000001001000;
    rom[16351] = 25'b1111111111110111111000000;
    rom[16352] = 25'b1111111111110111100110111;
    rom[16353] = 25'b1111111111110111010101110;
    rom[16354] = 25'b1111111111110111000100110;
    rom[16355] = 25'b1111111111110110110011100;
    rom[16356] = 25'b1111111111110110100010011;
    rom[16357] = 25'b1111111111110110010001010;
    rom[16358] = 25'b1111111111110110000000001;
    rom[16359] = 25'b1111111111110101101111000;
    rom[16360] = 25'b1111111111110101011101111;
    rom[16361] = 25'b1111111111110101001100101;
    rom[16362] = 25'b1111111111110100111011100;
    rom[16363] = 25'b1111111111110100101010011;
    rom[16364] = 25'b1111111111110100011001001;
    rom[16365] = 25'b1111111111110100001000000;
    rom[16366] = 25'b1111111111110011110110101;
    rom[16367] = 25'b1111111111110011100101100;
    rom[16368] = 25'b1111111111110011010100010;
    rom[16369] = 25'b1111111111110011000011000;
    rom[16370] = 25'b1111111111110010110001110;
    rom[16371] = 25'b1111111111110010100000101;
    rom[16372] = 25'b1111111111110010001111010;
    rom[16373] = 25'b1111111111110001111110000;
    rom[16374] = 25'b1111111111110001101100110;
    rom[16375] = 25'b1111111111110001011011100;
    rom[16376] = 25'b1111111111110001001010010;
    rom[16377] = 25'b1111111111110000111000111;
    rom[16378] = 25'b1111111111110000100111100;
    rom[16379] = 25'b1111111111110000010110010;
    rom[16380] = 25'b1111111111110000000101000;
    rom[16381] = 25'b1111111111101111110011101;
    rom[16382] = 25'b1111111111101111100010010;
    rom[16383] = 25'b1111111111101111010001000;
    rom[16384] = 25'b1111111111101110111111101;
    rom[16385] = 25'b1111111111101110101110010;
    rom[16386] = 25'b1111111111101110011100111;
    rom[16387] = 25'b1111111111101110001011100;
    rom[16388] = 25'b1111111111101101111010001;
    rom[16389] = 25'b1111111111101101101000110;
    rom[16390] = 25'b1111111111101101010111010;
    rom[16391] = 25'b1111111111101101000101111;
    rom[16392] = 25'b1111111111101100110100100;
    rom[16393] = 25'b1111111111101100100011001;
    rom[16394] = 25'b1111111111101100010001101;
    rom[16395] = 25'b1111111111101100000000001;
    rom[16396] = 25'b1111111111101011101110110;
    rom[16397] = 25'b1111111111101011011101011;
    rom[16398] = 25'b1111111111101011001011111;
    rom[16399] = 25'b1111111111101010111010011;
    rom[16400] = 25'b1111111111101010101000111;
    rom[16401] = 25'b1111111111101010010111011;
    rom[16402] = 25'b1111111111101010000101111;
    rom[16403] = 25'b1111111111101001110100100;
    rom[16404] = 25'b1111111111101001100010111;
    rom[16405] = 25'b1111111111101001010001011;
    rom[16406] = 25'b1111111111101000111111111;
    rom[16407] = 25'b1111111111101000101110011;
    rom[16408] = 25'b1111111111101000011100110;
    rom[16409] = 25'b1111111111101000001011010;
    rom[16410] = 25'b1111111111100111111001110;
    rom[16411] = 25'b1111111111100111101000010;
    rom[16412] = 25'b1111111111100111010110101;
    rom[16413] = 25'b1111111111100111000101000;
    rom[16414] = 25'b1111111111100110110011011;
    rom[16415] = 25'b1111111111100110100001111;
    rom[16416] = 25'b1111111111100110010000010;
    rom[16417] = 25'b1111111111100101111110101;
    rom[16418] = 25'b1111111111100101101101000;
    rom[16419] = 25'b1111111111100101011011100;
    rom[16420] = 25'b1111111111100101001001110;
    rom[16421] = 25'b1111111111100100111000001;
    rom[16422] = 25'b1111111111100100100110100;
    rom[16423] = 25'b1111111111100100010100111;
    rom[16424] = 25'b1111111111100100000011010;
    rom[16425] = 25'b1111111111100011110001100;
    rom[16426] = 25'b1111111111100011011111111;
    rom[16427] = 25'b1111111111100011001110010;
    rom[16428] = 25'b1111111111100010111100100;
    rom[16429] = 25'b1111111111100010101010111;
    rom[16430] = 25'b1111111111100010011001010;
    rom[16431] = 25'b1111111111100010000111100;
    rom[16432] = 25'b1111111111100001110101110;
    rom[16433] = 25'b1111111111100001100100001;
    rom[16434] = 25'b1111111111100001010010011;
    rom[16435] = 25'b1111111111100001000000101;
    rom[16436] = 25'b1111111111100000101110111;
    rom[16437] = 25'b1111111111100000011101001;
    rom[16438] = 25'b1111111111100000001011011;
    rom[16439] = 25'b1111111111011111111001101;
    rom[16440] = 25'b1111111111011111100111111;
    rom[16441] = 25'b1111111111011111010110001;
    rom[16442] = 25'b1111111111011111000100010;
    rom[16443] = 25'b1111111111011110110010100;
    rom[16444] = 25'b1111111111011110100000110;
    rom[16445] = 25'b1111111111011110001111000;
    rom[16446] = 25'b1111111111011101111101001;
    rom[16447] = 25'b1111111111011101101011010;
    rom[16448] = 25'b1111111111011101011001100;
    rom[16449] = 25'b1111111111011101000111110;
    rom[16450] = 25'b1111111111011100110101111;
    rom[16451] = 25'b1111111111011100100100000;
    rom[16452] = 25'b1111111111011100010010010;
    rom[16453] = 25'b1111111111011100000000011;
    rom[16454] = 25'b1111111111011011101110100;
    rom[16455] = 25'b1111111111011011011100101;
    rom[16456] = 25'b1111111111011011001010110;
    rom[16457] = 25'b1111111111011010111000111;
    rom[16458] = 25'b1111111111011010100111000;
    rom[16459] = 25'b1111111111011010010101001;
    rom[16460] = 25'b1111111111011010000011010;
    rom[16461] = 25'b1111111111011001110001010;
    rom[16462] = 25'b1111111111011001011111100;
    rom[16463] = 25'b1111111111011001001101100;
    rom[16464] = 25'b1111111111011000111011101;
    rom[16465] = 25'b1111111111011000101001101;
    rom[16466] = 25'b1111111111011000010111110;
    rom[16467] = 25'b1111111111011000000101110;
    rom[16468] = 25'b1111111111010111110011111;
    rom[16469] = 25'b1111111111010111100001111;
    rom[16470] = 25'b1111111111010111001111111;
    rom[16471] = 25'b1111111111010110111110000;
    rom[16472] = 25'b1111111111010110101100000;
    rom[16473] = 25'b1111111111010110011010000;
    rom[16474] = 25'b1111111111010110001000001;
    rom[16475] = 25'b1111111111010101110110001;
    rom[16476] = 25'b1111111111010101100100000;
    rom[16477] = 25'b1111111111010101010010001;
    rom[16478] = 25'b1111111111010101000000001;
    rom[16479] = 25'b1111111111010100101110001;
    rom[16480] = 25'b1111111111010100011100000;
    rom[16481] = 25'b1111111111010100001010000;
    rom[16482] = 25'b1111111111010011111000000;
    rom[16483] = 25'b1111111111010011100110000;
    rom[16484] = 25'b1111111111010011010100000;
    rom[16485] = 25'b1111111111010011000001111;
    rom[16486] = 25'b1111111111010010101111111;
    rom[16487] = 25'b1111111111010010011101110;
    rom[16488] = 25'b1111111111010010001011110;
    rom[16489] = 25'b1111111111010001111001101;
    rom[16490] = 25'b1111111111010001100111101;
    rom[16491] = 25'b1111111111010001010101100;
    rom[16492] = 25'b1111111111010001000011011;
    rom[16493] = 25'b1111111111010000110001011;
    rom[16494] = 25'b1111111111010000011111010;
    rom[16495] = 25'b1111111111010000001101001;
    rom[16496] = 25'b1111111111001111111011000;
    rom[16497] = 25'b1111111111001111101000111;
    rom[16498] = 25'b1111111111001111010110110;
    rom[16499] = 25'b1111111111001111000100101;
    rom[16500] = 25'b1111111111001110110010100;
    rom[16501] = 25'b1111111111001110100000011;
    rom[16502] = 25'b1111111111001110001110011;
    rom[16503] = 25'b1111111111001101111100001;
    rom[16504] = 25'b1111111111001101101010000;
    rom[16505] = 25'b1111111111001101010111111;
    rom[16506] = 25'b1111111111001101000101101;
    rom[16507] = 25'b1111111111001100110011100;
    rom[16508] = 25'b1111111111001100100001011;
    rom[16509] = 25'b1111111111001100001111010;
    rom[16510] = 25'b1111111111001011111101000;
    rom[16511] = 25'b1111111111001011101010110;
    rom[16512] = 25'b1111111111001011011000101;
    rom[16513] = 25'b1111111111001011000110100;
    rom[16514] = 25'b1111111111001010110100010;
    rom[16515] = 25'b1111111111001010100010000;
    rom[16516] = 25'b1111111111001010001111111;
    rom[16517] = 25'b1111111111001001111101101;
    rom[16518] = 25'b1111111111001001101011011;
    rom[16519] = 25'b1111111111001001011001001;
    rom[16520] = 25'b1111111111001001000110111;
    rom[16521] = 25'b1111111111001000110100110;
    rom[16522] = 25'b1111111111001000100010100;
    rom[16523] = 25'b1111111111001000010000001;
    rom[16524] = 25'b1111111111000111111110000;
    rom[16525] = 25'b1111111111000111101011101;
    rom[16526] = 25'b1111111111000111011001100;
    rom[16527] = 25'b1111111111000111000111001;
    rom[16528] = 25'b1111111111000110110100111;
    rom[16529] = 25'b1111111111000110100010101;
    rom[16530] = 25'b1111111111000110010000011;
    rom[16531] = 25'b1111111111000101111110000;
    rom[16532] = 25'b1111111111000101101011110;
    rom[16533] = 25'b1111111111000101011001100;
    rom[16534] = 25'b1111111111000101000111010;
    rom[16535] = 25'b1111111111000100110100111;
    rom[16536] = 25'b1111111111000100100010101;
    rom[16537] = 25'b1111111111000100010000010;
    rom[16538] = 25'b1111111111000011111101111;
    rom[16539] = 25'b1111111111000011101011101;
    rom[16540] = 25'b1111111111000011011001010;
    rom[16541] = 25'b1111111111000011000111000;
    rom[16542] = 25'b1111111111000010110100101;
    rom[16543] = 25'b1111111111000010100010010;
    rom[16544] = 25'b1111111111000010010000000;
    rom[16545] = 25'b1111111111000001111101101;
    rom[16546] = 25'b1111111111000001101011010;
    rom[16547] = 25'b1111111111000001011000111;
    rom[16548] = 25'b1111111111000001000110100;
    rom[16549] = 25'b1111111111000000110100001;
    rom[16550] = 25'b1111111111000000100001110;
    rom[16551] = 25'b1111111111000000001111011;
    rom[16552] = 25'b1111111110111111111101001;
    rom[16553] = 25'b1111111110111111101010110;
    rom[16554] = 25'b1111111110111111011000010;
    rom[16555] = 25'b1111111110111111000101111;
    rom[16556] = 25'b1111111110111110110011100;
    rom[16557] = 25'b1111111110111110100001001;
    rom[16558] = 25'b1111111110111110001110110;
    rom[16559] = 25'b1111111110111101111100010;
    rom[16560] = 25'b1111111110111101101001111;
    rom[16561] = 25'b1111111110111101010111011;
    rom[16562] = 25'b1111111110111101000101000;
    rom[16563] = 25'b1111111110111100110010101;
    rom[16564] = 25'b1111111110111100100000010;
    rom[16565] = 25'b1111111110111100001101110;
    rom[16566] = 25'b1111111110111011111011011;
    rom[16567] = 25'b1111111110111011101000111;
    rom[16568] = 25'b1111111110111011010110100;
    rom[16569] = 25'b1111111110111011000100000;
    rom[16570] = 25'b1111111110111010110001101;
    rom[16571] = 25'b1111111110111010011111001;
    rom[16572] = 25'b1111111110111010001100101;
    rom[16573] = 25'b1111111110111001111010001;
    rom[16574] = 25'b1111111110111001100111110;
    rom[16575] = 25'b1111111110111001010101010;
    rom[16576] = 25'b1111111110111001000010110;
    rom[16577] = 25'b1111111110111000110000011;
    rom[16578] = 25'b1111111110111000011101111;
    rom[16579] = 25'b1111111110111000001011011;
    rom[16580] = 25'b1111111110110111111000111;
    rom[16581] = 25'b1111111110110111100110011;
    rom[16582] = 25'b1111111110110111010011111;
    rom[16583] = 25'b1111111110110111000001011;
    rom[16584] = 25'b1111111110110110101110111;
    rom[16585] = 25'b1111111110110110011100011;
    rom[16586] = 25'b1111111110110110001001111;
    rom[16587] = 25'b1111111110110101110111011;
    rom[16588] = 25'b1111111110110101100100111;
    rom[16589] = 25'b1111111110110101010010011;
    rom[16590] = 25'b1111111110110100111111111;
    rom[16591] = 25'b1111111110110100101101010;
    rom[16592] = 25'b1111111110110100011010110;
    rom[16593] = 25'b1111111110110100001000001;
    rom[16594] = 25'b1111111110110011110101110;
    rom[16595] = 25'b1111111110110011100011010;
    rom[16596] = 25'b1111111110110011010000101;
    rom[16597] = 25'b1111111110110010111110000;
    rom[16598] = 25'b1111111110110010101011100;
    rom[16599] = 25'b1111111110110010011001000;
    rom[16600] = 25'b1111111110110010000110100;
    rom[16601] = 25'b1111111110110001110011111;
    rom[16602] = 25'b1111111110110001100001010;
    rom[16603] = 25'b1111111110110001001110110;
    rom[16604] = 25'b1111111110110000111100010;
    rom[16605] = 25'b1111111110110000101001101;
    rom[16606] = 25'b1111111110110000010111000;
    rom[16607] = 25'b1111111110110000000100100;
    rom[16608] = 25'b1111111110101111110001111;
    rom[16609] = 25'b1111111110101111011111010;
    rom[16610] = 25'b1111111110101111001100110;
    rom[16611] = 25'b1111111110101110111010001;
    rom[16612] = 25'b1111111110101110100111100;
    rom[16613] = 25'b1111111110101110010101000;
    rom[16614] = 25'b1111111110101110000010011;
    rom[16615] = 25'b1111111110101101101111110;
    rom[16616] = 25'b1111111110101101011101010;
    rom[16617] = 25'b1111111110101101001010101;
    rom[16618] = 25'b1111111110101100111000000;
    rom[16619] = 25'b1111111110101100100101011;
    rom[16620] = 25'b1111111110101100010010110;
    rom[16621] = 25'b1111111110101100000000010;
    rom[16622] = 25'b1111111110101011101101100;
    rom[16623] = 25'b1111111110101011011011000;
    rom[16624] = 25'b1111111110101011001000011;
    rom[16625] = 25'b1111111110101010110101101;
    rom[16626] = 25'b1111111110101010100011001;
    rom[16627] = 25'b1111111110101010010000011;
    rom[16628] = 25'b1111111110101001111101111;
    rom[16629] = 25'b1111111110101001101011010;
    rom[16630] = 25'b1111111110101001011000101;
    rom[16631] = 25'b1111111110101001000101111;
    rom[16632] = 25'b1111111110101000110011011;
    rom[16633] = 25'b1111111110101000100000101;
    rom[16634] = 25'b1111111110101000001110000;
    rom[16635] = 25'b1111111110100111111011011;
    rom[16636] = 25'b1111111110100111101000110;
    rom[16637] = 25'b1111111110100111010110001;
    rom[16638] = 25'b1111111110100111000011100;
    rom[16639] = 25'b1111111110100110110000110;
    rom[16640] = 25'b1111111110100110011110001;
    rom[16641] = 25'b1111111110100110001011100;
    rom[16642] = 25'b1111111110100101111000111;
    rom[16643] = 25'b1111111110100101100110001;
    rom[16644] = 25'b1111111110100101010011100;
    rom[16645] = 25'b1111111110100101000000111;
    rom[16646] = 25'b1111111110100100101110010;
    rom[16647] = 25'b1111111110100100011011100;
    rom[16648] = 25'b1111111110100100001000111;
    rom[16649] = 25'b1111111110100011110110001;
    rom[16650] = 25'b1111111110100011100011100;
    rom[16651] = 25'b1111111110100011010000111;
    rom[16652] = 25'b1111111110100010111110001;
    rom[16653] = 25'b1111111110100010101011100;
    rom[16654] = 25'b1111111110100010011000110;
    rom[16655] = 25'b1111111110100010000110001;
    rom[16656] = 25'b1111111110100001110011011;
    rom[16657] = 25'b1111111110100001100000110;
    rom[16658] = 25'b1111111110100001001110001;
    rom[16659] = 25'b1111111110100000111011011;
    rom[16660] = 25'b1111111110100000101000101;
    rom[16661] = 25'b1111111110100000010110000;
    rom[16662] = 25'b1111111110100000000011010;
    rom[16663] = 25'b1111111110011111110000101;
    rom[16664] = 25'b1111111110011111011101111;
    rom[16665] = 25'b1111111110011111001011010;
    rom[16666] = 25'b1111111110011110111000100;
    rom[16667] = 25'b1111111110011110100101110;
    rom[16668] = 25'b1111111110011110010011001;
    rom[16669] = 25'b1111111110011110000000100;
    rom[16670] = 25'b1111111110011101101101101;
    rom[16671] = 25'b1111111110011101011011000;
    rom[16672] = 25'b1111111110011101001000011;
    rom[16673] = 25'b1111111110011100110101100;
    rom[16674] = 25'b1111111110011100100010111;
    rom[16675] = 25'b1111111110011100010000010;
    rom[16676] = 25'b1111111110011011111101011;
    rom[16677] = 25'b1111111110011011101010110;
    rom[16678] = 25'b1111111110011011011000000;
    rom[16679] = 25'b1111111110011011000101010;
    rom[16680] = 25'b1111111110011010110010101;
    rom[16681] = 25'b1111111110011010011111111;
    rom[16682] = 25'b1111111110011010001101001;
    rom[16683] = 25'b1111111110011001111010011;
    rom[16684] = 25'b1111111110011001100111110;
    rom[16685] = 25'b1111111110011001010101000;
    rom[16686] = 25'b1111111110011001000010010;
    rom[16687] = 25'b1111111110011000101111101;
    rom[16688] = 25'b1111111110011000011100111;
    rom[16689] = 25'b1111111110011000001010001;
    rom[16690] = 25'b1111111110010111110111011;
    rom[16691] = 25'b1111111110010111100100110;
    rom[16692] = 25'b1111111110010111010001111;
    rom[16693] = 25'b1111111110010110111111010;
    rom[16694] = 25'b1111111110010110101100100;
    rom[16695] = 25'b1111111110010110011001110;
    rom[16696] = 25'b1111111110010110000111000;
    rom[16697] = 25'b1111111110010101110100010;
    rom[16698] = 25'b1111111110010101100001101;
    rom[16699] = 25'b1111111110010101001110110;
    rom[16700] = 25'b1111111110010100111100001;
    rom[16701] = 25'b1111111110010100101001011;
    rom[16702] = 25'b1111111110010100010110101;
    rom[16703] = 25'b1111111110010100000011111;
    rom[16704] = 25'b1111111110010011110001001;
    rom[16705] = 25'b1111111110010011011110100;
    rom[16706] = 25'b1111111110010011001011110;
    rom[16707] = 25'b1111111110010010111001000;
    rom[16708] = 25'b1111111110010010100110010;
    rom[16709] = 25'b1111111110010010010011100;
    rom[16710] = 25'b1111111110010010000000110;
    rom[16711] = 25'b1111111110010001101110000;
    rom[16712] = 25'b1111111110010001011011010;
    rom[16713] = 25'b1111111110010001001000101;
    rom[16714] = 25'b1111111110010000110101110;
    rom[16715] = 25'b1111111110010000100011001;
    rom[16716] = 25'b1111111110010000010000011;
    rom[16717] = 25'b1111111110001111111101101;
    rom[16718] = 25'b1111111110001111101010111;
    rom[16719] = 25'b1111111110001111011000001;
    rom[16720] = 25'b1111111110001111000101011;
    rom[16721] = 25'b1111111110001110110010110;
    rom[16722] = 25'b1111111110001110011111111;
    rom[16723] = 25'b1111111110001110001101010;
    rom[16724] = 25'b1111111110001101111010100;
    rom[16725] = 25'b1111111110001101100111110;
    rom[16726] = 25'b1111111110001101010101000;
    rom[16727] = 25'b1111111110001101000010010;
    rom[16728] = 25'b1111111110001100101111101;
    rom[16729] = 25'b1111111110001100011100110;
    rom[16730] = 25'b1111111110001100001010000;
    rom[16731] = 25'b1111111110001011110111011;
    rom[16732] = 25'b1111111110001011100100101;
    rom[16733] = 25'b1111111110001011010001111;
    rom[16734] = 25'b1111111110001010111111001;
    rom[16735] = 25'b1111111110001010101100011;
    rom[16736] = 25'b1111111110001010011001110;
    rom[16737] = 25'b1111111110001010000110111;
    rom[16738] = 25'b1111111110001001110100010;
    rom[16739] = 25'b1111111110001001100001100;
    rom[16740] = 25'b1111111110001001001110110;
    rom[16741] = 25'b1111111110001000111100000;
    rom[16742] = 25'b1111111110001000101001010;
    rom[16743] = 25'b1111111110001000010110101;
    rom[16744] = 25'b1111111110001000000011110;
    rom[16745] = 25'b1111111110000111110001001;
    rom[16746] = 25'b1111111110000111011110011;
    rom[16747] = 25'b1111111110000111001011101;
    rom[16748] = 25'b1111111110000110111000111;
    rom[16749] = 25'b1111111110000110100110010;
    rom[16750] = 25'b1111111110000110010011100;
    rom[16751] = 25'b1111111110000110000000110;
    rom[16752] = 25'b1111111110000101101110000;
    rom[16753] = 25'b1111111110000101011011011;
    rom[16754] = 25'b1111111110000101001000101;
    rom[16755] = 25'b1111111110000100110101111;
    rom[16756] = 25'b1111111110000100100011001;
    rom[16757] = 25'b1111111110000100010000100;
    rom[16758] = 25'b1111111110000011111101110;
    rom[16759] = 25'b1111111110000011101011000;
    rom[16760] = 25'b1111111110000011011000011;
    rom[16761] = 25'b1111111110000011000101100;
    rom[16762] = 25'b1111111110000010110010111;
    rom[16763] = 25'b1111111110000010100000001;
    rom[16764] = 25'b1111111110000010001101011;
    rom[16765] = 25'b1111111110000001111010110;
    rom[16766] = 25'b1111111110000001101000000;
    rom[16767] = 25'b1111111110000001010101010;
    rom[16768] = 25'b1111111110000001000010101;
    rom[16769] = 25'b1111111110000000101111111;
    rom[16770] = 25'b1111111110000000011101010;
    rom[16771] = 25'b1111111110000000001010100;
    rom[16772] = 25'b1111111101111111110111110;
    rom[16773] = 25'b1111111101111111100101001;
    rom[16774] = 25'b1111111101111111010010100;
    rom[16775] = 25'b1111111101111110111111110;
    rom[16776] = 25'b1111111101111110101101000;
    rom[16777] = 25'b1111111101111110011010011;
    rom[16778] = 25'b1111111101111110000111101;
    rom[16779] = 25'b1111111101111101110101000;
    rom[16780] = 25'b1111111101111101100010010;
    rom[16781] = 25'b1111111101111101001111101;
    rom[16782] = 25'b1111111101111100111101000;
    rom[16783] = 25'b1111111101111100101010010;
    rom[16784] = 25'b1111111101111100010111101;
    rom[16785] = 25'b1111111101111100000100111;
    rom[16786] = 25'b1111111101111011110010010;
    rom[16787] = 25'b1111111101111011011111100;
    rom[16788] = 25'b1111111101111011001100111;
    rom[16789] = 25'b1111111101111010111010010;
    rom[16790] = 25'b1111111101111010100111100;
    rom[16791] = 25'b1111111101111010010100111;
    rom[16792] = 25'b1111111101111010000010001;
    rom[16793] = 25'b1111111101111001101111100;
    rom[16794] = 25'b1111111101111001011100111;
    rom[16795] = 25'b1111111101111001001010010;
    rom[16796] = 25'b1111111101111000110111100;
    rom[16797] = 25'b1111111101111000100100111;
    rom[16798] = 25'b1111111101111000010010010;
    rom[16799] = 25'b1111111101110111111111101;
    rom[16800] = 25'b1111111101110111101100111;
    rom[16801] = 25'b1111111101110111011010010;
    rom[16802] = 25'b1111111101110111000111101;
    rom[16803] = 25'b1111111101110110110101000;
    rom[16804] = 25'b1111111101110110100010011;
    rom[16805] = 25'b1111111101110110001111110;
    rom[16806] = 25'b1111111101110101111101000;
    rom[16807] = 25'b1111111101110101101010100;
    rom[16808] = 25'b1111111101110101010111110;
    rom[16809] = 25'b1111111101110101000101010;
    rom[16810] = 25'b1111111101110100110010100;
    rom[16811] = 25'b1111111101110100100000000;
    rom[16812] = 25'b1111111101110100001101011;
    rom[16813] = 25'b1111111101110011111010110;
    rom[16814] = 25'b1111111101110011101000001;
    rom[16815] = 25'b1111111101110011010101100;
    rom[16816] = 25'b1111111101110011000010111;
    rom[16817] = 25'b1111111101110010110000010;
    rom[16818] = 25'b1111111101110010011101101;
    rom[16819] = 25'b1111111101110010001011001;
    rom[16820] = 25'b1111111101110001111000011;
    rom[16821] = 25'b1111111101110001100101111;
    rom[16822] = 25'b1111111101110001010011010;
    rom[16823] = 25'b1111111101110001000000101;
    rom[16824] = 25'b1111111101110000101110001;
    rom[16825] = 25'b1111111101110000011011100;
    rom[16826] = 25'b1111111101110000001000111;
    rom[16827] = 25'b1111111101101111110110011;
    rom[16828] = 25'b1111111101101111100011110;
    rom[16829] = 25'b1111111101101111010001001;
    rom[16830] = 25'b1111111101101110111110101;
    rom[16831] = 25'b1111111101101110101100001;
    rom[16832] = 25'b1111111101101110011001100;
    rom[16833] = 25'b1111111101101110000110111;
    rom[16834] = 25'b1111111101101101110100011;
    rom[16835] = 25'b1111111101101101100001111;
    rom[16836] = 25'b1111111101101101001111010;
    rom[16837] = 25'b1111111101101100111100101;
    rom[16838] = 25'b1111111101101100101010001;
    rom[16839] = 25'b1111111101101100010111101;
    rom[16840] = 25'b1111111101101100000101001;
    rom[16841] = 25'b1111111101101011110010100;
    rom[16842] = 25'b1111111101101011100000000;
    rom[16843] = 25'b1111111101101011001101100;
    rom[16844] = 25'b1111111101101010111011000;
    rom[16845] = 25'b1111111101101010101000011;
    rom[16846] = 25'b1111111101101010010101111;
    rom[16847] = 25'b1111111101101010000011011;
    rom[16848] = 25'b1111111101101001110000111;
    rom[16849] = 25'b1111111101101001011110011;
    rom[16850] = 25'b1111111101101001001011111;
    rom[16851] = 25'b1111111101101000111001011;
    rom[16852] = 25'b1111111101101000100110111;
    rom[16853] = 25'b1111111101101000010100011;
    rom[16854] = 25'b1111111101101000000001111;
    rom[16855] = 25'b1111111101100111101111011;
    rom[16856] = 25'b1111111101100111011100111;
    rom[16857] = 25'b1111111101100111001010011;
    rom[16858] = 25'b1111111101100110110111111;
    rom[16859] = 25'b1111111101100110100101100;
    rom[16860] = 25'b1111111101100110010011000;
    rom[16861] = 25'b1111111101100110000000100;
    rom[16862] = 25'b1111111101100101101110000;
    rom[16863] = 25'b1111111101100101011011101;
    rom[16864] = 25'b1111111101100101001001001;
    rom[16865] = 25'b1111111101100100110110110;
    rom[16866] = 25'b1111111101100100100100010;
    rom[16867] = 25'b1111111101100100010001111;
    rom[16868] = 25'b1111111101100011111111011;
    rom[16869] = 25'b1111111101100011101101000;
    rom[16870] = 25'b1111111101100011011010101;
    rom[16871] = 25'b1111111101100011001000001;
    rom[16872] = 25'b1111111101100010110101110;
    rom[16873] = 25'b1111111101100010100011010;
    rom[16874] = 25'b1111111101100010010000111;
    rom[16875] = 25'b1111111101100001111110100;
    rom[16876] = 25'b1111111101100001101100000;
    rom[16877] = 25'b1111111101100001011001101;
    rom[16878] = 25'b1111111101100001000111010;
    rom[16879] = 25'b1111111101100000110100111;
    rom[16880] = 25'b1111111101100000100010100;
    rom[16881] = 25'b1111111101100000010000001;
    rom[16882] = 25'b1111111101011111111101110;
    rom[16883] = 25'b1111111101011111101011011;
    rom[16884] = 25'b1111111101011111011001000;
    rom[16885] = 25'b1111111101011111000110101;
    rom[16886] = 25'b1111111101011110110100010;
    rom[16887] = 25'b1111111101011110100001111;
    rom[16888] = 25'b1111111101011110001111100;
    rom[16889] = 25'b1111111101011101111101010;
    rom[16890] = 25'b1111111101011101101010111;
    rom[16891] = 25'b1111111101011101011000100;
    rom[16892] = 25'b1111111101011101000110010;
    rom[16893] = 25'b1111111101011100110011111;
    rom[16894] = 25'b1111111101011100100001100;
    rom[16895] = 25'b1111111101011100001111010;
    rom[16896] = 25'b1111111101011011111100111;
    rom[16897] = 25'b1111111101011011101010101;
    rom[16898] = 25'b1111111101011011011000010;
    rom[16899] = 25'b1111111101011011000110000;
    rom[16900] = 25'b1111111101011010110011101;
    rom[16901] = 25'b1111111101011010100001100;
    rom[16902] = 25'b1111111101011010001111001;
    rom[16903] = 25'b1111111101011001111100111;
    rom[16904] = 25'b1111111101011001101010101;
    rom[16905] = 25'b1111111101011001011000011;
    rom[16906] = 25'b1111111101011001000110000;
    rom[16907] = 25'b1111111101011000110011111;
    rom[16908] = 25'b1111111101011000100001100;
    rom[16909] = 25'b1111111101011000001111011;
    rom[16910] = 25'b1111111101010111111101001;
    rom[16911] = 25'b1111111101010111101010110;
    rom[16912] = 25'b1111111101010111011000101;
    rom[16913] = 25'b1111111101010111000110011;
    rom[16914] = 25'b1111111101010110110100001;
    rom[16915] = 25'b1111111101010110100010000;
    rom[16916] = 25'b1111111101010110001111110;
    rom[16917] = 25'b1111111101010101111101100;
    rom[16918] = 25'b1111111101010101101011011;
    rom[16919] = 25'b1111111101010101011001001;
    rom[16920] = 25'b1111111101010101000110111;
    rom[16921] = 25'b1111111101010100110100110;
    rom[16922] = 25'b1111111101010100100010101;
    rom[16923] = 25'b1111111101010100010000011;
    rom[16924] = 25'b1111111101010011111110010;
    rom[16925] = 25'b1111111101010011101100001;
    rom[16926] = 25'b1111111101010011011001111;
    rom[16927] = 25'b1111111101010011000111111;
    rom[16928] = 25'b1111111101010010110101110;
    rom[16929] = 25'b1111111101010010100011100;
    rom[16930] = 25'b1111111101010010010001011;
    rom[16931] = 25'b1111111101010001111111010;
    rom[16932] = 25'b1111111101010001101101001;
    rom[16933] = 25'b1111111101010001011011000;
    rom[16934] = 25'b1111111101010001001000111;
    rom[16935] = 25'b1111111101010000110110110;
    rom[16936] = 25'b1111111101010000100100110;
    rom[16937] = 25'b1111111101010000010010101;
    rom[16938] = 25'b1111111101010000000000100;
    rom[16939] = 25'b1111111101001111101110100;
    rom[16940] = 25'b1111111101001111011100011;
    rom[16941] = 25'b1111111101001111001010011;
    rom[16942] = 25'b1111111101001110111000010;
    rom[16943] = 25'b1111111101001110100110010;
    rom[16944] = 25'b1111111101001110010100010;
    rom[16945] = 25'b1111111101001110000010001;
    rom[16946] = 25'b1111111101001101110000001;
    rom[16947] = 25'b1111111101001101011110001;
    rom[16948] = 25'b1111111101001101001100001;
    rom[16949] = 25'b1111111101001100111010001;
    rom[16950] = 25'b1111111101001100101000000;
    rom[16951] = 25'b1111111101001100010110000;
    rom[16952] = 25'b1111111101001100000100000;
    rom[16953] = 25'b1111111101001011110010001;
    rom[16954] = 25'b1111111101001011100000000;
    rom[16955] = 25'b1111111101001011001110001;
    rom[16956] = 25'b1111111101001010111100001;
    rom[16957] = 25'b1111111101001010101010001;
    rom[16958] = 25'b1111111101001010011000010;
    rom[16959] = 25'b1111111101001010000110010;
    rom[16960] = 25'b1111111101001001110100010;
    rom[16961] = 25'b1111111101001001100010011;
    rom[16962] = 25'b1111111101001001010000011;
    rom[16963] = 25'b1111111101001000111110100;
    rom[16964] = 25'b1111111101001000101100101;
    rom[16965] = 25'b1111111101001000011010110;
    rom[16966] = 25'b1111111101001000001000110;
    rom[16967] = 25'b1111111101000111110110111;
    rom[16968] = 25'b1111111101000111100101000;
    rom[16969] = 25'b1111111101000111010011001;
    rom[16970] = 25'b1111111101000111000001010;
    rom[16971] = 25'b1111111101000110101111011;
    rom[16972] = 25'b1111111101000110011101100;
    rom[16973] = 25'b1111111101000110001011101;
    rom[16974] = 25'b1111111101000101111001111;
    rom[16975] = 25'b1111111101000101101000000;
    rom[16976] = 25'b1111111101000101010110001;
    rom[16977] = 25'b1111111101000101000100011;
    rom[16978] = 25'b1111111101000100110010100;
    rom[16979] = 25'b1111111101000100100000110;
    rom[16980] = 25'b1111111101000100001110111;
    rom[16981] = 25'b1111111101000011111101000;
    rom[16982] = 25'b1111111101000011101011011;
    rom[16983] = 25'b1111111101000011011001101;
    rom[16984] = 25'b1111111101000011000111110;
    rom[16985] = 25'b1111111101000010110110000;
    rom[16986] = 25'b1111111101000010100100010;
    rom[16987] = 25'b1111111101000010010010100;
    rom[16988] = 25'b1111111101000010000000110;
    rom[16989] = 25'b1111111101000001101111000;
    rom[16990] = 25'b1111111101000001011101010;
    rom[16991] = 25'b1111111101000001001011100;
    rom[16992] = 25'b1111111101000000111001110;
    rom[16993] = 25'b1111111101000000101000001;
    rom[16994] = 25'b1111111101000000010110011;
    rom[16995] = 25'b1111111101000000000100110;
    rom[16996] = 25'b1111111100111111110011001;
    rom[16997] = 25'b1111111100111111100001011;
    rom[16998] = 25'b1111111100111111001111110;
    rom[16999] = 25'b1111111100111110111110000;
    rom[17000] = 25'b1111111100111110101100011;
    rom[17001] = 25'b1111111100111110011010110;
    rom[17002] = 25'b1111111100111110001001001;
    rom[17003] = 25'b1111111100111101110111100;
    rom[17004] = 25'b1111111100111101100101111;
    rom[17005] = 25'b1111111100111101010100010;
    rom[17006] = 25'b1111111100111101000010101;
    rom[17007] = 25'b1111111100111100110001000;
    rom[17008] = 25'b1111111100111100011111100;
    rom[17009] = 25'b1111111100111100001101111;
    rom[17010] = 25'b1111111100111011111100010;
    rom[17011] = 25'b1111111100111011101010110;
    rom[17012] = 25'b1111111100111011011001001;
    rom[17013] = 25'b1111111100111011000111101;
    rom[17014] = 25'b1111111100111010110110001;
    rom[17015] = 25'b1111111100111010100100101;
    rom[17016] = 25'b1111111100111010010011000;
    rom[17017] = 25'b1111111100111010000001100;
    rom[17018] = 25'b1111111100111001110000000;
    rom[17019] = 25'b1111111100111001011110100;
    rom[17020] = 25'b1111111100111001001101000;
    rom[17021] = 25'b1111111100111000111011100;
    rom[17022] = 25'b1111111100111000101010000;
    rom[17023] = 25'b1111111100111000011000101;
    rom[17024] = 25'b1111111100111000000111001;
    rom[17025] = 25'b1111111100110111110101101;
    rom[17026] = 25'b1111111100110111100100010;
    rom[17027] = 25'b1111111100110111010010111;
    rom[17028] = 25'b1111111100110111000001011;
    rom[17029] = 25'b1111111100110110110000000;
    rom[17030] = 25'b1111111100110110011110101;
    rom[17031] = 25'b1111111100110110001101001;
    rom[17032] = 25'b1111111100110101111011110;
    rom[17033] = 25'b1111111100110101101010011;
    rom[17034] = 25'b1111111100110101011001000;
    rom[17035] = 25'b1111111100110101000111101;
    rom[17036] = 25'b1111111100110100110110011;
    rom[17037] = 25'b1111111100110100100101000;
    rom[17038] = 25'b1111111100110100010011101;
    rom[17039] = 25'b1111111100110100000010011;
    rom[17040] = 25'b1111111100110011110001000;
    rom[17041] = 25'b1111111100110011011111110;
    rom[17042] = 25'b1111111100110011001110100;
    rom[17043] = 25'b1111111100110010111101001;
    rom[17044] = 25'b1111111100110010101011111;
    rom[17045] = 25'b1111111100110010011010101;
    rom[17046] = 25'b1111111100110010001001011;
    rom[17047] = 25'b1111111100110001111000001;
    rom[17048] = 25'b1111111100110001100110110;
    rom[17049] = 25'b1111111100110001010101101;
    rom[17050] = 25'b1111111100110001000100011;
    rom[17051] = 25'b1111111100110000110011001;
    rom[17052] = 25'b1111111100110000100010000;
    rom[17053] = 25'b1111111100110000010000110;
    rom[17054] = 25'b1111111100101111111111101;
    rom[17055] = 25'b1111111100101111101110011;
    rom[17056] = 25'b1111111100101111011101010;
    rom[17057] = 25'b1111111100101111001100001;
    rom[17058] = 25'b1111111100101110111010111;
    rom[17059] = 25'b1111111100101110101001110;
    rom[17060] = 25'b1111111100101110011000101;
    rom[17061] = 25'b1111111100101110000111100;
    rom[17062] = 25'b1111111100101101110110011;
    rom[17063] = 25'b1111111100101101100101011;
    rom[17064] = 25'b1111111100101101010100010;
    rom[17065] = 25'b1111111100101101000011001;
    rom[17066] = 25'b1111111100101100110010001;
    rom[17067] = 25'b1111111100101100100001000;
    rom[17068] = 25'b1111111100101100010000000;
    rom[17069] = 25'b1111111100101011111110111;
    rom[17070] = 25'b1111111100101011101101111;
    rom[17071] = 25'b1111111100101011011100111;
    rom[17072] = 25'b1111111100101011001011111;
    rom[17073] = 25'b1111111100101010111010111;
    rom[17074] = 25'b1111111100101010101001111;
    rom[17075] = 25'b1111111100101010011000111;
    rom[17076] = 25'b1111111100101010000111111;
    rom[17077] = 25'b1111111100101001110110111;
    rom[17078] = 25'b1111111100101001100110000;
    rom[17079] = 25'b1111111100101001010101000;
    rom[17080] = 25'b1111111100101001000100001;
    rom[17081] = 25'b1111111100101000110011010;
    rom[17082] = 25'b1111111100101000100010011;
    rom[17083] = 25'b1111111100101000010001011;
    rom[17084] = 25'b1111111100101000000000100;
    rom[17085] = 25'b1111111100100111101111101;
    rom[17086] = 25'b1111111100100111011110110;
    rom[17087] = 25'b1111111100100111001101111;
    rom[17088] = 25'b1111111100100110111101000;
    rom[17089] = 25'b1111111100100110101100001;
    rom[17090] = 25'b1111111100100110011011011;
    rom[17091] = 25'b1111111100100110001010101;
    rom[17092] = 25'b1111111100100101111001110;
    rom[17093] = 25'b1111111100100101101001000;
    rom[17094] = 25'b1111111100100101011000001;
    rom[17095] = 25'b1111111100100101000111011;
    rom[17096] = 25'b1111111100100100110110101;
    rom[17097] = 25'b1111111100100100100101111;
    rom[17098] = 25'b1111111100100100010101001;
    rom[17099] = 25'b1111111100100100000100011;
    rom[17100] = 25'b1111111100100011110011101;
    rom[17101] = 25'b1111111100100011100010111;
    rom[17102] = 25'b1111111100100011010010010;
    rom[17103] = 25'b1111111100100011000001100;
    rom[17104] = 25'b1111111100100010110000111;
    rom[17105] = 25'b1111111100100010100000001;
    rom[17106] = 25'b1111111100100010001111100;
    rom[17107] = 25'b1111111100100001111110111;
    rom[17108] = 25'b1111111100100001101110010;
    rom[17109] = 25'b1111111100100001011101101;
    rom[17110] = 25'b1111111100100001001101000;
    rom[17111] = 25'b1111111100100000111100011;
    rom[17112] = 25'b1111111100100000101011110;
    rom[17113] = 25'b1111111100100000011011010;
    rom[17114] = 25'b1111111100100000001010101;
    rom[17115] = 25'b1111111100011111111010001;
    rom[17116] = 25'b1111111100011111101001101;
    rom[17117] = 25'b1111111100011111011001000;
    rom[17118] = 25'b1111111100011111001000100;
    rom[17119] = 25'b1111111100011110111000000;
    rom[17120] = 25'b1111111100011110100111100;
    rom[17121] = 25'b1111111100011110010111000;
    rom[17122] = 25'b1111111100011110000110100;
    rom[17123] = 25'b1111111100011101110110001;
    rom[17124] = 25'b1111111100011101100101101;
    rom[17125] = 25'b1111111100011101010101001;
    rom[17126] = 25'b1111111100011101000100101;
    rom[17127] = 25'b1111111100011100110100011;
    rom[17128] = 25'b1111111100011100100011111;
    rom[17129] = 25'b1111111100011100010011100;
    rom[17130] = 25'b1111111100011100000011001;
    rom[17131] = 25'b1111111100011011110010101;
    rom[17132] = 25'b1111111100011011100010011;
    rom[17133] = 25'b1111111100011011010010000;
    rom[17134] = 25'b1111111100011011000001101;
    rom[17135] = 25'b1111111100011010110001010;
    rom[17136] = 25'b1111111100011010100001000;
    rom[17137] = 25'b1111111100011010010000110;
    rom[17138] = 25'b1111111100011010000000100;
    rom[17139] = 25'b1111111100011001110000001;
    rom[17140] = 25'b1111111100011001011111111;
    rom[17141] = 25'b1111111100011001001111101;
    rom[17142] = 25'b1111111100011000111111011;
    rom[17143] = 25'b1111111100011000101111001;
    rom[17144] = 25'b1111111100011000011110111;
    rom[17145] = 25'b1111111100011000001110110;
    rom[17146] = 25'b1111111100010111111110100;
    rom[17147] = 25'b1111111100010111101110010;
    rom[17148] = 25'b1111111100010111011110001;
    rom[17149] = 25'b1111111100010111001110000;
    rom[17150] = 25'b1111111100010110111101111;
    rom[17151] = 25'b1111111100010110101101110;
    rom[17152] = 25'b1111111100010110011101100;
    rom[17153] = 25'b1111111100010110001101100;
    rom[17154] = 25'b1111111100010101111101011;
    rom[17155] = 25'b1111111100010101101101010;
    rom[17156] = 25'b1111111100010101011101010;
    rom[17157] = 25'b1111111100010101001101001;
    rom[17158] = 25'b1111111100010100111101001;
    rom[17159] = 25'b1111111100010100101101001;
    rom[17160] = 25'b1111111100010100011101000;
    rom[17161] = 25'b1111111100010100001101000;
    rom[17162] = 25'b1111111100010011111101000;
    rom[17163] = 25'b1111111100010011101101000;
    rom[17164] = 25'b1111111100010011011101000;
    rom[17165] = 25'b1111111100010011001101001;
    rom[17166] = 25'b1111111100010010111101001;
    rom[17167] = 25'b1111111100010010101101001;
    rom[17168] = 25'b1111111100010010011101010;
    rom[17169] = 25'b1111111100010010001101011;
    rom[17170] = 25'b1111111100010001111101011;
    rom[17171] = 25'b1111111100010001101101100;
    rom[17172] = 25'b1111111100010001011101101;
    rom[17173] = 25'b1111111100010001001101110;
    rom[17174] = 25'b1111111100010000111110000;
    rom[17175] = 25'b1111111100010000101110001;
    rom[17176] = 25'b1111111100010000011110011;
    rom[17177] = 25'b1111111100010000001110100;
    rom[17178] = 25'b1111111100001111111110110;
    rom[17179] = 25'b1111111100001111101110111;
    rom[17180] = 25'b1111111100001111011111001;
    rom[17181] = 25'b1111111100001111001111100;
    rom[17182] = 25'b1111111100001110111111101;
    rom[17183] = 25'b1111111100001110110000000;
    rom[17184] = 25'b1111111100001110100000010;
    rom[17185] = 25'b1111111100001110010000100;
    rom[17186] = 25'b1111111100001110000000111;
    rom[17187] = 25'b1111111100001101110001001;
    rom[17188] = 25'b1111111100001101100001100;
    rom[17189] = 25'b1111111100001101010001111;
    rom[17190] = 25'b1111111100001101000010010;
    rom[17191] = 25'b1111111100001100110010101;
    rom[17192] = 25'b1111111100001100100011000;
    rom[17193] = 25'b1111111100001100010011011;
    rom[17194] = 25'b1111111100001100000011110;
    rom[17195] = 25'b1111111100001011110100010;
    rom[17196] = 25'b1111111100001011100100101;
    rom[17197] = 25'b1111111100001011010101001;
    rom[17198] = 25'b1111111100001011000101101;
    rom[17199] = 25'b1111111100001010110110001;
    rom[17200] = 25'b1111111100001010100110101;
    rom[17201] = 25'b1111111100001010010111001;
    rom[17202] = 25'b1111111100001010000111101;
    rom[17203] = 25'b1111111100001001111000001;
    rom[17204] = 25'b1111111100001001101000110;
    rom[17205] = 25'b1111111100001001011001010;
    rom[17206] = 25'b1111111100001001001001111;
    rom[17207] = 25'b1111111100001000111010011;
    rom[17208] = 25'b1111111100001000101011000;
    rom[17209] = 25'b1111111100001000011011110;
    rom[17210] = 25'b1111111100001000001100010;
    rom[17211] = 25'b1111111100000111111101000;
    rom[17212] = 25'b1111111100000111101101101;
    rom[17213] = 25'b1111111100000111011110011;
    rom[17214] = 25'b1111111100000111001111000;
    rom[17215] = 25'b1111111100000110111111110;
    rom[17216] = 25'b1111111100000110110000011;
    rom[17217] = 25'b1111111100000110100001001;
    rom[17218] = 25'b1111111100000110010010000;
    rom[17219] = 25'b1111111100000110000010101;
    rom[17220] = 25'b1111111100000101110011011;
    rom[17221] = 25'b1111111100000101100100010;
    rom[17222] = 25'b1111111100000101010101001;
    rom[17223] = 25'b1111111100000101000101111;
    rom[17224] = 25'b1111111100000100110110110;
    rom[17225] = 25'b1111111100000100100111101;
    rom[17226] = 25'b1111111100000100011000100;
    rom[17227] = 25'b1111111100000100001001011;
    rom[17228] = 25'b1111111100000011111010010;
    rom[17229] = 25'b1111111100000011101011001;
    rom[17230] = 25'b1111111100000011011100000;
    rom[17231] = 25'b1111111100000011001100111;
    rom[17232] = 25'b1111111100000010111101111;
    rom[17233] = 25'b1111111100000010101110111;
    rom[17234] = 25'b1111111100000010011111110;
    rom[17235] = 25'b1111111100000010010000111;
    rom[17236] = 25'b1111111100000010000001111;
    rom[17237] = 25'b1111111100000001110010111;
    rom[17238] = 25'b1111111100000001100100000;
    rom[17239] = 25'b1111111100000001010101000;
    rom[17240] = 25'b1111111100000001000110001;
    rom[17241] = 25'b1111111100000000110111001;
    rom[17242] = 25'b1111111100000000101000001;
    rom[17243] = 25'b1111111100000000011001011;
    rom[17244] = 25'b1111111100000000001010100;
    rom[17245] = 25'b1111111011111111111011101;
    rom[17246] = 25'b1111111011111111101100110;
    rom[17247] = 25'b1111111011111111011110000;
    rom[17248] = 25'b1111111011111111001111001;
    rom[17249] = 25'b1111111011111111000000011;
    rom[17250] = 25'b1111111011111110110001101;
    rom[17251] = 25'b1111111011111110100010110;
    rom[17252] = 25'b1111111011111110010100000;
    rom[17253] = 25'b1111111011111110000101011;
    rom[17254] = 25'b1111111011111101110110100;
    rom[17255] = 25'b1111111011111101100111111;
    rom[17256] = 25'b1111111011111101011001001;
    rom[17257] = 25'b1111111011111101001010100;
    rom[17258] = 25'b1111111011111100111011111;
    rom[17259] = 25'b1111111011111100101101001;
    rom[17260] = 25'b1111111011111100011110101;
    rom[17261] = 25'b1111111011111100001111111;
    rom[17262] = 25'b1111111011111100000001011;
    rom[17263] = 25'b1111111011111011110010110;
    rom[17264] = 25'b1111111011111011100100010;
    rom[17265] = 25'b1111111011111011010101101;
    rom[17266] = 25'b1111111011111011000111001;
    rom[17267] = 25'b1111111011111010111000101;
    rom[17268] = 25'b1111111011111010101010000;
    rom[17269] = 25'b1111111011111010011011101;
    rom[17270] = 25'b1111111011111010001101001;
    rom[17271] = 25'b1111111011111001111110101;
    rom[17272] = 25'b1111111011111001110000010;
    rom[17273] = 25'b1111111011111001100001110;
    rom[17274] = 25'b1111111011111001010011011;
    rom[17275] = 25'b1111111011111001000101000;
    rom[17276] = 25'b1111111011111000110110101;
    rom[17277] = 25'b1111111011111000101000010;
    rom[17278] = 25'b1111111011111000011001111;
    rom[17279] = 25'b1111111011111000001011101;
    rom[17280] = 25'b1111111011110111111101001;
    rom[17281] = 25'b1111111011110111101110111;
    rom[17282] = 25'b1111111011110111100000101;
    rom[17283] = 25'b1111111011110111010010011;
    rom[17284] = 25'b1111111011110111000100001;
    rom[17285] = 25'b1111111011110110110101111;
    rom[17286] = 25'b1111111011110110100111101;
    rom[17287] = 25'b1111111011110110011001100;
    rom[17288] = 25'b1111111011110110001011010;
    rom[17289] = 25'b1111111011110101111101001;
    rom[17290] = 25'b1111111011110101101111000;
    rom[17291] = 25'b1111111011110101100000111;
    rom[17292] = 25'b1111111011110101010010101;
    rom[17293] = 25'b1111111011110101000100100;
    rom[17294] = 25'b1111111011110100110110100;
    rom[17295] = 25'b1111111011110100101000100;
    rom[17296] = 25'b1111111011110100011010011;
    rom[17297] = 25'b1111111011110100001100011;
    rom[17298] = 25'b1111111011110011111110011;
    rom[17299] = 25'b1111111011110011110000011;
    rom[17300] = 25'b1111111011110011100010011;
    rom[17301] = 25'b1111111011110011010100010;
    rom[17302] = 25'b1111111011110011000110011;
    rom[17303] = 25'b1111111011110010111000011;
    rom[17304] = 25'b1111111011110010101010100;
    rom[17305] = 25'b1111111011110010011100100;
    rom[17306] = 25'b1111111011110010001110110;
    rom[17307] = 25'b1111111011110010000000111;
    rom[17308] = 25'b1111111011110001110011000;
    rom[17309] = 25'b1111111011110001100101001;
    rom[17310] = 25'b1111111011110001010111010;
    rom[17311] = 25'b1111111011110001001001100;
    rom[17312] = 25'b1111111011110000111011110;
    rom[17313] = 25'b1111111011110000101101111;
    rom[17314] = 25'b1111111011110000100000001;
    rom[17315] = 25'b1111111011110000010010011;
    rom[17316] = 25'b1111111011110000000100110;
    rom[17317] = 25'b1111111011101111110111000;
    rom[17318] = 25'b1111111011101111101001011;
    rom[17319] = 25'b1111111011101111011011101;
    rom[17320] = 25'b1111111011101111001110000;
    rom[17321] = 25'b1111111011101111000000011;
    rom[17322] = 25'b1111111011101110110010110;
    rom[17323] = 25'b1111111011101110100101001;
    rom[17324] = 25'b1111111011101110010111100;
    rom[17325] = 25'b1111111011101110001010000;
    rom[17326] = 25'b1111111011101101111100100;
    rom[17327] = 25'b1111111011101101101110111;
    rom[17328] = 25'b1111111011101101100001011;
    rom[17329] = 25'b1111111011101101010011111;
    rom[17330] = 25'b1111111011101101000110011;
    rom[17331] = 25'b1111111011101100111000111;
    rom[17332] = 25'b1111111011101100101011100;
    rom[17333] = 25'b1111111011101100011110000;
    rom[17334] = 25'b1111111011101100010000101;
    rom[17335] = 25'b1111111011101100000011010;
    rom[17336] = 25'b1111111011101011110101111;
    rom[17337] = 25'b1111111011101011101000100;
    rom[17338] = 25'b1111111011101011011011001;
    rom[17339] = 25'b1111111011101011001101111;
    rom[17340] = 25'b1111111011101011000000100;
    rom[17341] = 25'b1111111011101010110011010;
    rom[17342] = 25'b1111111011101010100110000;
    rom[17343] = 25'b1111111011101010011000101;
    rom[17344] = 25'b1111111011101010001011011;
    rom[17345] = 25'b1111111011101001111110010;
    rom[17346] = 25'b1111111011101001110001001;
    rom[17347] = 25'b1111111011101001100011111;
    rom[17348] = 25'b1111111011101001010110101;
    rom[17349] = 25'b1111111011101001001001101;
    rom[17350] = 25'b1111111011101000111100011;
    rom[17351] = 25'b1111111011101000101111011;
    rom[17352] = 25'b1111111011101000100010001;
    rom[17353] = 25'b1111111011101000010101001;
    rom[17354] = 25'b1111111011101000001000001;
    rom[17355] = 25'b1111111011100111111011000;
    rom[17356] = 25'b1111111011100111101110000;
    rom[17357] = 25'b1111111011100111100001000;
    rom[17358] = 25'b1111111011100111010100000;
    rom[17359] = 25'b1111111011100111000111000;
    rom[17360] = 25'b1111111011100110111010001;
    rom[17361] = 25'b1111111011100110101101001;
    rom[17362] = 25'b1111111011100110100000010;
    rom[17363] = 25'b1111111011100110010011011;
    rom[17364] = 25'b1111111011100110000110100;
    rom[17365] = 25'b1111111011100101111001101;
    rom[17366] = 25'b1111111011100101101100111;
    rom[17367] = 25'b1111111011100101100000000;
    rom[17368] = 25'b1111111011100101010011010;
    rom[17369] = 25'b1111111011100101000110011;
    rom[17370] = 25'b1111111011100100111001101;
    rom[17371] = 25'b1111111011100100101100111;
    rom[17372] = 25'b1111111011100100100000001;
    rom[17373] = 25'b1111111011100100010011100;
    rom[17374] = 25'b1111111011100100000110110;
    rom[17375] = 25'b1111111011100011111010000;
    rom[17376] = 25'b1111111011100011101101100;
    rom[17377] = 25'b1111111011100011100000111;
    rom[17378] = 25'b1111111011100011010100010;
    rom[17379] = 25'b1111111011100011000111101;
    rom[17380] = 25'b1111111011100010111011000;
    rom[17381] = 25'b1111111011100010101110011;
    rom[17382] = 25'b1111111011100010100001111;
    rom[17383] = 25'b1111111011100010010101011;
    rom[17384] = 25'b1111111011100010001000111;
    rom[17385] = 25'b1111111011100001111100100;
    rom[17386] = 25'b1111111011100001101111111;
    rom[17387] = 25'b1111111011100001100011100;
    rom[17388] = 25'b1111111011100001010111001;
    rom[17389] = 25'b1111111011100001001010101;
    rom[17390] = 25'b1111111011100000111110010;
    rom[17391] = 25'b1111111011100000110001111;
    rom[17392] = 25'b1111111011100000100101100;
    rom[17393] = 25'b1111111011100000011001001;
    rom[17394] = 25'b1111111011100000001100111;
    rom[17395] = 25'b1111111011100000000000101;
    rom[17396] = 25'b1111111011011111110100010;
    rom[17397] = 25'b1111111011011111101000000;
    rom[17398] = 25'b1111111011011111011011111;
    rom[17399] = 25'b1111111011011111001111101;
    rom[17400] = 25'b1111111011011111000011100;
    rom[17401] = 25'b1111111011011110110111010;
    rom[17402] = 25'b1111111011011110101011001;
    rom[17403] = 25'b1111111011011110011110111;
    rom[17404] = 25'b1111111011011110010010110;
    rom[17405] = 25'b1111111011011110000110110;
    rom[17406] = 25'b1111111011011101111010101;
    rom[17407] = 25'b1111111011011101101110100;
    rom[17408] = 25'b1111111011011101100010100;
    rom[17409] = 25'b1111111011011101010110100;
    rom[17410] = 25'b1111111011011101001010100;
    rom[17411] = 25'b1111111011011100111110100;
    rom[17412] = 25'b1111111011011100110010101;
    rom[17413] = 25'b1111111011011100100110101;
    rom[17414] = 25'b1111111011011100011010110;
    rom[17415] = 25'b1111111011011100001110110;
    rom[17416] = 25'b1111111011011100000010111;
    rom[17417] = 25'b1111111011011011110111000;
    rom[17418] = 25'b1111111011011011101011001;
    rom[17419] = 25'b1111111011011011011111011;
    rom[17420] = 25'b1111111011011011010011100;
    rom[17421] = 25'b1111111011011011000111110;
    rom[17422] = 25'b1111111011011010111100000;
    rom[17423] = 25'b1111111011011010110000010;
    rom[17424] = 25'b1111111011011010100100100;
    rom[17425] = 25'b1111111011011010011000110;
    rom[17426] = 25'b1111111011011010001101001;
    rom[17427] = 25'b1111111011011010000001100;
    rom[17428] = 25'b1111111011011001110101111;
    rom[17429] = 25'b1111111011011001101010010;
    rom[17430] = 25'b1111111011011001011110101;
    rom[17431] = 25'b1111111011011001010011000;
    rom[17432] = 25'b1111111011011001000111100;
    rom[17433] = 25'b1111111011011000111011111;
    rom[17434] = 25'b1111111011011000110000011;
    rom[17435] = 25'b1111111011011000100100111;
    rom[17436] = 25'b1111111011011000011001011;
    rom[17437] = 25'b1111111011011000001101111;
    rom[17438] = 25'b1111111011011000000010011;
    rom[17439] = 25'b1111111011010111110111000;
    rom[17440] = 25'b1111111011010111101011101;
    rom[17441] = 25'b1111111011010111100000010;
    rom[17442] = 25'b1111111011010111010100111;
    rom[17443] = 25'b1111111011010111001001101;
    rom[17444] = 25'b1111111011010110111110010;
    rom[17445] = 25'b1111111011010110110011000;
    rom[17446] = 25'b1111111011010110100111101;
    rom[17447] = 25'b1111111011010110011100011;
    rom[17448] = 25'b1111111011010110010001001;
    rom[17449] = 25'b1111111011010110000110000;
    rom[17450] = 25'b1111111011010101111010110;
    rom[17451] = 25'b1111111011010101101111100;
    rom[17452] = 25'b1111111011010101100100011;
    rom[17453] = 25'b1111111011010101011001010;
    rom[17454] = 25'b1111111011010101001110001;
    rom[17455] = 25'b1111111011010101000011001;
    rom[17456] = 25'b1111111011010100111000000;
    rom[17457] = 25'b1111111011010100101101000;
    rom[17458] = 25'b1111111011010100100001111;
    rom[17459] = 25'b1111111011010100010110111;
    rom[17460] = 25'b1111111011010100001011111;
    rom[17461] = 25'b1111111011010100000000111;
    rom[17462] = 25'b1111111011010011110110000;
    rom[17463] = 25'b1111111011010011101011000;
    rom[17464] = 25'b1111111011010011100000001;
    rom[17465] = 25'b1111111011010011010101010;
    rom[17466] = 25'b1111111011010011001010011;
    rom[17467] = 25'b1111111011010010111111100;
    rom[17468] = 25'b1111111011010010110100101;
    rom[17469] = 25'b1111111011010010101001111;
    rom[17470] = 25'b1111111011010010011111001;
    rom[17471] = 25'b1111111011010010010100011;
    rom[17472] = 25'b1111111011010010001001101;
    rom[17473] = 25'b1111111011010001111110111;
    rom[17474] = 25'b1111111011010001110100010;
    rom[17475] = 25'b1111111011010001101001101;
    rom[17476] = 25'b1111111011010001011110111;
    rom[17477] = 25'b1111111011010001010100010;
    rom[17478] = 25'b1111111011010001001001101;
    rom[17479] = 25'b1111111011010000111111001;
    rom[17480] = 25'b1111111011010000110100100;
    rom[17481] = 25'b1111111011010000101010000;
    rom[17482] = 25'b1111111011010000011111100;
    rom[17483] = 25'b1111111011010000010100111;
    rom[17484] = 25'b1111111011010000001010011;
    rom[17485] = 25'b1111111011010000000000000;
    rom[17486] = 25'b1111111011001111110101100;
    rom[17487] = 25'b1111111011001111101011001;
    rom[17488] = 25'b1111111011001111100000110;
    rom[17489] = 25'b1111111011001111010110011;
    rom[17490] = 25'b1111111011001111001100000;
    rom[17491] = 25'b1111111011001111000001101;
    rom[17492] = 25'b1111111011001110110111011;
    rom[17493] = 25'b1111111011001110101101001;
    rom[17494] = 25'b1111111011001110100010111;
    rom[17495] = 25'b1111111011001110011000101;
    rom[17496] = 25'b1111111011001110001110011;
    rom[17497] = 25'b1111111011001110000100001;
    rom[17498] = 25'b1111111011001101111010000;
    rom[17499] = 25'b1111111011001101101111111;
    rom[17500] = 25'b1111111011001101100101110;
    rom[17501] = 25'b1111111011001101011011101;
    rom[17502] = 25'b1111111011001101010001100;
    rom[17503] = 25'b1111111011001101000111011;
    rom[17504] = 25'b1111111011001100111101011;
    rom[17505] = 25'b1111111011001100110011011;
    rom[17506] = 25'b1111111011001100101001011;
    rom[17507] = 25'b1111111011001100011111011;
    rom[17508] = 25'b1111111011001100010101100;
    rom[17509] = 25'b1111111011001100001011100;
    rom[17510] = 25'b1111111011001100000001101;
    rom[17511] = 25'b1111111011001011110111101;
    rom[17512] = 25'b1111111011001011101101110;
    rom[17513] = 25'b1111111011001011100100000;
    rom[17514] = 25'b1111111011001011011010001;
    rom[17515] = 25'b1111111011001011010000011;
    rom[17516] = 25'b1111111011001011000110100;
    rom[17517] = 25'b1111111011001010111100111;
    rom[17518] = 25'b1111111011001010110011000;
    rom[17519] = 25'b1111111011001010101001011;
    rom[17520] = 25'b1111111011001010011111110;
    rom[17521] = 25'b1111111011001010010110000;
    rom[17522] = 25'b1111111011001010001100011;
    rom[17523] = 25'b1111111011001010000010110;
    rom[17524] = 25'b1111111011001001111001001;
    rom[17525] = 25'b1111111011001001101111101;
    rom[17526] = 25'b1111111011001001100110000;
    rom[17527] = 25'b1111111011001001011100100;
    rom[17528] = 25'b1111111011001001010011000;
    rom[17529] = 25'b1111111011001001001001100;
    rom[17530] = 25'b1111111011001001000000001;
    rom[17531] = 25'b1111111011001000110110100;
    rom[17532] = 25'b1111111011001000101101010;
    rom[17533] = 25'b1111111011001000100011110;
    rom[17534] = 25'b1111111011001000011010100;
    rom[17535] = 25'b1111111011001000010001001;
    rom[17536] = 25'b1111111011001000000111110;
    rom[17537] = 25'b1111111011000111111110011;
    rom[17538] = 25'b1111111011000111110101001;
    rom[17539] = 25'b1111111011000111101100000;
    rom[17540] = 25'b1111111011000111100010110;
    rom[17541] = 25'b1111111011000111011001100;
    rom[17542] = 25'b1111111011000111010000010;
    rom[17543] = 25'b1111111011000111000111001;
    rom[17544] = 25'b1111111011000110111110000;
    rom[17545] = 25'b1111111011000110110100111;
    rom[17546] = 25'b1111111011000110101011110;
    rom[17547] = 25'b1111111011000110100010101;
    rom[17548] = 25'b1111111011000110011001101;
    rom[17549] = 25'b1111111011000110010000101;
    rom[17550] = 25'b1111111011000110000111100;
    rom[17551] = 25'b1111111011000101111110101;
    rom[17552] = 25'b1111111011000101110101101;
    rom[17553] = 25'b1111111011000101101100110;
    rom[17554] = 25'b1111111011000101100011110;
    rom[17555] = 25'b1111111011000101011010111;
    rom[17556] = 25'b1111111011000101010010000;
    rom[17557] = 25'b1111111011000101001001010;
    rom[17558] = 25'b1111111011000101000000011;
    rom[17559] = 25'b1111111011000100110111101;
    rom[17560] = 25'b1111111011000100101110111;
    rom[17561] = 25'b1111111011000100100110000;
    rom[17562] = 25'b1111111011000100011101011;
    rom[17563] = 25'b1111111011000100010100101;
    rom[17564] = 25'b1111111011000100001100000;
    rom[17565] = 25'b1111111011000100000011011;
    rom[17566] = 25'b1111111011000011111010110;
    rom[17567] = 25'b1111111011000011110010001;
    rom[17568] = 25'b1111111011000011101001100;
    rom[17569] = 25'b1111111011000011100001000;
    rom[17570] = 25'b1111111011000011011000100;
    rom[17571] = 25'b1111111011000011010000000;
    rom[17572] = 25'b1111111011000011000111100;
    rom[17573] = 25'b1111111011000010111111000;
    rom[17574] = 25'b1111111011000010110110100;
    rom[17575] = 25'b1111111011000010101110001;
    rom[17576] = 25'b1111111011000010100101110;
    rom[17577] = 25'b1111111011000010011101011;
    rom[17578] = 25'b1111111011000010010101000;
    rom[17579] = 25'b1111111011000010001100110;
    rom[17580] = 25'b1111111011000010000100011;
    rom[17581] = 25'b1111111011000001111100001;
    rom[17582] = 25'b1111111011000001110011111;
    rom[17583] = 25'b1111111011000001101011101;
    rom[17584] = 25'b1111111011000001100011011;
    rom[17585] = 25'b1111111011000001011011010;
    rom[17586] = 25'b1111111011000001010011001;
    rom[17587] = 25'b1111111011000001001011000;
    rom[17588] = 25'b1111111011000001000010111;
    rom[17589] = 25'b1111111011000000111010110;
    rom[17590] = 25'b1111111011000000110010110;
    rom[17591] = 25'b1111111011000000101010110;
    rom[17592] = 25'b1111111011000000100010110;
    rom[17593] = 25'b1111111011000000011010110;
    rom[17594] = 25'b1111111011000000010010110;
    rom[17595] = 25'b1111111011000000001010111;
    rom[17596] = 25'b1111111011000000000011000;
    rom[17597] = 25'b1111111010111111111011000;
    rom[17598] = 25'b1111111010111111110011001;
    rom[17599] = 25'b1111111010111111101011011;
    rom[17600] = 25'b1111111010111111100011101;
    rom[17601] = 25'b1111111010111111011011110;
    rom[17602] = 25'b1111111010111111010100000;
    rom[17603] = 25'b1111111010111111001100010;
    rom[17604] = 25'b1111111010111111000100101;
    rom[17605] = 25'b1111111010111110111100111;
    rom[17606] = 25'b1111111010111110110101001;
    rom[17607] = 25'b1111111010111110101101100;
    rom[17608] = 25'b1111111010111110100110000;
    rom[17609] = 25'b1111111010111110011110011;
    rom[17610] = 25'b1111111010111110010110111;
    rom[17611] = 25'b1111111010111110001111010;
    rom[17612] = 25'b1111111010111110000111110;
    rom[17613] = 25'b1111111010111110000000010;
    rom[17614] = 25'b1111111010111101111000110;
    rom[17615] = 25'b1111111010111101110001010;
    rom[17616] = 25'b1111111010111101101001111;
    rom[17617] = 25'b1111111010111101100010100;
    rom[17618] = 25'b1111111010111101011011001;
    rom[17619] = 25'b1111111010111101010011110;
    rom[17620] = 25'b1111111010111101001100100;
    rom[17621] = 25'b1111111010111101000101010;
    rom[17622] = 25'b1111111010111100111101111;
    rom[17623] = 25'b1111111010111100110110101;
    rom[17624] = 25'b1111111010111100101111100;
    rom[17625] = 25'b1111111010111100101000010;
    rom[17626] = 25'b1111111010111100100001001;
    rom[17627] = 25'b1111111010111100011010000;
    rom[17628] = 25'b1111111010111100010010111;
    rom[17629] = 25'b1111111010111100001011110;
    rom[17630] = 25'b1111111010111100000100101;
    rom[17631] = 25'b1111111010111011111101101;
    rom[17632] = 25'b1111111010111011110110101;
    rom[17633] = 25'b1111111010111011101111101;
    rom[17634] = 25'b1111111010111011101000101;
    rom[17635] = 25'b1111111010111011100001110;
    rom[17636] = 25'b1111111010111011011010110;
    rom[17637] = 25'b1111111010111011010011111;
    rom[17638] = 25'b1111111010111011001101000;
    rom[17639] = 25'b1111111010111011000110010;
    rom[17640] = 25'b1111111010111010111111011;
    rom[17641] = 25'b1111111010111010111000101;
    rom[17642] = 25'b1111111010111010110001111;
    rom[17643] = 25'b1111111010111010101011001;
    rom[17644] = 25'b1111111010111010100100011;
    rom[17645] = 25'b1111111010111010011101101;
    rom[17646] = 25'b1111111010111010010111000;
    rom[17647] = 25'b1111111010111010010000011;
    rom[17648] = 25'b1111111010111010001001110;
    rom[17649] = 25'b1111111010111010000011001;
    rom[17650] = 25'b1111111010111001111100101;
    rom[17651] = 25'b1111111010111001110110001;
    rom[17652] = 25'b1111111010111001101111100;
    rom[17653] = 25'b1111111010111001101001001;
    rom[17654] = 25'b1111111010111001100010101;
    rom[17655] = 25'b1111111010111001011100010;
    rom[17656] = 25'b1111111010111001010101110;
    rom[17657] = 25'b1111111010111001001111011;
    rom[17658] = 25'b1111111010111001001001000;
    rom[17659] = 25'b1111111010111001000010110;
    rom[17660] = 25'b1111111010111000111100011;
    rom[17661] = 25'b1111111010111000110110001;
    rom[17662] = 25'b1111111010111000101111111;
    rom[17663] = 25'b1111111010111000101001101;
    rom[17664] = 25'b1111111010111000100011011;
    rom[17665] = 25'b1111111010111000011101010;
    rom[17666] = 25'b1111111010111000010111001;
    rom[17667] = 25'b1111111010111000010001000;
    rom[17668] = 25'b1111111010111000001010111;
    rom[17669] = 25'b1111111010111000000100110;
    rom[17670] = 25'b1111111010110111111110111;
    rom[17671] = 25'b1111111010110111111000110;
    rom[17672] = 25'b1111111010110111110010110;
    rom[17673] = 25'b1111111010110111101100110;
    rom[17674] = 25'b1111111010110111100110111;
    rom[17675] = 25'b1111111010110111100000111;
    rom[17676] = 25'b1111111010110111011011000;
    rom[17677] = 25'b1111111010110111010101001;
    rom[17678] = 25'b1111111010110111001111011;
    rom[17679] = 25'b1111111010110111001001100;
    rom[17680] = 25'b1111111010110111000011110;
    rom[17681] = 25'b1111111010110110111110000;
    rom[17682] = 25'b1111111010110110111000010;
    rom[17683] = 25'b1111111010110110110010100;
    rom[17684] = 25'b1111111010110110101100111;
    rom[17685] = 25'b1111111010110110100111010;
    rom[17686] = 25'b1111111010110110100001101;
    rom[17687] = 25'b1111111010110110011100000;
    rom[17688] = 25'b1111111010110110010110011;
    rom[17689] = 25'b1111111010110110010000111;
    rom[17690] = 25'b1111111010110110001011011;
    rom[17691] = 25'b1111111010110110000101111;
    rom[17692] = 25'b1111111010110110000000011;
    rom[17693] = 25'b1111111010110101111011000;
    rom[17694] = 25'b1111111010110101110101100;
    rom[17695] = 25'b1111111010110101110000001;
    rom[17696] = 25'b1111111010110101101010110;
    rom[17697] = 25'b1111111010110101100101100;
    rom[17698] = 25'b1111111010110101100000001;
    rom[17699] = 25'b1111111010110101011010111;
    rom[17700] = 25'b1111111010110101010101101;
    rom[17701] = 25'b1111111010110101010000011;
    rom[17702] = 25'b1111111010110101001011001;
    rom[17703] = 25'b1111111010110101000110000;
    rom[17704] = 25'b1111111010110101000000111;
    rom[17705] = 25'b1111111010110100111011110;
    rom[17706] = 25'b1111111010110100110110101;
    rom[17707] = 25'b1111111010110100110001100;
    rom[17708] = 25'b1111111010110100101100100;
    rom[17709] = 25'b1111111010110100100111100;
    rom[17710] = 25'b1111111010110100100010100;
    rom[17711] = 25'b1111111010110100011101101;
    rom[17712] = 25'b1111111010110100011000101;
    rom[17713] = 25'b1111111010110100010011110;
    rom[17714] = 25'b1111111010110100001110110;
    rom[17715] = 25'b1111111010110100001010000;
    rom[17716] = 25'b1111111010110100000101010;
    rom[17717] = 25'b1111111010110100000000011;
    rom[17718] = 25'b1111111010110011111011101;
    rom[17719] = 25'b1111111010110011110110110;
    rom[17720] = 25'b1111111010110011110010001;
    rom[17721] = 25'b1111111010110011101101100;
    rom[17722] = 25'b1111111010110011101000110;
    rom[17723] = 25'b1111111010110011100100001;
    rom[17724] = 25'b1111111010110011011111100;
    rom[17725] = 25'b1111111010110011011011000;
    rom[17726] = 25'b1111111010110011010110011;
    rom[17727] = 25'b1111111010110011010001111;
    rom[17728] = 25'b1111111010110011001101011;
    rom[17729] = 25'b1111111010110011001000111;
    rom[17730] = 25'b1111111010110011000100100;
    rom[17731] = 25'b1111111010110011000000000;
    rom[17732] = 25'b1111111010110010111011101;
    rom[17733] = 25'b1111111010110010110111010;
    rom[17734] = 25'b1111111010110010110010111;
    rom[17735] = 25'b1111111010110010101110101;
    rom[17736] = 25'b1111111010110010101010011;
    rom[17737] = 25'b1111111010110010100110001;
    rom[17738] = 25'b1111111010110010100001111;
    rom[17739] = 25'b1111111010110010011101101;
    rom[17740] = 25'b1111111010110010011001100;
    rom[17741] = 25'b1111111010110010010101011;
    rom[17742] = 25'b1111111010110010010001010;
    rom[17743] = 25'b1111111010110010001101001;
    rom[17744] = 25'b1111111010110010001001001;
    rom[17745] = 25'b1111111010110010000101001;
    rom[17746] = 25'b1111111010110010000001000;
    rom[17747] = 25'b1111111010110001111101000;
    rom[17748] = 25'b1111111010110001111001001;
    rom[17749] = 25'b1111111010110001110101010;
    rom[17750] = 25'b1111111010110001110001010;
    rom[17751] = 25'b1111111010110001101101100;
    rom[17752] = 25'b1111111010110001101001101;
    rom[17753] = 25'b1111111010110001100101110;
    rom[17754] = 25'b1111111010110001100010000;
    rom[17755] = 25'b1111111010110001011110010;
    rom[17756] = 25'b1111111010110001011010100;
    rom[17757] = 25'b1111111010110001010110111;
    rom[17758] = 25'b1111111010110001010011001;
    rom[17759] = 25'b1111111010110001001111100;
    rom[17760] = 25'b1111111010110001001011111;
    rom[17761] = 25'b1111111010110001001000010;
    rom[17762] = 25'b1111111010110001000100110;
    rom[17763] = 25'b1111111010110001000001001;
    rom[17764] = 25'b1111111010110000111101101;
    rom[17765] = 25'b1111111010110000111010001;
    rom[17766] = 25'b1111111010110000110110110;
    rom[17767] = 25'b1111111010110000110011011;
    rom[17768] = 25'b1111111010110000101111111;
    rom[17769] = 25'b1111111010110000101100100;
    rom[17770] = 25'b1111111010110000101001001;
    rom[17771] = 25'b1111111010110000100101111;
    rom[17772] = 25'b1111111010110000100010101;
    rom[17773] = 25'b1111111010110000011111011;
    rom[17774] = 25'b1111111010110000011100001;
    rom[17775] = 25'b1111111010110000011000111;
    rom[17776] = 25'b1111111010110000010101110;
    rom[17777] = 25'b1111111010110000010010101;
    rom[17778] = 25'b1111111010110000001111100;
    rom[17779] = 25'b1111111010110000001100011;
    rom[17780] = 25'b1111111010110000001001011;
    rom[17781] = 25'b1111111010110000000110011;
    rom[17782] = 25'b1111111010110000000011011;
    rom[17783] = 25'b1111111010110000000000011;
    rom[17784] = 25'b1111111010101111111101100;
    rom[17785] = 25'b1111111010101111111010100;
    rom[17786] = 25'b1111111010101111110111101;
    rom[17787] = 25'b1111111010101111110100110;
    rom[17788] = 25'b1111111010101111110010000;
    rom[17789] = 25'b1111111010101111101111001;
    rom[17790] = 25'b1111111010101111101100011;
    rom[17791] = 25'b1111111010101111101001101;
    rom[17792] = 25'b1111111010101111100110111;
    rom[17793] = 25'b1111111010101111100100010;
    rom[17794] = 25'b1111111010101111100001100;
    rom[17795] = 25'b1111111010101111011110111;
    rom[17796] = 25'b1111111010101111011100011;
    rom[17797] = 25'b1111111010101111011001110;
    rom[17798] = 25'b1111111010101111010111001;
    rom[17799] = 25'b1111111010101111010100101;
    rom[17800] = 25'b1111111010101111010010010;
    rom[17801] = 25'b1111111010101111001111110;
    rom[17802] = 25'b1111111010101111001101010;
    rom[17803] = 25'b1111111010101111001011000;
    rom[17804] = 25'b1111111010101111001000100;
    rom[17805] = 25'b1111111010101111000110001;
    rom[17806] = 25'b1111111010101111000011111;
    rom[17807] = 25'b1111111010101111000001101;
    rom[17808] = 25'b1111111010101110111111011;
    rom[17809] = 25'b1111111010101110111101001;
    rom[17810] = 25'b1111111010101110111010111;
    rom[17811] = 25'b1111111010101110111000110;
    rom[17812] = 25'b1111111010101110110110101;
    rom[17813] = 25'b1111111010101110110100100;
    rom[17814] = 25'b1111111010101110110010011;
    rom[17815] = 25'b1111111010101110110000011;
    rom[17816] = 25'b1111111010101110101110010;
    rom[17817] = 25'b1111111010101110101100011;
    rom[17818] = 25'b1111111010101110101010011;
    rom[17819] = 25'b1111111010101110101000011;
    rom[17820] = 25'b1111111010101110100110100;
    rom[17821] = 25'b1111111010101110100100101;
    rom[17822] = 25'b1111111010101110100010110;
    rom[17823] = 25'b1111111010101110100000111;
    rom[17824] = 25'b1111111010101110011111001;
    rom[17825] = 25'b1111111010101110011101011;
    rom[17826] = 25'b1111111010101110011011101;
    rom[17827] = 25'b1111111010101110011001111;
    rom[17828] = 25'b1111111010101110011000010;
    rom[17829] = 25'b1111111010101110010110100;
    rom[17830] = 25'b1111111010101110010101000;
    rom[17831] = 25'b1111111010101110010011011;
    rom[17832] = 25'b1111111010101110010001110;
    rom[17833] = 25'b1111111010101110010000010;
    rom[17834] = 25'b1111111010101110001110110;
    rom[17835] = 25'b1111111010101110001101010;
    rom[17836] = 25'b1111111010101110001011111;
    rom[17837] = 25'b1111111010101110001010011;
    rom[17838] = 25'b1111111010101110001001001;
    rom[17839] = 25'b1111111010101110000111110;
    rom[17840] = 25'b1111111010101110000110011;
    rom[17841] = 25'b1111111010101110000101001;
    rom[17842] = 25'b1111111010101110000011110;
    rom[17843] = 25'b1111111010101110000010101;
    rom[17844] = 25'b1111111010101110000001011;
    rom[17845] = 25'b1111111010101110000000001;
    rom[17846] = 25'b1111111010101101111111000;
    rom[17847] = 25'b1111111010101101111101111;
    rom[17848] = 25'b1111111010101101111100110;
    rom[17849] = 25'b1111111010101101111011110;
    rom[17850] = 25'b1111111010101101111010110;
    rom[17851] = 25'b1111111010101101111001110;
    rom[17852] = 25'b1111111010101101111000110;
    rom[17853] = 25'b1111111010101101110111111;
    rom[17854] = 25'b1111111010101101110110111;
    rom[17855] = 25'b1111111010101101110110000;
    rom[17856] = 25'b1111111010101101110101001;
    rom[17857] = 25'b1111111010101101110100010;
    rom[17858] = 25'b1111111010101101110011100;
    rom[17859] = 25'b1111111010101101110010110;
    rom[17860] = 25'b1111111010101101110010000;
    rom[17861] = 25'b1111111010101101110001010;
    rom[17862] = 25'b1111111010101101110000101;
    rom[17863] = 25'b1111111010101101110000000;
    rom[17864] = 25'b1111111010101101101111011;
    rom[17865] = 25'b1111111010101101101110110;
    rom[17866] = 25'b1111111010101101101110010;
    rom[17867] = 25'b1111111010101101101101101;
    rom[17868] = 25'b1111111010101101101101001;
    rom[17869] = 25'b1111111010101101101100110;
    rom[17870] = 25'b1111111010101101101100010;
    rom[17871] = 25'b1111111010101101101011111;
    rom[17872] = 25'b1111111010101101101011100;
    rom[17873] = 25'b1111111010101101101011001;
    rom[17874] = 25'b1111111010101101101010110;
    rom[17875] = 25'b1111111010101101101010100;
    rom[17876] = 25'b1111111010101101101010010;
    rom[17877] = 25'b1111111010101101101010000;
    rom[17878] = 25'b1111111010101101101001111;
    rom[17879] = 25'b1111111010101101101001101;
    rom[17880] = 25'b1111111010101101101001100;
    rom[17881] = 25'b1111111010101101101001011;
    rom[17882] = 25'b1111111010101101101001010;
    rom[17883] = 25'b1111111010101101101001010;
    rom[17884] = 25'b1111111010101101101001010;
    rom[17885] = 25'b1111111010101101101001010;
    rom[17886] = 25'b1111111010101101101001010;
    rom[17887] = 25'b1111111010101101101001011;
    rom[17888] = 25'b1111111010101101101001100;
    rom[17889] = 25'b1111111010101101101001100;
    rom[17890] = 25'b1111111010101101101001110;
    rom[17891] = 25'b1111111010101101101001111;
    rom[17892] = 25'b1111111010101101101010010;
    rom[17893] = 25'b1111111010101101101010011;
    rom[17894] = 25'b1111111010101101101010101;
    rom[17895] = 25'b1111111010101101101011000;
    rom[17896] = 25'b1111111010101101101011011;
    rom[17897] = 25'b1111111010101101101011110;
    rom[17898] = 25'b1111111010101101101100001;
    rom[17899] = 25'b1111111010101101101100100;
    rom[17900] = 25'b1111111010101101101101000;
    rom[17901] = 25'b1111111010101101101101100;
    rom[17902] = 25'b1111111010101101101110000;
    rom[17903] = 25'b1111111010101101101110101;
    rom[17904] = 25'b1111111010101101101111001;
    rom[17905] = 25'b1111111010101101101111110;
    rom[17906] = 25'b1111111010101101110000011;
    rom[17907] = 25'b1111111010101101110001001;
    rom[17908] = 25'b1111111010101101110001110;
    rom[17909] = 25'b1111111010101101110010100;
    rom[17910] = 25'b1111111010101101110011010;
    rom[17911] = 25'b1111111010101101110100001;
    rom[17912] = 25'b1111111010101101110100111;
    rom[17913] = 25'b1111111010101101110101110;
    rom[17914] = 25'b1111111010101101110110101;
    rom[17915] = 25'b1111111010101101110111100;
    rom[17916] = 25'b1111111010101101111000100;
    rom[17917] = 25'b1111111010101101111001100;
    rom[17918] = 25'b1111111010101101111010100;
    rom[17919] = 25'b1111111010101101111011101;
    rom[17920] = 25'b1111111010101101111100101;
    rom[17921] = 25'b1111111010101101111101110;
    rom[17922] = 25'b1111111010101101111110111;
    rom[17923] = 25'b1111111010101110000000000;
    rom[17924] = 25'b1111111010101110000001001;
    rom[17925] = 25'b1111111010101110000010011;
    rom[17926] = 25'b1111111010101110000011110;
    rom[17927] = 25'b1111111010101110000101000;
    rom[17928] = 25'b1111111010101110000110010;
    rom[17929] = 25'b1111111010101110000111101;
    rom[17930] = 25'b1111111010101110001001000;
    rom[17931] = 25'b1111111010101110001010011;
    rom[17932] = 25'b1111111010101110001011111;
    rom[17933] = 25'b1111111010101110001101010;
    rom[17934] = 25'b1111111010101110001110110;
    rom[17935] = 25'b1111111010101110010000011;
    rom[17936] = 25'b1111111010101110010001111;
    rom[17937] = 25'b1111111010101110010011100;
    rom[17938] = 25'b1111111010101110010101001;
    rom[17939] = 25'b1111111010101110010110110;
    rom[17940] = 25'b1111111010101110011000011;
    rom[17941] = 25'b1111111010101110011010010;
    rom[17942] = 25'b1111111010101110011100000;
    rom[17943] = 25'b1111111010101110011101110;
    rom[17944] = 25'b1111111010101110011111100;
    rom[17945] = 25'b1111111010101110100001011;
    rom[17946] = 25'b1111111010101110100011010;
    rom[17947] = 25'b1111111010101110100101001;
    rom[17948] = 25'b1111111010101110100111001;
    rom[17949] = 25'b1111111010101110101001000;
    rom[17950] = 25'b1111111010101110101011000;
    rom[17951] = 25'b1111111010101110101101000;
    rom[17952] = 25'b1111111010101110101111001;
    rom[17953] = 25'b1111111010101110110001001;
    rom[17954] = 25'b1111111010101110110011011;
    rom[17955] = 25'b1111111010101110110101100;
    rom[17956] = 25'b1111111010101110110111101;
    rom[17957] = 25'b1111111010101110111001111;
    rom[17958] = 25'b1111111010101110111100001;
    rom[17959] = 25'b1111111010101110111110011;
    rom[17960] = 25'b1111111010101111000000101;
    rom[17961] = 25'b1111111010101111000011000;
    rom[17962] = 25'b1111111010101111000101011;
    rom[17963] = 25'b1111111010101111000111110;
    rom[17964] = 25'b1111111010101111001010010;
    rom[17965] = 25'b1111111010101111001100101;
    rom[17966] = 25'b1111111010101111001111001;
    rom[17967] = 25'b1111111010101111010001101;
    rom[17968] = 25'b1111111010101111010100010;
    rom[17969] = 25'b1111111010101111010110110;
    rom[17970] = 25'b1111111010101111011001011;
    rom[17971] = 25'b1111111010101111011100000;
    rom[17972] = 25'b1111111010101111011110110;
    rom[17973] = 25'b1111111010101111100001100;
    rom[17974] = 25'b1111111010101111100100010;
    rom[17975] = 25'b1111111010101111100111000;
    rom[17976] = 25'b1111111010101111101001110;
    rom[17977] = 25'b1111111010101111101100101;
    rom[17978] = 25'b1111111010101111101111100;
    rom[17979] = 25'b1111111010101111110010011;
    rom[17980] = 25'b1111111010101111110101011;
    rom[17981] = 25'b1111111010101111111000010;
    rom[17982] = 25'b1111111010101111111011010;
    rom[17983] = 25'b1111111010101111111110010;
    rom[17984] = 25'b1111111010110000000001011;
    rom[17985] = 25'b1111111010110000000100100;
    rom[17986] = 25'b1111111010110000000111100;
    rom[17987] = 25'b1111111010110000001010110;
    rom[17988] = 25'b1111111010110000001101111;
    rom[17989] = 25'b1111111010110000010001001;
    rom[17990] = 25'b1111111010110000010100011;
    rom[17991] = 25'b1111111010110000010111101;
    rom[17992] = 25'b1111111010110000011010111;
    rom[17993] = 25'b1111111010110000011110010;
    rom[17994] = 25'b1111111010110000100001101;
    rom[17995] = 25'b1111111010110000100101001;
    rom[17996] = 25'b1111111010110000101000011;
    rom[17997] = 25'b1111111010110000101100000;
    rom[17998] = 25'b1111111010110000101111011;
    rom[17999] = 25'b1111111010110000110011000;
    rom[18000] = 25'b1111111010110000110110100;
    rom[18001] = 25'b1111111010110000111010001;
    rom[18002] = 25'b1111111010110000111101110;
    rom[18003] = 25'b1111111010110001000001011;
    rom[18004] = 25'b1111111010110001000101001;
    rom[18005] = 25'b1111111010110001001000111;
    rom[18006] = 25'b1111111010110001001100101;
    rom[18007] = 25'b1111111010110001010000010;
    rom[18008] = 25'b1111111010110001010100001;
    rom[18009] = 25'b1111111010110001011000000;
    rom[18010] = 25'b1111111010110001011011111;
    rom[18011] = 25'b1111111010110001011111110;
    rom[18012] = 25'b1111111010110001100011110;
    rom[18013] = 25'b1111111010110001100111101;
    rom[18014] = 25'b1111111010110001101011101;
    rom[18015] = 25'b1111111010110001101111101;
    rom[18016] = 25'b1111111010110001110011110;
    rom[18017] = 25'b1111111010110001110111111;
    rom[18018] = 25'b1111111010110001111100000;
    rom[18019] = 25'b1111111010110010000000010;
    rom[18020] = 25'b1111111010110010000100011;
    rom[18021] = 25'b1111111010110010001000101;
    rom[18022] = 25'b1111111010110010001100111;
    rom[18023] = 25'b1111111010110010010001001;
    rom[18024] = 25'b1111111010110010010101011;
    rom[18025] = 25'b1111111010110010011001110;
    rom[18026] = 25'b1111111010110010011110001;
    rom[18027] = 25'b1111111010110010100010101;
    rom[18028] = 25'b1111111010110010100111000;
    rom[18029] = 25'b1111111010110010101011100;
    rom[18030] = 25'b1111111010110010110000000;
    rom[18031] = 25'b1111111010110010110100101;
    rom[18032] = 25'b1111111010110010111001001;
    rom[18033] = 25'b1111111010110010111101110;
    rom[18034] = 25'b1111111010110011000010011;
    rom[18035] = 25'b1111111010110011000111001;
    rom[18036] = 25'b1111111010110011001011110;
    rom[18037] = 25'b1111111010110011010000100;
    rom[18038] = 25'b1111111010110011010101010;
    rom[18039] = 25'b1111111010110011011010000;
    rom[18040] = 25'b1111111010110011011110111;
    rom[18041] = 25'b1111111010110011100011110;
    rom[18042] = 25'b1111111010110011101000110;
    rom[18043] = 25'b1111111010110011101101101;
    rom[18044] = 25'b1111111010110011110010101;
    rom[18045] = 25'b1111111010110011110111100;
    rom[18046] = 25'b1111111010110011111100101;
    rom[18047] = 25'b1111111010110100000001101;
    rom[18048] = 25'b1111111010110100000110101;
    rom[18049] = 25'b1111111010110100001011111;
    rom[18050] = 25'b1111111010110100010001000;
    rom[18051] = 25'b1111111010110100010110010;
    rom[18052] = 25'b1111111010110100011011011;
    rom[18053] = 25'b1111111010110100100000101;
    rom[18054] = 25'b1111111010110100100110000;
    rom[18055] = 25'b1111111010110100101011010;
    rom[18056] = 25'b1111111010110100110000101;
    rom[18057] = 25'b1111111010110100110110000;
    rom[18058] = 25'b1111111010110100111011011;
    rom[18059] = 25'b1111111010110101000000111;
    rom[18060] = 25'b1111111010110101000110010;
    rom[18061] = 25'b1111111010110101001011110;
    rom[18062] = 25'b1111111010110101010001010;
    rom[18063] = 25'b1111111010110101010110111;
    rom[18064] = 25'b1111111010110101011100100;
    rom[18065] = 25'b1111111010110101100010001;
    rom[18066] = 25'b1111111010110101100111110;
    rom[18067] = 25'b1111111010110101101101100;
    rom[18068] = 25'b1111111010110101110011010;
    rom[18069] = 25'b1111111010110101111001000;
    rom[18070] = 25'b1111111010110101111110110;
    rom[18071] = 25'b1111111010110110000100101;
    rom[18072] = 25'b1111111010110110001010100;
    rom[18073] = 25'b1111111010110110010000011;
    rom[18074] = 25'b1111111010110110010110011;
    rom[18075] = 25'b1111111010110110011100010;
    rom[18076] = 25'b1111111010110110100010010;
    rom[18077] = 25'b1111111010110110101000010;
    rom[18078] = 25'b1111111010110110101110011;
    rom[18079] = 25'b1111111010110110110100011;
    rom[18080] = 25'b1111111010110110111010100;
    rom[18081] = 25'b1111111010110111000000110;
    rom[18082] = 25'b1111111010110111000110111;
    rom[18083] = 25'b1111111010110111001101001;
    rom[18084] = 25'b1111111010110111010011011;
    rom[18085] = 25'b1111111010110111011001101;
    rom[18086] = 25'b1111111010110111011111111;
    rom[18087] = 25'b1111111010110111100110010;
    rom[18088] = 25'b1111111010110111101100110;
    rom[18089] = 25'b1111111010110111110011000;
    rom[18090] = 25'b1111111010110111111001100;
    rom[18091] = 25'b1111111010111000000000000;
    rom[18092] = 25'b1111111010111000000110100;
    rom[18093] = 25'b1111111010111000001101000;
    rom[18094] = 25'b1111111010111000010011101;
    rom[18095] = 25'b1111111010111000011010010;
    rom[18096] = 25'b1111111010111000100000111;
    rom[18097] = 25'b1111111010111000100111100;
    rom[18098] = 25'b1111111010111000101110010;
    rom[18099] = 25'b1111111010111000110101000;
    rom[18100] = 25'b1111111010111000111011110;
    rom[18101] = 25'b1111111010111001000010100;
    rom[18102] = 25'b1111111010111001001001011;
    rom[18103] = 25'b1111111010111001010000010;
    rom[18104] = 25'b1111111010111001010111001;
    rom[18105] = 25'b1111111010111001011110001;
    rom[18106] = 25'b1111111010111001100101001;
    rom[18107] = 25'b1111111010111001101100001;
    rom[18108] = 25'b1111111010111001110011001;
    rom[18109] = 25'b1111111010111001111010001;
    rom[18110] = 25'b1111111010111010000001001;
    rom[18111] = 25'b1111111010111010001000011;
    rom[18112] = 25'b1111111010111010001111100;
    rom[18113] = 25'b1111111010111010010110101;
    rom[18114] = 25'b1111111010111010011110000;
    rom[18115] = 25'b1111111010111010100101001;
    rom[18116] = 25'b1111111010111010101100100;
    rom[18117] = 25'b1111111010111010110011110;
    rom[18118] = 25'b1111111010111010111011001;
    rom[18119] = 25'b1111111010111011000010100;
    rom[18120] = 25'b1111111010111011001001111;
    rom[18121] = 25'b1111111010111011010001011;
    rom[18122] = 25'b1111111010111011011000111;
    rom[18123] = 25'b1111111010111011100000100;
    rom[18124] = 25'b1111111010111011101000000;
    rom[18125] = 25'b1111111010111011101111101;
    rom[18126] = 25'b1111111010111011110111001;
    rom[18127] = 25'b1111111010111011111110110;
    rom[18128] = 25'b1111111010111100000110100;
    rom[18129] = 25'b1111111010111100001110010;
    rom[18130] = 25'b1111111010111100010110000;
    rom[18131] = 25'b1111111010111100011101110;
    rom[18132] = 25'b1111111010111100100101100;
    rom[18133] = 25'b1111111010111100101101011;
    rom[18134] = 25'b1111111010111100110101010;
    rom[18135] = 25'b1111111010111100111101001;
    rom[18136] = 25'b1111111010111101000101001;
    rom[18137] = 25'b1111111010111101001101000;
    rom[18138] = 25'b1111111010111101010101001;
    rom[18139] = 25'b1111111010111101011101001;
    rom[18140] = 25'b1111111010111101100101010;
    rom[18141] = 25'b1111111010111101101101011;
    rom[18142] = 25'b1111111010111101110101100;
    rom[18143] = 25'b1111111010111101111101101;
    rom[18144] = 25'b1111111010111110000101111;
    rom[18145] = 25'b1111111010111110001110000;
    rom[18146] = 25'b1111111010111110010110011;
    rom[18147] = 25'b1111111010111110011110101;
    rom[18148] = 25'b1111111010111110100111000;
    rom[18149] = 25'b1111111010111110101111011;
    rom[18150] = 25'b1111111010111110110111110;
    rom[18151] = 25'b1111111010111111000000010;
    rom[18152] = 25'b1111111010111111001000110;
    rom[18153] = 25'b1111111010111111010001010;
    rom[18154] = 25'b1111111010111111011001110;
    rom[18155] = 25'b1111111010111111100010010;
    rom[18156] = 25'b1111111010111111101010111;
    rom[18157] = 25'b1111111010111111110011100;
    rom[18158] = 25'b1111111010111111111100001;
    rom[18159] = 25'b1111111011000000000100111;
    rom[18160] = 25'b1111111011000000001101101;
    rom[18161] = 25'b1111111011000000010110011;
    rom[18162] = 25'b1111111011000000011111001;
    rom[18163] = 25'b1111111011000000101000000;
    rom[18164] = 25'b1111111011000000110000111;
    rom[18165] = 25'b1111111011000000111001110;
    rom[18166] = 25'b1111111011000001000010101;
    rom[18167] = 25'b1111111011000001001011101;
    rom[18168] = 25'b1111111011000001010100101;
    rom[18169] = 25'b1111111011000001011101101;
    rom[18170] = 25'b1111111011000001100110110;
    rom[18171] = 25'b1111111011000001101111110;
    rom[18172] = 25'b1111111011000001111000111;
    rom[18173] = 25'b1111111011000010000010001;
    rom[18174] = 25'b1111111011000010001011010;
    rom[18175] = 25'b1111111011000010010100100;
    rom[18176] = 25'b1111111011000010011101110;
    rom[18177] = 25'b1111111011000010100111000;
    rom[18178] = 25'b1111111011000010110000011;
    rom[18179] = 25'b1111111011000010111001110;
    rom[18180] = 25'b1111111011000011000011001;
    rom[18181] = 25'b1111111011000011001100100;
    rom[18182] = 25'b1111111011000011010101111;
    rom[18183] = 25'b1111111011000011011111100;
    rom[18184] = 25'b1111111011000011101001000;
    rom[18185] = 25'b1111111011000011110010100;
    rom[18186] = 25'b1111111011000011111100001;
    rom[18187] = 25'b1111111011000100000101110;
    rom[18188] = 25'b1111111011000100001111011;
    rom[18189] = 25'b1111111011000100011001001;
    rom[18190] = 25'b1111111011000100100010110;
    rom[18191] = 25'b1111111011000100101100100;
    rom[18192] = 25'b1111111011000100110110010;
    rom[18193] = 25'b1111111011000101000000001;
    rom[18194] = 25'b1111111011000101001010000;
    rom[18195] = 25'b1111111011000101010011111;
    rom[18196] = 25'b1111111011000101011101110;
    rom[18197] = 25'b1111111011000101100111110;
    rom[18198] = 25'b1111111011000101110001110;
    rom[18199] = 25'b1111111011000101111011110;
    rom[18200] = 25'b1111111011000110000101110;
    rom[18201] = 25'b1111111011000110001111111;
    rom[18202] = 25'b1111111011000110011010000;
    rom[18203] = 25'b1111111011000110100100001;
    rom[18204] = 25'b1111111011000110101110010;
    rom[18205] = 25'b1111111011000110111000100;
    rom[18206] = 25'b1111111011000111000010110;
    rom[18207] = 25'b1111111011000111001101000;
    rom[18208] = 25'b1111111011000111010111010;
    rom[18209] = 25'b1111111011000111100001101;
    rom[18210] = 25'b1111111011000111101100000;
    rom[18211] = 25'b1111111011000111110110100;
    rom[18212] = 25'b1111111011001000000001000;
    rom[18213] = 25'b1111111011001000001011011;
    rom[18214] = 25'b1111111011001000010101111;
    rom[18215] = 25'b1111111011001000100000011;
    rom[18216] = 25'b1111111011001000101011001;
    rom[18217] = 25'b1111111011001000110101101;
    rom[18218] = 25'b1111111011001001000000010;
    rom[18219] = 25'b1111111011001001001010111;
    rom[18220] = 25'b1111111011001001010101101;
    rom[18221] = 25'b1111111011001001100000011;
    rom[18222] = 25'b1111111011001001101011001;
    rom[18223] = 25'b1111111011001001110110000;
    rom[18224] = 25'b1111111011001010000000110;
    rom[18225] = 25'b1111111011001010001011110;
    rom[18226] = 25'b1111111011001010010110100;
    rom[18227] = 25'b1111111011001010100001101;
    rom[18228] = 25'b1111111011001010101100100;
    rom[18229] = 25'b1111111011001010110111100;
    rom[18230] = 25'b1111111011001011000010100;
    rom[18231] = 25'b1111111011001011001101101;
    rom[18232] = 25'b1111111011001011011000110;
    rom[18233] = 25'b1111111011001011100011111;
    rom[18234] = 25'b1111111011001011101111001;
    rom[18235] = 25'b1111111011001011111010010;
    rom[18236] = 25'b1111111011001100000101100;
    rom[18237] = 25'b1111111011001100010000110;
    rom[18238] = 25'b1111111011001100011100001;
    rom[18239] = 25'b1111111011001100100111011;
    rom[18240] = 25'b1111111011001100110010110;
    rom[18241] = 25'b1111111011001100111110010;
    rom[18242] = 25'b1111111011001101001001101;
    rom[18243] = 25'b1111111011001101010101001;
    rom[18244] = 25'b1111111011001101100000100;
    rom[18245] = 25'b1111111011001101101100001;
    rom[18246] = 25'b1111111011001101110111110;
    rom[18247] = 25'b1111111011001110000011010;
    rom[18248] = 25'b1111111011001110001110111;
    rom[18249] = 25'b1111111011001110011010100;
    rom[18250] = 25'b1111111011001110100110011;
    rom[18251] = 25'b1111111011001110110010000;
    rom[18252] = 25'b1111111011001110111101110;
    rom[18253] = 25'b1111111011001111001001101;
    rom[18254] = 25'b1111111011001111010101011;
    rom[18255] = 25'b1111111011001111100001010;
    rom[18256] = 25'b1111111011001111101101010;
    rom[18257] = 25'b1111111011001111111001000;
    rom[18258] = 25'b1111111011010000000101001;
    rom[18259] = 25'b1111111011010000010001000;
    rom[18260] = 25'b1111111011010000011101001;
    rom[18261] = 25'b1111111011010000101001001;
    rom[18262] = 25'b1111111011010000110101010;
    rom[18263] = 25'b1111111011010001000001011;
    rom[18264] = 25'b1111111011010001001101101;
    rom[18265] = 25'b1111111011010001011001110;
    rom[18266] = 25'b1111111011010001100110000;
    rom[18267] = 25'b1111111011010001110010010;
    rom[18268] = 25'b1111111011010001111110100;
    rom[18269] = 25'b1111111011010010001010111;
    rom[18270] = 25'b1111111011010010010111010;
    rom[18271] = 25'b1111111011010010100011101;
    rom[18272] = 25'b1111111011010010110000000;
    rom[18273] = 25'b1111111011010010111100100;
    rom[18274] = 25'b1111111011010011001001000;
    rom[18275] = 25'b1111111011010011010101100;
    rom[18276] = 25'b1111111011010011100010000;
    rom[18277] = 25'b1111111011010011101110101;
    rom[18278] = 25'b1111111011010011111011010;
    rom[18279] = 25'b1111111011010100001000000;
    rom[18280] = 25'b1111111011010100010100101;
    rom[18281] = 25'b1111111011010100100001011;
    rom[18282] = 25'b1111111011010100101110001;
    rom[18283] = 25'b1111111011010100111011000;
    rom[18284] = 25'b1111111011010101000111110;
    rom[18285] = 25'b1111111011010101010100101;
    rom[18286] = 25'b1111111011010101100001100;
    rom[18287] = 25'b1111111011010101101110011;
    rom[18288] = 25'b1111111011010101111011011;
    rom[18289] = 25'b1111111011010110001000011;
    rom[18290] = 25'b1111111011010110010101011;
    rom[18291] = 25'b1111111011010110100010011;
    rom[18292] = 25'b1111111011010110101111100;
    rom[18293] = 25'b1111111011010110111100101;
    rom[18294] = 25'b1111111011010111001001111;
    rom[18295] = 25'b1111111011010111010111000;
    rom[18296] = 25'b1111111011010111100100010;
    rom[18297] = 25'b1111111011010111110001100;
    rom[18298] = 25'b1111111011010111111110110;
    rom[18299] = 25'b1111111011011000001100000;
    rom[18300] = 25'b1111111011011000011001011;
    rom[18301] = 25'b1111111011011000100110111;
    rom[18302] = 25'b1111111011011000110100010;
    rom[18303] = 25'b1111111011011001000001101;
    rom[18304] = 25'b1111111011011001001111010;
    rom[18305] = 25'b1111111011011001011100110;
    rom[18306] = 25'b1111111011011001101010010;
    rom[18307] = 25'b1111111011011001110111111;
    rom[18308] = 25'b1111111011011010000101100;
    rom[18309] = 25'b1111111011011010010011001;
    rom[18310] = 25'b1111111011011010100000111;
    rom[18311] = 25'b1111111011011010101110100;
    rom[18312] = 25'b1111111011011010111100010;
    rom[18313] = 25'b1111111011011011001010000;
    rom[18314] = 25'b1111111011011011010111111;
    rom[18315] = 25'b1111111011011011100101110;
    rom[18316] = 25'b1111111011011011110011100;
    rom[18317] = 25'b1111111011011100000001100;
    rom[18318] = 25'b1111111011011100001111100;
    rom[18319] = 25'b1111111011011100011101011;
    rom[18320] = 25'b1111111011011100101011011;
    rom[18321] = 25'b1111111011011100111001100;
    rom[18322] = 25'b1111111011011101000111101;
    rom[18323] = 25'b1111111011011101010101110;
    rom[18324] = 25'b1111111011011101100011110;
    rom[18325] = 25'b1111111011011101110010000;
    rom[18326] = 25'b1111111011011110000000010;
    rom[18327] = 25'b1111111011011110001110100;
    rom[18328] = 25'b1111111011011110011100110;
    rom[18329] = 25'b1111111011011110101011001;
    rom[18330] = 25'b1111111011011110111001011;
    rom[18331] = 25'b1111111011011111000111110;
    rom[18332] = 25'b1111111011011111010110010;
    rom[18333] = 25'b1111111011011111100100101;
    rom[18334] = 25'b1111111011011111110011001;
    rom[18335] = 25'b1111111011100000000001101;
    rom[18336] = 25'b1111111011100000010000001;
    rom[18337] = 25'b1111111011100000011110101;
    rom[18338] = 25'b1111111011100000101101011;
    rom[18339] = 25'b1111111011100000111100000;
    rom[18340] = 25'b1111111011100001001010101;
    rom[18341] = 25'b1111111011100001011001011;
    rom[18342] = 25'b1111111011100001101000001;
    rom[18343] = 25'b1111111011100001110110111;
    rom[18344] = 25'b1111111011100010000101101;
    rom[18345] = 25'b1111111011100010010100100;
    rom[18346] = 25'b1111111011100010100011011;
    rom[18347] = 25'b1111111011100010110010010;
    rom[18348] = 25'b1111111011100011000001001;
    rom[18349] = 25'b1111111011100011010000010;
    rom[18350] = 25'b1111111011100011011111001;
    rom[18351] = 25'b1111111011100011101110001;
    rom[18352] = 25'b1111111011100011111101011;
    rom[18353] = 25'b1111111011100100001100011;
    rom[18354] = 25'b1111111011100100011011100;
    rom[18355] = 25'b1111111011100100101010110;
    rom[18356] = 25'b1111111011100100111001111;
    rom[18357] = 25'b1111111011100101001001001;
    rom[18358] = 25'b1111111011100101011000011;
    rom[18359] = 25'b1111111011100101100111101;
    rom[18360] = 25'b1111111011100101110111000;
    rom[18361] = 25'b1111111011100110000110011;
    rom[18362] = 25'b1111111011100110010101110;
    rom[18363] = 25'b1111111011100110100101010;
    rom[18364] = 25'b1111111011100110110100101;
    rom[18365] = 25'b1111111011100111000100001;
    rom[18366] = 25'b1111111011100111010011101;
    rom[18367] = 25'b1111111011100111100011010;
    rom[18368] = 25'b1111111011100111110010111;
    rom[18369] = 25'b1111111011101000000010011;
    rom[18370] = 25'b1111111011101000010010001;
    rom[18371] = 25'b1111111011101000100001110;
    rom[18372] = 25'b1111111011101000110001100;
    rom[18373] = 25'b1111111011101001000001010;
    rom[18374] = 25'b1111111011101001010001000;
    rom[18375] = 25'b1111111011101001100000111;
    rom[18376] = 25'b1111111011101001110000110;
    rom[18377] = 25'b1111111011101010000000101;
    rom[18378] = 25'b1111111011101010010000100;
    rom[18379] = 25'b1111111011101010100000100;
    rom[18380] = 25'b1111111011101010110000100;
    rom[18381] = 25'b1111111011101011000000100;
    rom[18382] = 25'b1111111011101011010000100;
    rom[18383] = 25'b1111111011101011100000101;
    rom[18384] = 25'b1111111011101011110000110;
    rom[18385] = 25'b1111111011101100000000111;
    rom[18386] = 25'b1111111011101100010001000;
    rom[18387] = 25'b1111111011101100100001010;
    rom[18388] = 25'b1111111011101100110001100;
    rom[18389] = 25'b1111111011101101000001110;
    rom[18390] = 25'b1111111011101101010010001;
    rom[18391] = 25'b1111111011101101100010100;
    rom[18392] = 25'b1111111011101101110010111;
    rom[18393] = 25'b1111111011101110000011010;
    rom[18394] = 25'b1111111011101110010011110;
    rom[18395] = 25'b1111111011101110100100010;
    rom[18396] = 25'b1111111011101110110100101;
    rom[18397] = 25'b1111111011101111000101010;
    rom[18398] = 25'b1111111011101111010101111;
    rom[18399] = 25'b1111111011101111100110100;
    rom[18400] = 25'b1111111011101111110111001;
    rom[18401] = 25'b1111111011110000000111110;
    rom[18402] = 25'b1111111011110000011000011;
    rom[18403] = 25'b1111111011110000101001001;
    rom[18404] = 25'b1111111011110000111001111;
    rom[18405] = 25'b1111111011110001001010110;
    rom[18406] = 25'b1111111011110001011011100;
    rom[18407] = 25'b1111111011110001101100100;
    rom[18408] = 25'b1111111011110001111101011;
    rom[18409] = 25'b1111111011110010001110010;
    rom[18410] = 25'b1111111011110010011111010;
    rom[18411] = 25'b1111111011110010110000010;
    rom[18412] = 25'b1111111011110011000001010;
    rom[18413] = 25'b1111111011110011010010011;
    rom[18414] = 25'b1111111011110011100011011;
    rom[18415] = 25'b1111111011110011110100100;
    rom[18416] = 25'b1111111011110100000101110;
    rom[18417] = 25'b1111111011110100010110111;
    rom[18418] = 25'b1111111011110100101000001;
    rom[18419] = 25'b1111111011110100111001011;
    rom[18420] = 25'b1111111011110101001010101;
    rom[18421] = 25'b1111111011110101011100000;
    rom[18422] = 25'b1111111011110101101101011;
    rom[18423] = 25'b1111111011110101111110110;
    rom[18424] = 25'b1111111011110110010000001;
    rom[18425] = 25'b1111111011110110100001101;
    rom[18426] = 25'b1111111011110110110011001;
    rom[18427] = 25'b1111111011110111000100101;
    rom[18428] = 25'b1111111011110111010110001;
    rom[18429] = 25'b1111111011110111100111110;
    rom[18430] = 25'b1111111011110111111001011;
    rom[18431] = 25'b1111111011111000001011000;
    rom[18432] = 25'b1111111011111000011100101;
    rom[18433] = 25'b1111111011111000101110011;
    rom[18434] = 25'b1111111011111001000000001;
    rom[18435] = 25'b1111111011111001010001111;
    rom[18436] = 25'b1111111011111001100011110;
    rom[18437] = 25'b1111111011111001110101100;
    rom[18438] = 25'b1111111011111010000111011;
    rom[18439] = 25'b1111111011111010011001011;
    rom[18440] = 25'b1111111011111010101011010;
    rom[18441] = 25'b1111111011111010111101001;
    rom[18442] = 25'b1111111011111011001111010;
    rom[18443] = 25'b1111111011111011100001010;
    rom[18444] = 25'b1111111011111011110011011;
    rom[18445] = 25'b1111111011111100000101100;
    rom[18446] = 25'b1111111011111100010111101;
    rom[18447] = 25'b1111111011111100101001110;
    rom[18448] = 25'b1111111011111100111011111;
    rom[18449] = 25'b1111111011111101001110001;
    rom[18450] = 25'b1111111011111101100000011;
    rom[18451] = 25'b1111111011111101110010110;
    rom[18452] = 25'b1111111011111110000101000;
    rom[18453] = 25'b1111111011111110010111011;
    rom[18454] = 25'b1111111011111110101001110;
    rom[18455] = 25'b1111111011111110111100001;
    rom[18456] = 25'b1111111011111111001110101;
    rom[18457] = 25'b1111111011111111100001001;
    rom[18458] = 25'b1111111011111111110011101;
    rom[18459] = 25'b1111111100000000000110010;
    rom[18460] = 25'b1111111100000000011000110;
    rom[18461] = 25'b1111111100000000101011011;
    rom[18462] = 25'b1111111100000000111110000;
    rom[18463] = 25'b1111111100000001010000110;
    rom[18464] = 25'b1111111100000001100011011;
    rom[18465] = 25'b1111111100000001110110001;
    rom[18466] = 25'b1111111100000010001000111;
    rom[18467] = 25'b1111111100000010011011110;
    rom[18468] = 25'b1111111100000010101110101;
    rom[18469] = 25'b1111111100000011000001011;
    rom[18470] = 25'b1111111100000011010100010;
    rom[18471] = 25'b1111111100000011100111010;
    rom[18472] = 25'b1111111100000011111010010;
    rom[18473] = 25'b1111111100000100001101010;
    rom[18474] = 25'b1111111100000100100000010;
    rom[18475] = 25'b1111111100000100110011010;
    rom[18476] = 25'b1111111100000101000110011;
    rom[18477] = 25'b1111111100000101011001100;
    rom[18478] = 25'b1111111100000101101100110;
    rom[18479] = 25'b1111111100000101111111111;
    rom[18480] = 25'b1111111100000110010011001;
    rom[18481] = 25'b1111111100000110100110011;
    rom[18482] = 25'b1111111100000110111001101;
    rom[18483] = 25'b1111111100000111001101000;
    rom[18484] = 25'b1111111100000111100000011;
    rom[18485] = 25'b1111111100000111110011101;
    rom[18486] = 25'b1111111100001000000111001;
    rom[18487] = 25'b1111111100001000011010100;
    rom[18488] = 25'b1111111100001000101110000;
    rom[18489] = 25'b1111111100001001000001100;
    rom[18490] = 25'b1111111100001001010101000;
    rom[18491] = 25'b1111111100001001101000101;
    rom[18492] = 25'b1111111100001001111100001;
    rom[18493] = 25'b1111111100001010001111111;
    rom[18494] = 25'b1111111100001010100011100;
    rom[18495] = 25'b1111111100001010110111010;
    rom[18496] = 25'b1111111100001011001010111;
    rom[18497] = 25'b1111111100001011011110110;
    rom[18498] = 25'b1111111100001011110010100;
    rom[18499] = 25'b1111111100001100000110010;
    rom[18500] = 25'b1111111100001100011010010;
    rom[18501] = 25'b1111111100001100101110001;
    rom[18502] = 25'b1111111100001101000010000;
    rom[18503] = 25'b1111111100001101010110000;
    rom[18504] = 25'b1111111100001101101010000;
    rom[18505] = 25'b1111111100001101111101111;
    rom[18506] = 25'b1111111100001110010010000;
    rom[18507] = 25'b1111111100001110100110001;
    rom[18508] = 25'b1111111100001110111010001;
    rom[18509] = 25'b1111111100001111001110011;
    rom[18510] = 25'b1111111100001111100010100;
    rom[18511] = 25'b1111111100001111110110101;
    rom[18512] = 25'b1111111100010000001011000;
    rom[18513] = 25'b1111111100010000011111010;
    rom[18514] = 25'b1111111100010000110011100;
    rom[18515] = 25'b1111111100010001000111111;
    rom[18516] = 25'b1111111100010001011100001;
    rom[18517] = 25'b1111111100010001110000100;
    rom[18518] = 25'b1111111100010010000101000;
    rom[18519] = 25'b1111111100010010011001100;
    rom[18520] = 25'b1111111100010010101101111;
    rom[18521] = 25'b1111111100010011000010100;
    rom[18522] = 25'b1111111100010011010111000;
    rom[18523] = 25'b1111111100010011101011100;
    rom[18524] = 25'b1111111100010100000000001;
    rom[18525] = 25'b1111111100010100010100111;
    rom[18526] = 25'b1111111100010100101001100;
    rom[18527] = 25'b1111111100010100111110001;
    rom[18528] = 25'b1111111100010101010010111;
    rom[18529] = 25'b1111111100010101100111110;
    rom[18530] = 25'b1111111100010101111100100;
    rom[18531] = 25'b1111111100010110010001011;
    rom[18532] = 25'b1111111100010110100110010;
    rom[18533] = 25'b1111111100010110111011001;
    rom[18534] = 25'b1111111100010111010000000;
    rom[18535] = 25'b1111111100010111100101000;
    rom[18536] = 25'b1111111100010111111010000;
    rom[18537] = 25'b1111111100011000001111000;
    rom[18538] = 25'b1111111100011000100100000;
    rom[18539] = 25'b1111111100011000111001001;
    rom[18540] = 25'b1111111100011001001110010;
    rom[18541] = 25'b1111111100011001100011011;
    rom[18542] = 25'b1111111100011001111000100;
    rom[18543] = 25'b1111111100011010001101110;
    rom[18544] = 25'b1111111100011010100011000;
    rom[18545] = 25'b1111111100011010111000010;
    rom[18546] = 25'b1111111100011011001101101;
    rom[18547] = 25'b1111111100011011100010111;
    rom[18548] = 25'b1111111100011011111000010;
    rom[18549] = 25'b1111111100011100001101101;
    rom[18550] = 25'b1111111100011100100011000;
    rom[18551] = 25'b1111111100011100111000100;
    rom[18552] = 25'b1111111100011101001110000;
    rom[18553] = 25'b1111111100011101100011100;
    rom[18554] = 25'b1111111100011101111001000;
    rom[18555] = 25'b1111111100011110001110101;
    rom[18556] = 25'b1111111100011110100100010;
    rom[18557] = 25'b1111111100011110111001111;
    rom[18558] = 25'b1111111100011111001111100;
    rom[18559] = 25'b1111111100011111100101010;
    rom[18560] = 25'b1111111100011111111011000;
    rom[18561] = 25'b1111111100100000010000110;
    rom[18562] = 25'b1111111100100000100110101;
    rom[18563] = 25'b1111111100100000111100011;
    rom[18564] = 25'b1111111100100001010010010;
    rom[18565] = 25'b1111111100100001101000001;
    rom[18566] = 25'b1111111100100001111110001;
    rom[18567] = 25'b1111111100100010010100000;
    rom[18568] = 25'b1111111100100010101010000;
    rom[18569] = 25'b1111111100100011000000000;
    rom[18570] = 25'b1111111100100011010110000;
    rom[18571] = 25'b1111111100100011101100001;
    rom[18572] = 25'b1111111100100100000010010;
    rom[18573] = 25'b1111111100100100011000011;
    rom[18574] = 25'b1111111100100100101110100;
    rom[18575] = 25'b1111111100100101000100110;
    rom[18576] = 25'b1111111100100101011010111;
    rom[18577] = 25'b1111111100100101110001001;
    rom[18578] = 25'b1111111100100110000111011;
    rom[18579] = 25'b1111111100100110011101110;
    rom[18580] = 25'b1111111100100110110100001;
    rom[18581] = 25'b1111111100100111001010100;
    rom[18582] = 25'b1111111100100111100000111;
    rom[18583] = 25'b1111111100100111110111011;
    rom[18584] = 25'b1111111100101000001101110;
    rom[18585] = 25'b1111111100101000100100010;
    rom[18586] = 25'b1111111100101000111010110;
    rom[18587] = 25'b1111111100101001010001011;
    rom[18588] = 25'b1111111100101001101000000;
    rom[18589] = 25'b1111111100101001111110101;
    rom[18590] = 25'b1111111100101010010101010;
    rom[18591] = 25'b1111111100101010101011111;
    rom[18592] = 25'b1111111100101011000010101;
    rom[18593] = 25'b1111111100101011011001011;
    rom[18594] = 25'b1111111100101011110000001;
    rom[18595] = 25'b1111111100101100000110111;
    rom[18596] = 25'b1111111100101100011101110;
    rom[18597] = 25'b1111111100101100110100101;
    rom[18598] = 25'b1111111100101101001011101;
    rom[18599] = 25'b1111111100101101100010100;
    rom[18600] = 25'b1111111100101101111001011;
    rom[18601] = 25'b1111111100101110010000011;
    rom[18602] = 25'b1111111100101110100111011;
    rom[18603] = 25'b1111111100101110111110011;
    rom[18604] = 25'b1111111100101111010101100;
    rom[18605] = 25'b1111111100101111101100101;
    rom[18606] = 25'b1111111100110000000011110;
    rom[18607] = 25'b1111111100110000011010111;
    rom[18608] = 25'b1111111100110000110010001;
    rom[18609] = 25'b1111111100110001001001011;
    rom[18610] = 25'b1111111100110001100000101;
    rom[18611] = 25'b1111111100110001110111111;
    rom[18612] = 25'b1111111100110010001111010;
    rom[18613] = 25'b1111111100110010100110101;
    rom[18614] = 25'b1111111100110010111110000;
    rom[18615] = 25'b1111111100110011010101010;
    rom[18616] = 25'b1111111100110011101100110;
    rom[18617] = 25'b1111111100110100000100010;
    rom[18618] = 25'b1111111100110100011011110;
    rom[18619] = 25'b1111111100110100110011010;
    rom[18620] = 25'b1111111100110101001010110;
    rom[18621] = 25'b1111111100110101100010011;
    rom[18622] = 25'b1111111100110101111010000;
    rom[18623] = 25'b1111111100110110010001101;
    rom[18624] = 25'b1111111100110110101001011;
    rom[18625] = 25'b1111111100110111000001000;
    rom[18626] = 25'b1111111100110111011000110;
    rom[18627] = 25'b1111111100110111110000100;
    rom[18628] = 25'b1111111100111000001000011;
    rom[18629] = 25'b1111111100111000100000001;
    rom[18630] = 25'b1111111100111000111000000;
    rom[18631] = 25'b1111111100111001001111111;
    rom[18632] = 25'b1111111100111001100111110;
    rom[18633] = 25'b1111111100111001111111110;
    rom[18634] = 25'b1111111100111010010111110;
    rom[18635] = 25'b1111111100111010101111110;
    rom[18636] = 25'b1111111100111011000111110;
    rom[18637] = 25'b1111111100111011011111110;
    rom[18638] = 25'b1111111100111011110111111;
    rom[18639] = 25'b1111111100111100010000000;
    rom[18640] = 25'b1111111100111100101000001;
    rom[18641] = 25'b1111111100111101000000011;
    rom[18642] = 25'b1111111100111101011000100;
    rom[18643] = 25'b1111111100111101110000111;
    rom[18644] = 25'b1111111100111110001001000;
    rom[18645] = 25'b1111111100111110100001011;
    rom[18646] = 25'b1111111100111110111001101;
    rom[18647] = 25'b1111111100111111010010000;
    rom[18648] = 25'b1111111100111111101010011;
    rom[18649] = 25'b1111111101000000000010110;
    rom[18650] = 25'b1111111101000000011011010;
    rom[18651] = 25'b1111111101000000110011110;
    rom[18652] = 25'b1111111101000001001100001;
    rom[18653] = 25'b1111111101000001100100110;
    rom[18654] = 25'b1111111101000001111101010;
    rom[18655] = 25'b1111111101000010010101111;
    rom[18656] = 25'b1111111101000010101110100;
    rom[18657] = 25'b1111111101000011000111001;
    rom[18658] = 25'b1111111101000011011111111;
    rom[18659] = 25'b1111111101000011111000101;
    rom[18660] = 25'b1111111101000100010001011;
    rom[18661] = 25'b1111111101000100101010001;
    rom[18662] = 25'b1111111101000101000010111;
    rom[18663] = 25'b1111111101000101011011101;
    rom[18664] = 25'b1111111101000101110100100;
    rom[18665] = 25'b1111111101000110001101011;
    rom[18666] = 25'b1111111101000110100110010;
    rom[18667] = 25'b1111111101000110111111010;
    rom[18668] = 25'b1111111101000111011000010;
    rom[18669] = 25'b1111111101000111110001001;
    rom[18670] = 25'b1111111101001000001010010;
    rom[18671] = 25'b1111111101001000100011011;
    rom[18672] = 25'b1111111101001000111100011;
    rom[18673] = 25'b1111111101001001010101100;
    rom[18674] = 25'b1111111101001001101110101;
    rom[18675] = 25'b1111111101001010000111110;
    rom[18676] = 25'b1111111101001010100001000;
    rom[18677] = 25'b1111111101001010111010010;
    rom[18678] = 25'b1111111101001011010011100;
    rom[18679] = 25'b1111111101001011101100110;
    rom[18680] = 25'b1111111101001100000110001;
    rom[18681] = 25'b1111111101001100011111011;
    rom[18682] = 25'b1111111101001100111000110;
    rom[18683] = 25'b1111111101001101010010001;
    rom[18684] = 25'b1111111101001101101011101;
    rom[18685] = 25'b1111111101001110000101001;
    rom[18686] = 25'b1111111101001110011110101;
    rom[18687] = 25'b1111111101001110111000000;
    rom[18688] = 25'b1111111101001111010001100;
    rom[18689] = 25'b1111111101001111101011001;
    rom[18690] = 25'b1111111101010000000100110;
    rom[18691] = 25'b1111111101010000011110011;
    rom[18692] = 25'b1111111101010000111000000;
    rom[18693] = 25'b1111111101010001010001101;
    rom[18694] = 25'b1111111101010001101011100;
    rom[18695] = 25'b1111111101010010000101001;
    rom[18696] = 25'b1111111101010010011110111;
    rom[18697] = 25'b1111111101010010111000110;
    rom[18698] = 25'b1111111101010011010010100;
    rom[18699] = 25'b1111111101010011101100011;
    rom[18700] = 25'b1111111101010100000110010;
    rom[18701] = 25'b1111111101010100100000010;
    rom[18702] = 25'b1111111101010100111010001;
    rom[18703] = 25'b1111111101010101010100001;
    rom[18704] = 25'b1111111101010101101110001;
    rom[18705] = 25'b1111111101010110001000001;
    rom[18706] = 25'b1111111101010110100010001;
    rom[18707] = 25'b1111111101010110111100010;
    rom[18708] = 25'b1111111101010111010110011;
    rom[18709] = 25'b1111111101010111110000100;
    rom[18710] = 25'b1111111101011000001010101;
    rom[18711] = 25'b1111111101011000100100111;
    rom[18712] = 25'b1111111101011000111111001;
    rom[18713] = 25'b1111111101011001011001011;
    rom[18714] = 25'b1111111101011001110011101;
    rom[18715] = 25'b1111111101011010001110000;
    rom[18716] = 25'b1111111101011010101000010;
    rom[18717] = 25'b1111111101011011000010101;
    rom[18718] = 25'b1111111101011011011101000;
    rom[18719] = 25'b1111111101011011110111011;
    rom[18720] = 25'b1111111101011100010001111;
    rom[18721] = 25'b1111111101011100101100011;
    rom[18722] = 25'b1111111101011101000110111;
    rom[18723] = 25'b1111111101011101100001011;
    rom[18724] = 25'b1111111101011101111011111;
    rom[18725] = 25'b1111111101011110010110100;
    rom[18726] = 25'b1111111101011110110001001;
    rom[18727] = 25'b1111111101011111001011110;
    rom[18728] = 25'b1111111101011111100110011;
    rom[18729] = 25'b1111111101100000000001001;
    rom[18730] = 25'b1111111101100000011011110;
    rom[18731] = 25'b1111111101100000110110101;
    rom[18732] = 25'b1111111101100001010001010;
    rom[18733] = 25'b1111111101100001101100001;
    rom[18734] = 25'b1111111101100010000111000;
    rom[18735] = 25'b1111111101100010100001110;
    rom[18736] = 25'b1111111101100010111100110;
    rom[18737] = 25'b1111111101100011010111101;
    rom[18738] = 25'b1111111101100011110010101;
    rom[18739] = 25'b1111111101100100001101101;
    rom[18740] = 25'b1111111101100100101000100;
    rom[18741] = 25'b1111111101100101000011100;
    rom[18742] = 25'b1111111101100101011110101;
    rom[18743] = 25'b1111111101100101111001110;
    rom[18744] = 25'b1111111101100110010100110;
    rom[18745] = 25'b1111111101100110101111111;
    rom[18746] = 25'b1111111101100111001011000;
    rom[18747] = 25'b1111111101100111100110010;
    rom[18748] = 25'b1111111101101000000001100;
    rom[18749] = 25'b1111111101101000011100101;
    rom[18750] = 25'b1111111101101000110111111;
    rom[18751] = 25'b1111111101101001010011010;
    rom[18752] = 25'b1111111101101001101110101;
    rom[18753] = 25'b1111111101101010001001111;
    rom[18754] = 25'b1111111101101010100101010;
    rom[18755] = 25'b1111111101101011000000110;
    rom[18756] = 25'b1111111101101011011100001;
    rom[18757] = 25'b1111111101101011110111101;
    rom[18758] = 25'b1111111101101100010011001;
    rom[18759] = 25'b1111111101101100101110101;
    rom[18760] = 25'b1111111101101101001010001;
    rom[18761] = 25'b1111111101101101100101101;
    rom[18762] = 25'b1111111101101110000001011;
    rom[18763] = 25'b1111111101101110011100111;
    rom[18764] = 25'b1111111101101110111000100;
    rom[18765] = 25'b1111111101101111010100010;
    rom[18766] = 25'b1111111101101111101111111;
    rom[18767] = 25'b1111111101110000001011101;
    rom[18768] = 25'b1111111101110000100111011;
    rom[18769] = 25'b1111111101110001000011001;
    rom[18770] = 25'b1111111101110001011111000;
    rom[18771] = 25'b1111111101110001111010111;
    rom[18772] = 25'b1111111101110010010110101;
    rom[18773] = 25'b1111111101110010110010100;
    rom[18774] = 25'b1111111101110011001110011;
    rom[18775] = 25'b1111111101110011101010011;
    rom[18776] = 25'b1111111101110100000110011;
    rom[18777] = 25'b1111111101110100100010011;
    rom[18778] = 25'b1111111101110100111110011;
    rom[18779] = 25'b1111111101110101011010011;
    rom[18780] = 25'b1111111101110101110110011;
    rom[18781] = 25'b1111111101110110010010100;
    rom[18782] = 25'b1111111101110110101110101;
    rom[18783] = 25'b1111111101110111001010111;
    rom[18784] = 25'b1111111101110111100111000;
    rom[18785] = 25'b1111111101111000000011001;
    rom[18786] = 25'b1111111101111000011111100;
    rom[18787] = 25'b1111111101111000111011101;
    rom[18788] = 25'b1111111101111001011000000;
    rom[18789] = 25'b1111111101111001110100010;
    rom[18790] = 25'b1111111101111010010000101;
    rom[18791] = 25'b1111111101111010101101000;
    rom[18792] = 25'b1111111101111011001001011;
    rom[18793] = 25'b1111111101111011100101110;
    rom[18794] = 25'b1111111101111100000010010;
    rom[18795] = 25'b1111111101111100011110101;
    rom[18796] = 25'b1111111101111100111011001;
    rom[18797] = 25'b1111111101111101010111101;
    rom[18798] = 25'b1111111101111101110100001;
    rom[18799] = 25'b1111111101111110010000110;
    rom[18800] = 25'b1111111101111110101101010;
    rom[18801] = 25'b1111111101111111001010000;
    rom[18802] = 25'b1111111101111111100110101;
    rom[18803] = 25'b1111111110000000000011010;
    rom[18804] = 25'b1111111110000000100000000;
    rom[18805] = 25'b1111111110000000111100101;
    rom[18806] = 25'b1111111110000001011001011;
    rom[18807] = 25'b1111111110000001110110001;
    rom[18808] = 25'b1111111110000010010011000;
    rom[18809] = 25'b1111111110000010101111110;
    rom[18810] = 25'b1111111110000011001100101;
    rom[18811] = 25'b1111111110000011101001100;
    rom[18812] = 25'b1111111110000100000110100;
    rom[18813] = 25'b1111111110000100100011010;
    rom[18814] = 25'b1111111110000101000000010;
    rom[18815] = 25'b1111111110000101011101010;
    rom[18816] = 25'b1111111110000101111010010;
    rom[18817] = 25'b1111111110000110010111010;
    rom[18818] = 25'b1111111110000110110100011;
    rom[18819] = 25'b1111111110000111010001011;
    rom[18820] = 25'b1111111110000111101110100;
    rom[18821] = 25'b1111111110001000001011101;
    rom[18822] = 25'b1111111110001000101000110;
    rom[18823] = 25'b1111111110001001000101111;
    rom[18824] = 25'b1111111110001001100011001;
    rom[18825] = 25'b1111111110001010000000011;
    rom[18826] = 25'b1111111110001010011101101;
    rom[18827] = 25'b1111111110001010111010111;
    rom[18828] = 25'b1111111110001011011000010;
    rom[18829] = 25'b1111111110001011110101101;
    rom[18830] = 25'b1111111110001100010010111;
    rom[18831] = 25'b1111111110001100110000011;
    rom[18832] = 25'b1111111110001101001101101;
    rom[18833] = 25'b1111111110001101101011001;
    rom[18834] = 25'b1111111110001110001000101;
    rom[18835] = 25'b1111111110001110100110001;
    rom[18836] = 25'b1111111110001111000011100;
    rom[18837] = 25'b1111111110001111100001001;
    rom[18838] = 25'b1111111110001111111110101;
    rom[18839] = 25'b1111111110010000011100010;
    rom[18840] = 25'b1111111110010000111001111;
    rom[18841] = 25'b1111111110010001010111011;
    rom[18842] = 25'b1111111110010001110101000;
    rom[18843] = 25'b1111111110010010010010110;
    rom[18844] = 25'b1111111110010010110000011;
    rom[18845] = 25'b1111111110010011001110001;
    rom[18846] = 25'b1111111110010011101011111;
    rom[18847] = 25'b1111111110010100001001110;
    rom[18848] = 25'b1111111110010100100111100;
    rom[18849] = 25'b1111111110010101000101010;
    rom[18850] = 25'b1111111110010101100011001;
    rom[18851] = 25'b1111111110010110000001000;
    rom[18852] = 25'b1111111110010110011110111;
    rom[18853] = 25'b1111111110010110111100111;
    rom[18854] = 25'b1111111110010111011010110;
    rom[18855] = 25'b1111111110010111111000110;
    rom[18856] = 25'b1111111110011000010110110;
    rom[18857] = 25'b1111111110011000110100110;
    rom[18858] = 25'b1111111110011001010010110;
    rom[18859] = 25'b1111111110011001110000111;
    rom[18860] = 25'b1111111110011010001111000;
    rom[18861] = 25'b1111111110011010101101000;
    rom[18862] = 25'b1111111110011011001011001;
    rom[18863] = 25'b1111111110011011101001011;
    rom[18864] = 25'b1111111110011100000111100;
    rom[18865] = 25'b1111111110011100100101110;
    rom[18866] = 25'b1111111110011101000011111;
    rom[18867] = 25'b1111111110011101100010001;
    rom[18868] = 25'b1111111110011110000000100;
    rom[18869] = 25'b1111111110011110011110110;
    rom[18870] = 25'b1111111110011110111101001;
    rom[18871] = 25'b1111111110011111011011100;
    rom[18872] = 25'b1111111110011111111001111;
    rom[18873] = 25'b1111111110100000011000010;
    rom[18874] = 25'b1111111110100000110110101;
    rom[18875] = 25'b1111111110100001010101001;
    rom[18876] = 25'b1111111110100001110011101;
    rom[18877] = 25'b1111111110100010010010001;
    rom[18878] = 25'b1111111110100010110000101;
    rom[18879] = 25'b1111111110100011001111001;
    rom[18880] = 25'b1111111110100011101101101;
    rom[18881] = 25'b1111111110100100001100010;
    rom[18882] = 25'b1111111110100100101010111;
    rom[18883] = 25'b1111111110100101001001101;
    rom[18884] = 25'b1111111110100101101000010;
    rom[18885] = 25'b1111111110100110000110111;
    rom[18886] = 25'b1111111110100110100101100;
    rom[18887] = 25'b1111111110100111000100010;
    rom[18888] = 25'b1111111110100111100011001;
    rom[18889] = 25'b1111111110101000000001111;
    rom[18890] = 25'b1111111110101000100000101;
    rom[18891] = 25'b1111111110101000111111100;
    rom[18892] = 25'b1111111110101001011110010;
    rom[18893] = 25'b1111111110101001111101001;
    rom[18894] = 25'b1111111110101010011100001;
    rom[18895] = 25'b1111111110101010111011000;
    rom[18896] = 25'b1111111110101011011001111;
    rom[18897] = 25'b1111111110101011111000111;
    rom[18898] = 25'b1111111110101100010111111;
    rom[18899] = 25'b1111111110101100110110111;
    rom[18900] = 25'b1111111110101101010101111;
    rom[18901] = 25'b1111111110101101110101000;
    rom[18902] = 25'b1111111110101110010100000;
    rom[18903] = 25'b1111111110101110110011000;
    rom[18904] = 25'b1111111110101111010010010;
    rom[18905] = 25'b1111111110101111110001011;
    rom[18906] = 25'b1111111110110000010000100;
    rom[18907] = 25'b1111111110110000101111110;
    rom[18908] = 25'b1111111110110001001110111;
    rom[18909] = 25'b1111111110110001101110001;
    rom[18910] = 25'b1111111110110010001101011;
    rom[18911] = 25'b1111111110110010101100101;
    rom[18912] = 25'b1111111110110011001100000;
    rom[18913] = 25'b1111111110110011101011011;
    rom[18914] = 25'b1111111110110100001010101;
    rom[18915] = 25'b1111111110110100101010000;
    rom[18916] = 25'b1111111110110101001001011;
    rom[18917] = 25'b1111111110110101101000111;
    rom[18918] = 25'b1111111110110110001000010;
    rom[18919] = 25'b1111111110110110100111110;
    rom[18920] = 25'b1111111110110111000111001;
    rom[18921] = 25'b1111111110110111100110101;
    rom[18922] = 25'b1111111110111000000110010;
    rom[18923] = 25'b1111111110111000100101110;
    rom[18924] = 25'b1111111110111001000101011;
    rom[18925] = 25'b1111111110111001100100111;
    rom[18926] = 25'b1111111110111010000100100;
    rom[18927] = 25'b1111111110111010100100001;
    rom[18928] = 25'b1111111110111011000011110;
    rom[18929] = 25'b1111111110111011100011011;
    rom[18930] = 25'b1111111110111100000011001;
    rom[18931] = 25'b1111111110111100100010111;
    rom[18932] = 25'b1111111110111101000010101;
    rom[18933] = 25'b1111111110111101100010011;
    rom[18934] = 25'b1111111110111110000010010;
    rom[18935] = 25'b1111111110111110100010000;
    rom[18936] = 25'b1111111110111111000001110;
    rom[18937] = 25'b1111111110111111100001101;
    rom[18938] = 25'b1111111111000000000001100;
    rom[18939] = 25'b1111111111000000100001011;
    rom[18940] = 25'b1111111111000001000001011;
    rom[18941] = 25'b1111111111000001100001010;
    rom[18942] = 25'b1111111111000010000001010;
    rom[18943] = 25'b1111111111000010100001001;
    rom[18944] = 25'b1111111111000011000001010;
    rom[18945] = 25'b1111111111000011100001010;
    rom[18946] = 25'b1111111111000100000001010;
    rom[18947] = 25'b1111111111000100100001010;
    rom[18948] = 25'b1111111111000101000001011;
    rom[18949] = 25'b1111111111000101100001100;
    rom[18950] = 25'b1111111111000110000001101;
    rom[18951] = 25'b1111111111000110100001110;
    rom[18952] = 25'b1111111111000111000010000;
    rom[18953] = 25'b1111111111000111100010001;
    rom[18954] = 25'b1111111111001000000010011;
    rom[18955] = 25'b1111111111001000100010101;
    rom[18956] = 25'b1111111111001001000010111;
    rom[18957] = 25'b1111111111001001100011001;
    rom[18958] = 25'b1111111111001010000011011;
    rom[18959] = 25'b1111111111001010100011110;
    rom[18960] = 25'b1111111111001011000100001;
    rom[18961] = 25'b1111111111001011100100100;
    rom[18962] = 25'b1111111111001100000100111;
    rom[18963] = 25'b1111111111001100100101010;
    rom[18964] = 25'b1111111111001101000101101;
    rom[18965] = 25'b1111111111001101100110001;
    rom[18966] = 25'b1111111111001110000110101;
    rom[18967] = 25'b1111111111001110100111001;
    rom[18968] = 25'b1111111111001111000111101;
    rom[18969] = 25'b1111111111001111101000001;
    rom[18970] = 25'b1111111111010000001000101;
    rom[18971] = 25'b1111111111010000101001001;
    rom[18972] = 25'b1111111111010001001001110;
    rom[18973] = 25'b1111111111010001101010011;
    rom[18974] = 25'b1111111111010010001011000;
    rom[18975] = 25'b1111111111010010101011101;
    rom[18976] = 25'b1111111111010011001100010;
    rom[18977] = 25'b1111111111010011101101000;
    rom[18978] = 25'b1111111111010100001101101;
    rom[18979] = 25'b1111111111010100101110100;
    rom[18980] = 25'b1111111111010101001111010;
    rom[18981] = 25'b1111111111010101110000000;
    rom[18982] = 25'b1111111111010110010000110;
    rom[18983] = 25'b1111111111010110110001101;
    rom[18984] = 25'b1111111111010111010010011;
    rom[18985] = 25'b1111111111010111110011010;
    rom[18986] = 25'b1111111111011000010100001;
    rom[18987] = 25'b1111111111011000110101000;
    rom[18988] = 25'b1111111111011001010101111;
    rom[18989] = 25'b1111111111011001110110110;
    rom[18990] = 25'b1111111111011010010111110;
    rom[18991] = 25'b1111111111011010111000110;
    rom[18992] = 25'b1111111111011011011001110;
    rom[18993] = 25'b1111111111011011111010110;
    rom[18994] = 25'b1111111111011100011011111;
    rom[18995] = 25'b1111111111011100111100110;
    rom[18996] = 25'b1111111111011101011101111;
    rom[18997] = 25'b1111111111011101111111000;
    rom[18998] = 25'b1111111111011110100000000;
    rom[18999] = 25'b1111111111011111000001010;
    rom[19000] = 25'b1111111111011111100010011;
    rom[19001] = 25'b1111111111100000000011100;
    rom[19002] = 25'b1111111111100000100100101;
    rom[19003] = 25'b1111111111100001000101111;
    rom[19004] = 25'b1111111111100001100111001;
    rom[19005] = 25'b1111111111100010001000011;
    rom[19006] = 25'b1111111111100010101001101;
    rom[19007] = 25'b1111111111100011001010111;
    rom[19008] = 25'b1111111111100011101100010;
    rom[19009] = 25'b1111111111100100001101100;
    rom[19010] = 25'b1111111111100100101110111;
    rom[19011] = 25'b1111111111100101010000001;
    rom[19012] = 25'b1111111111100101110001101;
    rom[19013] = 25'b1111111111100110010010111;
    rom[19014] = 25'b1111111111100110110100011;
    rom[19015] = 25'b1111111111100111010101110;
    rom[19016] = 25'b1111111111100111110111010;
    rom[19017] = 25'b1111111111101000011000110;
    rom[19018] = 25'b1111111111101000111010001;
    rom[19019] = 25'b1111111111101001011011110;
    rom[19020] = 25'b1111111111101001111101010;
    rom[19021] = 25'b1111111111101010011110110;
    rom[19022] = 25'b1111111111101011000000011;
    rom[19023] = 25'b1111111111101011100001111;
    rom[19024] = 25'b1111111111101100000011100;
    rom[19025] = 25'b1111111111101100100101001;
    rom[19026] = 25'b1111111111101101000110110;
    rom[19027] = 25'b1111111111101101101000100;
    rom[19028] = 25'b1111111111101110001010001;
    rom[19029] = 25'b1111111111101110101011110;
    rom[19030] = 25'b1111111111101111001101100;
    rom[19031] = 25'b1111111111101111101111010;
    rom[19032] = 25'b1111111111110000010001000;
    rom[19033] = 25'b1111111111110000110010110;
    rom[19034] = 25'b1111111111110001010100100;
    rom[19035] = 25'b1111111111110001110110011;
    rom[19036] = 25'b1111111111110010011000001;
    rom[19037] = 25'b1111111111110010111010000;
    rom[19038] = 25'b1111111111110011011011111;
    rom[19039] = 25'b1111111111110011111101101;
    rom[19040] = 25'b1111111111110100011111101;
    rom[19041] = 25'b1111111111110101000001100;
    rom[19042] = 25'b1111111111110101100011100;
    rom[19043] = 25'b1111111111110110000101011;
    rom[19044] = 25'b1111111111110110100111011;
    rom[19045] = 25'b1111111111110111001001011;
    rom[19046] = 25'b1111111111110111101011011;
    rom[19047] = 25'b1111111111111000001101011;
    rom[19048] = 25'b1111111111111000101111011;
    rom[19049] = 25'b1111111111111001010001011;
    rom[19050] = 25'b1111111111111001110011100;
    rom[19051] = 25'b1111111111111010010101101;
    rom[19052] = 25'b1111111111111010110111101;
    rom[19053] = 25'b1111111111111011011001110;
    rom[19054] = 25'b1111111111111011111100000;
    rom[19055] = 25'b1111111111111100011110001;
    rom[19056] = 25'b1111111111111101000000010;
    rom[19057] = 25'b1111111111111101100010100;
    rom[19058] = 25'b1111111111111110000100101;
    rom[19059] = 25'b1111111111111110100110111;
    rom[19060] = 25'b1111111111111111001001001;
    rom[19061] = 25'b1111111111111111101011011;
    rom[19062] = 25'b0000000000000000001101101;
    rom[19063] = 25'b0000000000000000101111111;
    rom[19064] = 25'b0000000000000001010010010;
    rom[19065] = 25'b0000000000000001110100100;
    rom[19066] = 25'b0000000000000010010110111;
    rom[19067] = 25'b0000000000000010111001010;
    rom[19068] = 25'b0000000000000011011011101;
    rom[19069] = 25'b0000000000000011111110000;
    rom[19070] = 25'b0000000000000100100000011;
    rom[19071] = 25'b0000000000000101000010110;
    rom[19072] = 25'b0000000000000101100101010;
    rom[19073] = 25'b0000000000000110000111110;
    rom[19074] = 25'b0000000000000110101010001;
    rom[19075] = 25'b0000000000000111001100110;
    rom[19076] = 25'b0000000000000111101111001;
    rom[19077] = 25'b0000000000001000010001110;
    rom[19078] = 25'b0000000000001000110100010;
    rom[19079] = 25'b0000000000001001010110111;
    rom[19080] = 25'b0000000000001001111001011;
    rom[19081] = 25'b0000000000001010011100000;
    rom[19082] = 25'b0000000000001010111110101;
    rom[19083] = 25'b0000000000001011100001010;
    rom[19084] = 25'b0000000000001100000011111;
    rom[19085] = 25'b0000000000001100100110100;
    rom[19086] = 25'b0000000000001101001001001;
    rom[19087] = 25'b0000000000001101101011111;
    rom[19088] = 25'b0000000000001110001110100;
    rom[19089] = 25'b0000000000001110110001010;
    rom[19090] = 25'b0000000000001111010100000;
    rom[19091] = 25'b0000000000001111110110110;
    rom[19092] = 25'b0000000000010000011001101;
    rom[19093] = 25'b0000000000010000111100011;
    rom[19094] = 25'b0000000000010001011111001;
    rom[19095] = 25'b0000000000010010000010000;
    rom[19096] = 25'b0000000000010010100100111;
    rom[19097] = 25'b0000000000010011000111101;
    rom[19098] = 25'b0000000000010011101010100;
    rom[19099] = 25'b0000000000010100001101100;
    rom[19100] = 25'b0000000000010100110000010;
    rom[19101] = 25'b0000000000010101010011010;
    rom[19102] = 25'b0000000000010101110110001;
    rom[19103] = 25'b0000000000010110011001000;
    rom[19104] = 25'b0000000000010110111100001;
    rom[19105] = 25'b0000000000010111011111000;
    rom[19106] = 25'b0000000000011000000010000;
    rom[19107] = 25'b0000000000011000100101000;
    rom[19108] = 25'b0000000000011001001000000;
    rom[19109] = 25'b0000000000011001101011001;
    rom[19110] = 25'b0000000000011010001110001;
    rom[19111] = 25'b0000000000011010110001001;
    rom[19112] = 25'b0000000000011011010100010;
    rom[19113] = 25'b0000000000011011110111011;
    rom[19114] = 25'b0000000000011100011010100;
    rom[19115] = 25'b0000000000011100111101101;
    rom[19116] = 25'b0000000000011101100000110;
    rom[19117] = 25'b0000000000011110000011110;
    rom[19118] = 25'b0000000000011110100111000;
    rom[19119] = 25'b0000000000011111001010010;
    rom[19120] = 25'b0000000000011111101101011;
    rom[19121] = 25'b0000000000100000010000101;
    rom[19122] = 25'b0000000000100000110011111;
    rom[19123] = 25'b0000000000100001010111000;
    rom[19124] = 25'b0000000000100001111010011;
    rom[19125] = 25'b0000000000100010011101100;
    rom[19126] = 25'b0000000000100011000000111;
    rom[19127] = 25'b0000000000100011100100001;
    rom[19128] = 25'b0000000000100100000111100;
    rom[19129] = 25'b0000000000100100101010111;
    rom[19130] = 25'b0000000000100101001110001;
    rom[19131] = 25'b0000000000100101110001100;
    rom[19132] = 25'b0000000000100110010100111;
    rom[19133] = 25'b0000000000100110111000010;
    rom[19134] = 25'b0000000000100111011011101;
    rom[19135] = 25'b0000000000100111111111001;
    rom[19136] = 25'b0000000000101000100010100;
    rom[19137] = 25'b0000000000101001000101111;
    rom[19138] = 25'b0000000000101001101001011;
    rom[19139] = 25'b0000000000101010001100111;
    rom[19140] = 25'b0000000000101010110000011;
    rom[19141] = 25'b0000000000101011010011111;
    rom[19142] = 25'b0000000000101011110111011;
    rom[19143] = 25'b0000000000101100011010111;
    rom[19144] = 25'b0000000000101100111110011;
    rom[19145] = 25'b0000000000101101100010000;
    rom[19146] = 25'b0000000000101110000101101;
    rom[19147] = 25'b0000000000101110101001001;
    rom[19148] = 25'b0000000000101111001100110;
    rom[19149] = 25'b0000000000101111110000010;
    rom[19150] = 25'b0000000000110000010011111;
    rom[19151] = 25'b0000000000110000110111100;
    rom[19152] = 25'b0000000000110001011011010;
    rom[19153] = 25'b0000000000110001111110111;
    rom[19154] = 25'b0000000000110010100010100;
    rom[19155] = 25'b0000000000110011000110010;
    rom[19156] = 25'b0000000000110011101001111;
    rom[19157] = 25'b0000000000110100001101101;
    rom[19158] = 25'b0000000000110100110001011;
    rom[19159] = 25'b0000000000110101010101001;
    rom[19160] = 25'b0000000000110101111000111;
    rom[19161] = 25'b0000000000110110011100101;
    rom[19162] = 25'b0000000000110111000000011;
    rom[19163] = 25'b0000000000110111100100010;
    rom[19164] = 25'b0000000000111000001000000;
    rom[19165] = 25'b0000000000111000101011111;
    rom[19166] = 25'b0000000000111001001111101;
    rom[19167] = 25'b0000000000111001110011100;
    rom[19168] = 25'b0000000000111010010111011;
    rom[19169] = 25'b0000000000111010111011001;
    rom[19170] = 25'b0000000000111011011111000;
    rom[19171] = 25'b0000000000111100000010111;
    rom[19172] = 25'b0000000000111100100110111;
    rom[19173] = 25'b0000000000111101001010111;
    rom[19174] = 25'b0000000000111101101110101;
    rom[19175] = 25'b0000000000111110010010101;
    rom[19176] = 25'b0000000000111110110110101;
    rom[19177] = 25'b0000000000111111011010100;
    rom[19178] = 25'b0000000000111111111110100;
    rom[19179] = 25'b0000000001000000100010100;
    rom[19180] = 25'b0000000001000001000110100;
    rom[19181] = 25'b0000000001000001101010100;
    rom[19182] = 25'b0000000001000010001110101;
    rom[19183] = 25'b0000000001000010110010101;
    rom[19184] = 25'b0000000001000011010110101;
    rom[19185] = 25'b0000000001000011111010110;
    rom[19186] = 25'b0000000001000100011110110;
    rom[19187] = 25'b0000000001000101000010111;
    rom[19188] = 25'b0000000001000101100111000;
    rom[19189] = 25'b0000000001000110001011001;
    rom[19190] = 25'b0000000001000110101111001;
    rom[19191] = 25'b0000000001000111010011010;
    rom[19192] = 25'b0000000001000111110111011;
    rom[19193] = 25'b0000000001001000011011101;
    rom[19194] = 25'b0000000001001000111111110;
    rom[19195] = 25'b0000000001001001100100000;
    rom[19196] = 25'b0000000001001010001000001;
    rom[19197] = 25'b0000000001001010101100011;
    rom[19198] = 25'b0000000001001011010000100;
    rom[19199] = 25'b0000000001001011110100110;
    rom[19200] = 25'b0000000001001100011001000;
    rom[19201] = 25'b0000000001001100111101010;
    rom[19202] = 25'b0000000001001101100001100;
    rom[19203] = 25'b0000000001001110000101111;
    rom[19204] = 25'b0000000001001110101010000;
    rom[19205] = 25'b0000000001001111001110011;
    rom[19206] = 25'b0000000001001111110010110;
    rom[19207] = 25'b0000000001010000010111000;
    rom[19208] = 25'b0000000001010000111011010;
    rom[19209] = 25'b0000000001010001011111110;
    rom[19210] = 25'b0000000001010010000100000;
    rom[19211] = 25'b0000000001010010101000011;
    rom[19212] = 25'b0000000001010011001100101;
    rom[19213] = 25'b0000000001010011110001001;
    rom[19214] = 25'b0000000001010100010101100;
    rom[19215] = 25'b0000000001010100111001111;
    rom[19216] = 25'b0000000001010101011110010;
    rom[19217] = 25'b0000000001010110000010110;
    rom[19218] = 25'b0000000001010110100111001;
    rom[19219] = 25'b0000000001010111001011100;
    rom[19220] = 25'b0000000001010111110000000;
    rom[19221] = 25'b0000000001011000010100100;
    rom[19222] = 25'b0000000001011000111001000;
    rom[19223] = 25'b0000000001011001011101011;
    rom[19224] = 25'b0000000001011010000001111;
    rom[19225] = 25'b0000000001011010100110011;
    rom[19226] = 25'b0000000001011011001011000;
    rom[19227] = 25'b0000000001011011101111100;
    rom[19228] = 25'b0000000001011100010100000;
    rom[19229] = 25'b0000000001011100111000101;
    rom[19230] = 25'b0000000001011101011101001;
    rom[19231] = 25'b0000000001011110000001101;
    rom[19232] = 25'b0000000001011110100110010;
    rom[19233] = 25'b0000000001011111001010111;
    rom[19234] = 25'b0000000001011111101111011;
    rom[19235] = 25'b0000000001100000010100000;
    rom[19236] = 25'b0000000001100000111000100;
    rom[19237] = 25'b0000000001100001011101010;
    rom[19238] = 25'b0000000001100010000001111;
    rom[19239] = 25'b0000000001100010100110100;
    rom[19240] = 25'b0000000001100011001011001;
    rom[19241] = 25'b0000000001100011101111110;
    rom[19242] = 25'b0000000001100100010100100;
    rom[19243] = 25'b0000000001100100111001001;
    rom[19244] = 25'b0000000001100101011101110;
    rom[19245] = 25'b0000000001100110000010100;
    rom[19246] = 25'b0000000001100110100111010;
    rom[19247] = 25'b0000000001100111001011111;
    rom[19248] = 25'b0000000001100111110000110;
    rom[19249] = 25'b0000000001101000010101011;
    rom[19250] = 25'b0000000001101000111010001;
    rom[19251] = 25'b0000000001101001011110111;
    rom[19252] = 25'b0000000001101010000011101;
    rom[19253] = 25'b0000000001101010101000011;
    rom[19254] = 25'b0000000001101011001101001;
    rom[19255] = 25'b0000000001101011110010000;
    rom[19256] = 25'b0000000001101100010110110;
    rom[19257] = 25'b0000000001101100111011100;
    rom[19258] = 25'b0000000001101101100000011;
    rom[19259] = 25'b0000000001101110000101001;
    rom[19260] = 25'b0000000001101110101010000;
    rom[19261] = 25'b0000000001101111001110111;
    rom[19262] = 25'b0000000001101111110011101;
    rom[19263] = 25'b0000000001110000011000100;
    rom[19264] = 25'b0000000001110000111101011;
    rom[19265] = 25'b0000000001110001100010010;
    rom[19266] = 25'b0000000001110010000111001;
    rom[19267] = 25'b0000000001110010101100000;
    rom[19268] = 25'b0000000001110011010000111;
    rom[19269] = 25'b0000000001110011110101110;
    rom[19270] = 25'b0000000001110100011010110;
    rom[19271] = 25'b0000000001110100111111101;
    rom[19272] = 25'b0000000001110101100100100;
    rom[19273] = 25'b0000000001110110001001100;
    rom[19274] = 25'b0000000001110110101110011;
    rom[19275] = 25'b0000000001110111010011011;
    rom[19276] = 25'b0000000001110111111000011;
    rom[19277] = 25'b0000000001111000011101010;
    rom[19278] = 25'b0000000001111001000010010;
    rom[19279] = 25'b0000000001111001100111001;
    rom[19280] = 25'b0000000001111010001100001;
    rom[19281] = 25'b0000000001111010110001001;
    rom[19282] = 25'b0000000001111011010110010;
    rom[19283] = 25'b0000000001111011111011010;
    rom[19284] = 25'b0000000001111100100000001;
    rom[19285] = 25'b0000000001111101000101010;
    rom[19286] = 25'b0000000001111101101010010;
    rom[19287] = 25'b0000000001111110001111011;
    rom[19288] = 25'b0000000001111110110100011;
    rom[19289] = 25'b0000000001111111011001011;
    rom[19290] = 25'b0000000001111111111110100;
    rom[19291] = 25'b0000000010000000100011100;
    rom[19292] = 25'b0000000010000001001000101;
    rom[19293] = 25'b0000000010000001101101101;
    rom[19294] = 25'b0000000010000010010010110;
    rom[19295] = 25'b0000000010000010110111111;
    rom[19296] = 25'b0000000010000011011101000;
    rom[19297] = 25'b0000000010000100000010000;
    rom[19298] = 25'b0000000010000100100111001;
    rom[19299] = 25'b0000000010000101001100010;
    rom[19300] = 25'b0000000010000101110001011;
    rom[19301] = 25'b0000000010000110010110100;
    rom[19302] = 25'b0000000010000110111011110;
    rom[19303] = 25'b0000000010000111100000110;
    rom[19304] = 25'b0000000010001000000110000;
    rom[19305] = 25'b0000000010001000101011001;
    rom[19306] = 25'b0000000010001001010000010;
    rom[19307] = 25'b0000000010001001110101100;
    rom[19308] = 25'b0000000010001010011010101;
    rom[19309] = 25'b0000000010001010111111110;
    rom[19310] = 25'b0000000010001011100101000;
    rom[19311] = 25'b0000000010001100001010010;
    rom[19312] = 25'b0000000010001100101111011;
    rom[19313] = 25'b0000000010001101010100101;
    rom[19314] = 25'b0000000010001101111001111;
    rom[19315] = 25'b0000000010001110011111001;
    rom[19316] = 25'b0000000010001111000100010;
    rom[19317] = 25'b0000000010001111101001100;
    rom[19318] = 25'b0000000010010000001110101;
    rom[19319] = 25'b0000000010010000110100000;
    rom[19320] = 25'b0000000010010001011001010;
    rom[19321] = 25'b0000000010010001111110100;
    rom[19322] = 25'b0000000010010010100011110;
    rom[19323] = 25'b0000000010010011001001000;
    rom[19324] = 25'b0000000010010011101110010;
    rom[19325] = 25'b0000000010010100010011100;
    rom[19326] = 25'b0000000010010100111000110;
    rom[19327] = 25'b0000000010010101011110001;
    rom[19328] = 25'b0000000010010110000011011;
    rom[19329] = 25'b0000000010010110101000101;
    rom[19330] = 25'b0000000010010111001110000;
    rom[19331] = 25'b0000000010010111110011010;
    rom[19332] = 25'b0000000010011000011000101;
    rom[19333] = 25'b0000000010011000111101111;
    rom[19334] = 25'b0000000010011001100011010;
    rom[19335] = 25'b0000000010011010001000100;
    rom[19336] = 25'b0000000010011010101101111;
    rom[19337] = 25'b0000000010011011010011010;
    rom[19338] = 25'b0000000010011011111000101;
    rom[19339] = 25'b0000000010011100011101111;
    rom[19340] = 25'b0000000010011101000011010;
    rom[19341] = 25'b0000000010011101101000101;
    rom[19342] = 25'b0000000010011110001110000;
    rom[19343] = 25'b0000000010011110110011011;
    rom[19344] = 25'b0000000010011111011000110;
    rom[19345] = 25'b0000000010011111111110000;
    rom[19346] = 25'b0000000010100000100011011;
    rom[19347] = 25'b0000000010100001001000110;
    rom[19348] = 25'b0000000010100001101110010;
    rom[19349] = 25'b0000000010100010010011100;
    rom[19350] = 25'b0000000010100010111000111;
    rom[19351] = 25'b0000000010100011011110011;
    rom[19352] = 25'b0000000010100100000011110;
    rom[19353] = 25'b0000000010100100101001001;
    rom[19354] = 25'b0000000010100101001110100;
    rom[19355] = 25'b0000000010100101110100000;
    rom[19356] = 25'b0000000010100110011001011;
    rom[19357] = 25'b0000000010100110111110110;
    rom[19358] = 25'b0000000010100111100100010;
    rom[19359] = 25'b0000000010101000001001101;
    rom[19360] = 25'b0000000010101000101111001;
    rom[19361] = 25'b0000000010101001010100100;
    rom[19362] = 25'b0000000010101001111001111;
    rom[19363] = 25'b0000000010101010011111011;
    rom[19364] = 25'b0000000010101011000100111;
    rom[19365] = 25'b0000000010101011101010010;
    rom[19366] = 25'b0000000010101100001111110;
    rom[19367] = 25'b0000000010101100110101001;
    rom[19368] = 25'b0000000010101101011010101;
    rom[19369] = 25'b0000000010101110000000000;
    rom[19370] = 25'b0000000010101110100101100;
    rom[19371] = 25'b0000000010101111001011000;
    rom[19372] = 25'b0000000010101111110000100;
    rom[19373] = 25'b0000000010110000010110000;
    rom[19374] = 25'b0000000010110000111011011;
    rom[19375] = 25'b0000000010110001100000111;
    rom[19376] = 25'b0000000010110010000110011;
    rom[19377] = 25'b0000000010110010101011111;
    rom[19378] = 25'b0000000010110011010001011;
    rom[19379] = 25'b0000000010110011110110111;
    rom[19380] = 25'b0000000010110100011100011;
    rom[19381] = 25'b0000000010110101000001110;
    rom[19382] = 25'b0000000010110101100111011;
    rom[19383] = 25'b0000000010110110001100110;
    rom[19384] = 25'b0000000010110110110010011;
    rom[19385] = 25'b0000000010110111010111110;
    rom[19386] = 25'b0000000010110111111101011;
    rom[19387] = 25'b0000000010111000100010110;
    rom[19388] = 25'b0000000010111001001000011;
    rom[19389] = 25'b0000000010111001101101111;
    rom[19390] = 25'b0000000010111010010011010;
    rom[19391] = 25'b0000000010111010111000111;
    rom[19392] = 25'b0000000010111011011110011;
    rom[19393] = 25'b0000000010111100000011111;
    rom[19394] = 25'b0000000010111100101001011;
    rom[19395] = 25'b0000000010111101001110111;
    rom[19396] = 25'b0000000010111101110100100;
    rom[19397] = 25'b0000000010111110011010000;
    rom[19398] = 25'b0000000010111110111111100;
    rom[19399] = 25'b0000000010111111100101001;
    rom[19400] = 25'b0000000011000000001010100;
    rom[19401] = 25'b0000000011000000110000001;
    rom[19402] = 25'b0000000011000001010101101;
    rom[19403] = 25'b0000000011000001111011001;
    rom[19404] = 25'b0000000011000010100000110;
    rom[19405] = 25'b0000000011000011000110010;
    rom[19406] = 25'b0000000011000011101011110;
    rom[19407] = 25'b0000000011000100010001011;
    rom[19408] = 25'b0000000011000100110110111;
    rom[19409] = 25'b0000000011000101011100011;
    rom[19410] = 25'b0000000011000110000010000;
    rom[19411] = 25'b0000000011000110100111100;
    rom[19412] = 25'b0000000011000111001101000;
    rom[19413] = 25'b0000000011000111110010101;
    rom[19414] = 25'b0000000011001000011000001;
    rom[19415] = 25'b0000000011001000111101101;
    rom[19416] = 25'b0000000011001001100011010;
    rom[19417] = 25'b0000000011001010001000110;
    rom[19418] = 25'b0000000011001010101110011;
    rom[19419] = 25'b0000000011001011010011111;
    rom[19420] = 25'b0000000011001011111001100;
    rom[19421] = 25'b0000000011001100011111000;
    rom[19422] = 25'b0000000011001101000100100;
    rom[19423] = 25'b0000000011001101101010001;
    rom[19424] = 25'b0000000011001110001111101;
    rom[19425] = 25'b0000000011001110110101001;
    rom[19426] = 25'b0000000011001111011010110;
    rom[19427] = 25'b0000000011010000000000010;
    rom[19428] = 25'b0000000011010000100101111;
    rom[19429] = 25'b0000000011010001001011011;
    rom[19430] = 25'b0000000011010001110001000;
    rom[19431] = 25'b0000000011010010010110100;
    rom[19432] = 25'b0000000011010010111100000;
    rom[19433] = 25'b0000000011010011100001101;
    rom[19434] = 25'b0000000011010100000111001;
    rom[19435] = 25'b0000000011010100101100101;
    rom[19436] = 25'b0000000011010101010010011;
    rom[19437] = 25'b0000000011010101110111111;
    rom[19438] = 25'b0000000011010110011101011;
    rom[19439] = 25'b0000000011010111000011000;
    rom[19440] = 25'b0000000011010111101000100;
    rom[19441] = 25'b0000000011011000001110000;
    rom[19442] = 25'b0000000011011000110011101;
    rom[19443] = 25'b0000000011011001011001001;
    rom[19444] = 25'b0000000011011001111110101;
    rom[19445] = 25'b0000000011011010100100010;
    rom[19446] = 25'b0000000011011011001001110;
    rom[19447] = 25'b0000000011011011101111010;
    rom[19448] = 25'b0000000011011100010100111;
    rom[19449] = 25'b0000000011011100111010011;
    rom[19450] = 25'b0000000011011101011111111;
    rom[19451] = 25'b0000000011011110000101100;
    rom[19452] = 25'b0000000011011110101011000;
    rom[19453] = 25'b0000000011011111010000100;
    rom[19454] = 25'b0000000011011111110110001;
    rom[19455] = 25'b0000000011100000011011101;
    rom[19456] = 25'b0000000011100001000001001;
    rom[19457] = 25'b0000000011100001100110110;
    rom[19458] = 25'b0000000011100010001100010;
    rom[19459] = 25'b0000000011100010110001110;
    rom[19460] = 25'b0000000011100011010111011;
    rom[19461] = 25'b0000000011100011111100110;
    rom[19462] = 25'b0000000011100100100010010;
    rom[19463] = 25'b0000000011100101000111111;
    rom[19464] = 25'b0000000011100101101101011;
    rom[19465] = 25'b0000000011100110010010111;
    rom[19466] = 25'b0000000011100110111000011;
    rom[19467] = 25'b0000000011100111011101111;
    rom[19468] = 25'b0000000011101000000011100;
    rom[19469] = 25'b0000000011101000101000111;
    rom[19470] = 25'b0000000011101001001110100;
    rom[19471] = 25'b0000000011101001110100000;
    rom[19472] = 25'b0000000011101010011001100;
    rom[19473] = 25'b0000000011101010111111000;
    rom[19474] = 25'b0000000011101011100100011;
    rom[19475] = 25'b0000000011101100001010000;
    rom[19476] = 25'b0000000011101100101111011;
    rom[19477] = 25'b0000000011101101010101000;
    rom[19478] = 25'b0000000011101101111010011;
    rom[19479] = 25'b0000000011101110100000000;
    rom[19480] = 25'b0000000011101111000101011;
    rom[19481] = 25'b0000000011101111101011000;
    rom[19482] = 25'b0000000011110000010000011;
    rom[19483] = 25'b0000000011110000110101111;
    rom[19484] = 25'b0000000011110001011011010;
    rom[19485] = 25'b0000000011110010000000111;
    rom[19486] = 25'b0000000011110010100110010;
    rom[19487] = 25'b0000000011110011001011110;
    rom[19488] = 25'b0000000011110011110001001;
    rom[19489] = 25'b0000000011110100010110101;
    rom[19490] = 25'b0000000011110100111100001;
    rom[19491] = 25'b0000000011110101100001100;
    rom[19492] = 25'b0000000011110110000111000;
    rom[19493] = 25'b0000000011110110101100011;
    rom[19494] = 25'b0000000011110111010001111;
    rom[19495] = 25'b0000000011110111110111010;
    rom[19496] = 25'b0000000011111000011100110;
    rom[19497] = 25'b0000000011111001000010010;
    rom[19498] = 25'b0000000011111001100111101;
    rom[19499] = 25'b0000000011111010001101000;
    rom[19500] = 25'b0000000011111010110010100;
    rom[19501] = 25'b0000000011111011010111111;
    rom[19502] = 25'b0000000011111011111101010;
    rom[19503] = 25'b0000000011111100100010110;
    rom[19504] = 25'b0000000011111101001000001;
    rom[19505] = 25'b0000000011111101101101100;
    rom[19506] = 25'b0000000011111110010011000;
    rom[19507] = 25'b0000000011111110111000011;
    rom[19508] = 25'b0000000011111111011101101;
    rom[19509] = 25'b0000000100000000000011001;
    rom[19510] = 25'b0000000100000000101000100;
    rom[19511] = 25'b0000000100000001001101111;
    rom[19512] = 25'b0000000100000001110011001;
    rom[19513] = 25'b0000000100000010011000100;
    rom[19514] = 25'b0000000100000010111101111;
    rom[19515] = 25'b0000000100000011100011011;
    rom[19516] = 25'b0000000100000100001000101;
    rom[19517] = 25'b0000000100000100101110000;
    rom[19518] = 25'b0000000100000101010011010;
    rom[19519] = 25'b0000000100000101111000101;
    rom[19520] = 25'b0000000100000110011110000;
    rom[19521] = 25'b0000000100000111000011011;
    rom[19522] = 25'b0000000100000111101000101;
    rom[19523] = 25'b0000000100001000001110000;
    rom[19524] = 25'b0000000100001000110011011;
    rom[19525] = 25'b0000000100001001011000101;
    rom[19526] = 25'b0000000100001001111101111;
    rom[19527] = 25'b0000000100001010100011010;
    rom[19528] = 25'b0000000100001011001000100;
    rom[19529] = 25'b0000000100001011101101111;
    rom[19530] = 25'b0000000100001100010011001;
    rom[19531] = 25'b0000000100001100111000011;
    rom[19532] = 25'b0000000100001101011101101;
    rom[19533] = 25'b0000000100001110000010111;
    rom[19534] = 25'b0000000100001110101000001;
    rom[19535] = 25'b0000000100001111001101011;
    rom[19536] = 25'b0000000100001111110010101;
    rom[19537] = 25'b0000000100010000010111111;
    rom[19538] = 25'b0000000100010000111101001;
    rom[19539] = 25'b0000000100010001100010011;
    rom[19540] = 25'b0000000100010010000111101;
    rom[19541] = 25'b0000000100010010101100110;
    rom[19542] = 25'b0000000100010011010010000;
    rom[19543] = 25'b0000000100010011110111010;
    rom[19544] = 25'b0000000100010100011100100;
    rom[19545] = 25'b0000000100010101000001101;
    rom[19546] = 25'b0000000100010101100110111;
    rom[19547] = 25'b0000000100010110001100000;
    rom[19548] = 25'b0000000100010110110001001;
    rom[19549] = 25'b0000000100010111010110011;
    rom[19550] = 25'b0000000100010111111011100;
    rom[19551] = 25'b0000000100011000100000101;
    rom[19552] = 25'b0000000100011001000101111;
    rom[19553] = 25'b0000000100011001101011000;
    rom[19554] = 25'b0000000100011010010000001;
    rom[19555] = 25'b0000000100011010110101010;
    rom[19556] = 25'b0000000100011011011010011;
    rom[19557] = 25'b0000000100011011111111100;
    rom[19558] = 25'b0000000100011100100100101;
    rom[19559] = 25'b0000000100011101001001110;
    rom[19560] = 25'b0000000100011101101110110;
    rom[19561] = 25'b0000000100011110010011111;
    rom[19562] = 25'b0000000100011110111001000;
    rom[19563] = 25'b0000000100011111011110000;
    rom[19564] = 25'b0000000100100000000011001;
    rom[19565] = 25'b0000000100100000101000001;
    rom[19566] = 25'b0000000100100001001101010;
    rom[19567] = 25'b0000000100100001110010011;
    rom[19568] = 25'b0000000100100010010111010;
    rom[19569] = 25'b0000000100100010111100011;
    rom[19570] = 25'b0000000100100011100001011;
    rom[19571] = 25'b0000000100100100000110011;
    rom[19572] = 25'b0000000100100100101011011;
    rom[19573] = 25'b0000000100100101010000011;
    rom[19574] = 25'b0000000100100101110101011;
    rom[19575] = 25'b0000000100100110011010011;
    rom[19576] = 25'b0000000100100110111111011;
    rom[19577] = 25'b0000000100100111100100011;
    rom[19578] = 25'b0000000100101000001001010;
    rom[19579] = 25'b0000000100101000101110010;
    rom[19580] = 25'b0000000100101001010011001;
    rom[19581] = 25'b0000000100101001111000001;
    rom[19582] = 25'b0000000100101010011101000;
    rom[19583] = 25'b0000000100101011000001111;
    rom[19584] = 25'b0000000100101011100110111;
    rom[19585] = 25'b0000000100101100001011110;
    rom[19586] = 25'b0000000100101100110000101;
    rom[19587] = 25'b0000000100101101010101101;
    rom[19588] = 25'b0000000100101101111010100;
    rom[19589] = 25'b0000000100101110011111011;
    rom[19590] = 25'b0000000100101111000100001;
    rom[19591] = 25'b0000000100101111101001000;
    rom[19592] = 25'b0000000100110000001101111;
    rom[19593] = 25'b0000000100110000110010110;
    rom[19594] = 25'b0000000100110001010111100;
    rom[19595] = 25'b0000000100110001111100010;
    rom[19596] = 25'b0000000100110010100001010;
    rom[19597] = 25'b0000000100110011000110000;
    rom[19598] = 25'b0000000100110011101010110;
    rom[19599] = 25'b0000000100110100001111100;
    rom[19600] = 25'b0000000100110100110100010;
    rom[19601] = 25'b0000000100110101011001001;
    rom[19602] = 25'b0000000100110101111101110;
    rom[19603] = 25'b0000000100110110100010101;
    rom[19604] = 25'b0000000100110111000111010;
    rom[19605] = 25'b0000000100110111101100000;
    rom[19606] = 25'b0000000100111000010000110;
    rom[19607] = 25'b0000000100111000110101100;
    rom[19608] = 25'b0000000100111001011010001;
    rom[19609] = 25'b0000000100111001111110110;
    rom[19610] = 25'b0000000100111010100011100;
    rom[19611] = 25'b0000000100111011001000001;
    rom[19612] = 25'b0000000100111011101100110;
    rom[19613] = 25'b0000000100111100010001100;
    rom[19614] = 25'b0000000100111100110110001;
    rom[19615] = 25'b0000000100111101011010110;
    rom[19616] = 25'b0000000100111101111111010;
    rom[19617] = 25'b0000000100111110100011111;
    rom[19618] = 25'b0000000100111111001000100;
    rom[19619] = 25'b0000000100111111101101001;
    rom[19620] = 25'b0000000101000000010001101;
    rom[19621] = 25'b0000000101000000110110010;
    rom[19622] = 25'b0000000101000001011010110;
    rom[19623] = 25'b0000000101000001111111011;
    rom[19624] = 25'b0000000101000010100011111;
    rom[19625] = 25'b0000000101000011001000011;
    rom[19626] = 25'b0000000101000011101100111;
    rom[19627] = 25'b0000000101000100010001011;
    rom[19628] = 25'b0000000101000100110110000;
    rom[19629] = 25'b0000000101000101011010011;
    rom[19630] = 25'b0000000101000101111110111;
    rom[19631] = 25'b0000000101000110100011010;
    rom[19632] = 25'b0000000101000111000111110;
    rom[19633] = 25'b0000000101000111101100001;
    rom[19634] = 25'b0000000101001000010000101;
    rom[19635] = 25'b0000000101001000110101000;
    rom[19636] = 25'b0000000101001001011001011;
    rom[19637] = 25'b0000000101001001111101111;
    rom[19638] = 25'b0000000101001010100010001;
    rom[19639] = 25'b0000000101001011000110101;
    rom[19640] = 25'b0000000101001011101010111;
    rom[19641] = 25'b0000000101001100001111010;
    rom[19642] = 25'b0000000101001100110011100;
    rom[19643] = 25'b0000000101001101010111111;
    rom[19644] = 25'b0000000101001101111100010;
    rom[19645] = 25'b0000000101001110100000100;
    rom[19646] = 25'b0000000101001111000100110;
    rom[19647] = 25'b0000000101001111101001001;
    rom[19648] = 25'b0000000101010000001101011;
    rom[19649] = 25'b0000000101010000110001101;
    rom[19650] = 25'b0000000101010001010101110;
    rom[19651] = 25'b0000000101010001111010000;
    rom[19652] = 25'b0000000101010010011110010;
    rom[19653] = 25'b0000000101010011000010100;
    rom[19654] = 25'b0000000101010011100110101;
    rom[19655] = 25'b0000000101010100001010111;
    rom[19656] = 25'b0000000101010100101111000;
    rom[19657] = 25'b0000000101010101010011001;
    rom[19658] = 25'b0000000101010101110111010;
    rom[19659] = 25'b0000000101010110011011100;
    rom[19660] = 25'b0000000101010110111111101;
    rom[19661] = 25'b0000000101010111100011101;
    rom[19662] = 25'b0000000101011000000111110;
    rom[19663] = 25'b0000000101011000101011111;
    rom[19664] = 25'b0000000101011001001111111;
    rom[19665] = 25'b0000000101011001110011111;
    rom[19666] = 25'b0000000101011010011000000;
    rom[19667] = 25'b0000000101011010111100000;
    rom[19668] = 25'b0000000101011011100000000;
    rom[19669] = 25'b0000000101011100000100000;
    rom[19670] = 25'b0000000101011100101000000;
    rom[19671] = 25'b0000000101011101001011111;
    rom[19672] = 25'b0000000101011101101111111;
    rom[19673] = 25'b0000000101011110010011111;
    rom[19674] = 25'b0000000101011110110111110;
    rom[19675] = 25'b0000000101011111011011110;
    rom[19676] = 25'b0000000101011111111111101;
    rom[19677] = 25'b0000000101100000100011100;
    rom[19678] = 25'b0000000101100001000111011;
    rom[19679] = 25'b0000000101100001101011010;
    rom[19680] = 25'b0000000101100010001111001;
    rom[19681] = 25'b0000000101100010110011000;
    rom[19682] = 25'b0000000101100011010110110;
    rom[19683] = 25'b0000000101100011111010101;
    rom[19684] = 25'b0000000101100100011110011;
    rom[19685] = 25'b0000000101100101000010001;
    rom[19686] = 25'b0000000101100101100101111;
    rom[19687] = 25'b0000000101100110001001110;
    rom[19688] = 25'b0000000101100110101101100;
    rom[19689] = 25'b0000000101100111010001001;
    rom[19690] = 25'b0000000101100111110100111;
    rom[19691] = 25'b0000000101101000011000101;
    rom[19692] = 25'b0000000101101000111100010;
    rom[19693] = 25'b0000000101101001011111111;
    rom[19694] = 25'b0000000101101010000011101;
    rom[19695] = 25'b0000000101101010100111001;
    rom[19696] = 25'b0000000101101011001010111;
    rom[19697] = 25'b0000000101101011101110011;
    rom[19698] = 25'b0000000101101100010010000;
    rom[19699] = 25'b0000000101101100110101101;
    rom[19700] = 25'b0000000101101101011001001;
    rom[19701] = 25'b0000000101101101111100110;
    rom[19702] = 25'b0000000101101110100000010;
    rom[19703] = 25'b0000000101101111000011110;
    rom[19704] = 25'b0000000101101111100111010;
    rom[19705] = 25'b0000000101110000001010110;
    rom[19706] = 25'b0000000101110000101110010;
    rom[19707] = 25'b0000000101110001010001101;
    rom[19708] = 25'b0000000101110001110101001;
    rom[19709] = 25'b0000000101110010011000100;
    rom[19710] = 25'b0000000101110010111100000;
    rom[19711] = 25'b0000000101110011011111011;
    rom[19712] = 25'b0000000101110100000010110;
    rom[19713] = 25'b0000000101110100100110001;
    rom[19714] = 25'b0000000101110101001001100;
    rom[19715] = 25'b0000000101110101101100111;
    rom[19716] = 25'b0000000101110110010000001;
    rom[19717] = 25'b0000000101110110110011011;
    rom[19718] = 25'b0000000101110111010110110;
    rom[19719] = 25'b0000000101110111111010000;
    rom[19720] = 25'b0000000101111000011101010;
    rom[19721] = 25'b0000000101111001000000100;
    rom[19722] = 25'b0000000101111001100011110;
    rom[19723] = 25'b0000000101111010000111000;
    rom[19724] = 25'b0000000101111010101010001;
    rom[19725] = 25'b0000000101111011001101010;
    rom[19726] = 25'b0000000101111011110000100;
    rom[19727] = 25'b0000000101111100010011101;
    rom[19728] = 25'b0000000101111100110110110;
    rom[19729] = 25'b0000000101111101011001110;
    rom[19730] = 25'b0000000101111101111100111;
    rom[19731] = 25'b0000000101111110100000000;
    rom[19732] = 25'b0000000101111111000011000;
    rom[19733] = 25'b0000000101111111100110001;
    rom[19734] = 25'b0000000110000000001001001;
    rom[19735] = 25'b0000000110000000101100001;
    rom[19736] = 25'b0000000110000001001111001;
    rom[19737] = 25'b0000000110000001110010001;
    rom[19738] = 25'b0000000110000010010101001;
    rom[19739] = 25'b0000000110000010111000000;
    rom[19740] = 25'b0000000110000011011011000;
    rom[19741] = 25'b0000000110000011111101111;
    rom[19742] = 25'b0000000110000100100000110;
    rom[19743] = 25'b0000000110000101000011101;
    rom[19744] = 25'b0000000110000101100110100;
    rom[19745] = 25'b0000000110000110001001010;
    rom[19746] = 25'b0000000110000110101100001;
    rom[19747] = 25'b0000000110000111001110111;
    rom[19748] = 25'b0000000110000111110001110;
    rom[19749] = 25'b0000000110001000010100100;
    rom[19750] = 25'b0000000110001000110111001;
    rom[19751] = 25'b0000000110001001011001111;
    rom[19752] = 25'b0000000110001001111100101;
    rom[19753] = 25'b0000000110001010011111010;
    rom[19754] = 25'b0000000110001011000010000;
    rom[19755] = 25'b0000000110001011100100110;
    rom[19756] = 25'b0000000110001100000111011;
    rom[19757] = 25'b0000000110001100101010000;
    rom[19758] = 25'b0000000110001101001100100;
    rom[19759] = 25'b0000000110001101101111001;
    rom[19760] = 25'b0000000110001110010001110;
    rom[19761] = 25'b0000000110001110110100010;
    rom[19762] = 25'b0000000110001111010110111;
    rom[19763] = 25'b0000000110001111111001010;
    rom[19764] = 25'b0000000110010000011011111;
    rom[19765] = 25'b0000000110010000111110011;
    rom[19766] = 25'b0000000110010001100000110;
    rom[19767] = 25'b0000000110010010000011001;
    rom[19768] = 25'b0000000110010010100101101;
    rom[19769] = 25'b0000000110010011001000000;
    rom[19770] = 25'b0000000110010011101010011;
    rom[19771] = 25'b0000000110010100001100110;
    rom[19772] = 25'b0000000110010100101111001;
    rom[19773] = 25'b0000000110010101010001011;
    rom[19774] = 25'b0000000110010101110011110;
    rom[19775] = 25'b0000000110010110010110001;
    rom[19776] = 25'b0000000110010110111000010;
    rom[19777] = 25'b0000000110010111011010100;
    rom[19778] = 25'b0000000110010111111100110;
    rom[19779] = 25'b0000000110011000011111000;
    rom[19780] = 25'b0000000110011001000001001;
    rom[19781] = 25'b0000000110011001100011011;
    rom[19782] = 25'b0000000110011010000101100;
    rom[19783] = 25'b0000000110011010100111101;
    rom[19784] = 25'b0000000110011011001001110;
    rom[19785] = 25'b0000000110011011101011111;
    rom[19786] = 25'b0000000110011100001110000;
    rom[19787] = 25'b0000000110011100110000000;
    rom[19788] = 25'b0000000110011101010010000;
    rom[19789] = 25'b0000000110011101110100000;
    rom[19790] = 25'b0000000110011110010110000;
    rom[19791] = 25'b0000000110011110111000000;
    rom[19792] = 25'b0000000110011111011001111;
    rom[19793] = 25'b0000000110011111111011111;
    rom[19794] = 25'b0000000110100000011101110;
    rom[19795] = 25'b0000000110100000111111110;
    rom[19796] = 25'b0000000110100001100001101;
    rom[19797] = 25'b0000000110100010000011011;
    rom[19798] = 25'b0000000110100010100101010;
    rom[19799] = 25'b0000000110100011000111001;
    rom[19800] = 25'b0000000110100011101000111;
    rom[19801] = 25'b0000000110100100001010101;
    rom[19802] = 25'b0000000110100100101100011;
    rom[19803] = 25'b0000000110100101001110001;
    rom[19804] = 25'b0000000110100101101111111;
    rom[19805] = 25'b0000000110100110010001100;
    rom[19806] = 25'b0000000110100110110011010;
    rom[19807] = 25'b0000000110100111010100111;
    rom[19808] = 25'b0000000110100111110110100;
    rom[19809] = 25'b0000000110101000011000000;
    rom[19810] = 25'b0000000110101000111001101;
    rom[19811] = 25'b0000000110101001011011010;
    rom[19812] = 25'b0000000110101001111100110;
    rom[19813] = 25'b0000000110101010011110010;
    rom[19814] = 25'b0000000110101010111111110;
    rom[19815] = 25'b0000000110101011100001010;
    rom[19816] = 25'b0000000110101100000010110;
    rom[19817] = 25'b0000000110101100100100001;
    rom[19818] = 25'b0000000110101101000101100;
    rom[19819] = 25'b0000000110101101100111000;
    rom[19820] = 25'b0000000110101110001000010;
    rom[19821] = 25'b0000000110101110101001101;
    rom[19822] = 25'b0000000110101111001011000;
    rom[19823] = 25'b0000000110101111101100010;
    rom[19824] = 25'b0000000110110000001101100;
    rom[19825] = 25'b0000000110110000101110110;
    rom[19826] = 25'b0000000110110001010000000;
    rom[19827] = 25'b0000000110110001110001010;
    rom[19828] = 25'b0000000110110010010010011;
    rom[19829] = 25'b0000000110110010110011101;
    rom[19830] = 25'b0000000110110011010100111;
    rom[19831] = 25'b0000000110110011110101111;
    rom[19832] = 25'b0000000110110100010111000;
    rom[19833] = 25'b0000000110110100111000001;
    rom[19834] = 25'b0000000110110101011001001;
    rom[19835] = 25'b0000000110110101111010010;
    rom[19836] = 25'b0000000110110110011011010;
    rom[19837] = 25'b0000000110110110111100010;
    rom[19838] = 25'b0000000110110111011101010;
    rom[19839] = 25'b0000000110110111111110001;
    rom[19840] = 25'b0000000110111000011111000;
    rom[19841] = 25'b0000000110111000111111111;
    rom[19842] = 25'b0000000110111001100000110;
    rom[19843] = 25'b0000000110111010000001101;
    rom[19844] = 25'b0000000110111010100010100;
    rom[19845] = 25'b0000000110111011000011011;
    rom[19846] = 25'b0000000110111011100100001;
    rom[19847] = 25'b0000000110111100000100111;
    rom[19848] = 25'b0000000110111100100101100;
    rom[19849] = 25'b0000000110111101000110011;
    rom[19850] = 25'b0000000110111101100111000;
    rom[19851] = 25'b0000000110111110000111110;
    rom[19852] = 25'b0000000110111110101000010;
    rom[19853] = 25'b0000000110111111001001000;
    rom[19854] = 25'b0000000110111111101001101;
    rom[19855] = 25'b0000000111000000001010001;
    rom[19856] = 25'b0000000111000000101010101;
    rom[19857] = 25'b0000000111000001001011001;
    rom[19858] = 25'b0000000111000001101011101;
    rom[19859] = 25'b0000000111000010001100001;
    rom[19860] = 25'b0000000111000010101100101;
    rom[19861] = 25'b0000000111000011001101001;
    rom[19862] = 25'b0000000111000011101101100;
    rom[19863] = 25'b0000000111000100001101111;
    rom[19864] = 25'b0000000111000100101110010;
    rom[19865] = 25'b0000000111000101001110100;
    rom[19866] = 25'b0000000111000101101110111;
    rom[19867] = 25'b0000000111000110001111001;
    rom[19868] = 25'b0000000111000110101111100;
    rom[19869] = 25'b0000000111000111001111101;
    rom[19870] = 25'b0000000111000111101111111;
    rom[19871] = 25'b0000000111001000010000000;
    rom[19872] = 25'b0000000111001000110000010;
    rom[19873] = 25'b0000000111001001010000011;
    rom[19874] = 25'b0000000111001001110000100;
    rom[19875] = 25'b0000000111001010010000100;
    rom[19876] = 25'b0000000111001010110000101;
    rom[19877] = 25'b0000000111001011010000101;
    rom[19878] = 25'b0000000111001011110000110;
    rom[19879] = 25'b0000000111001100010000101;
    rom[19880] = 25'b0000000111001100110000101;
    rom[19881] = 25'b0000000111001101010000100;
    rom[19882] = 25'b0000000111001101110000100;
    rom[19883] = 25'b0000000111001110010000011;
    rom[19884] = 25'b0000000111001110110000010;
    rom[19885] = 25'b0000000111001111010000001;
    rom[19886] = 25'b0000000111001111101111111;
    rom[19887] = 25'b0000000111010000001111101;
    rom[19888] = 25'b0000000111010000101111011;
    rom[19889] = 25'b0000000111010001001111001;
    rom[19890] = 25'b0000000111010001101110111;
    rom[19891] = 25'b0000000111010010001110101;
    rom[19892] = 25'b0000000111010010101110010;
    rom[19893] = 25'b0000000111010011001101110;
    rom[19894] = 25'b0000000111010011101101100;
    rom[19895] = 25'b0000000111010100001101000;
    rom[19896] = 25'b0000000111010100101100101;
    rom[19897] = 25'b0000000111010101001100001;
    rom[19898] = 25'b0000000111010101101011101;
    rom[19899] = 25'b0000000111010110001011001;
    rom[19900] = 25'b0000000111010110101010101;
    rom[19901] = 25'b0000000111010111001010000;
    rom[19902] = 25'b0000000111010111101001011;
    rom[19903] = 25'b0000000111011000001000110;
    rom[19904] = 25'b0000000111011000101000001;
    rom[19905] = 25'b0000000111011001000111011;
    rom[19906] = 25'b0000000111011001100110101;
    rom[19907] = 25'b0000000111011010000110000;
    rom[19908] = 25'b0000000111011010100101010;
    rom[19909] = 25'b0000000111011011000100011;
    rom[19910] = 25'b0000000111011011100011101;
    rom[19911] = 25'b0000000111011100000010110;
    rom[19912] = 25'b0000000111011100100001111;
    rom[19913] = 25'b0000000111011101000001000;
    rom[19914] = 25'b0000000111011101100000001;
    rom[19915] = 25'b0000000111011101111111001;
    rom[19916] = 25'b0000000111011110011110001;
    rom[19917] = 25'b0000000111011110111101001;
    rom[19918] = 25'b0000000111011111011100001;
    rom[19919] = 25'b0000000111011111111011000;
    rom[19920] = 25'b0000000111100000011001111;
    rom[19921] = 25'b0000000111100000111000111;
    rom[19922] = 25'b0000000111100001010111101;
    rom[19923] = 25'b0000000111100001110110100;
    rom[19924] = 25'b0000000111100010010101010;
    rom[19925] = 25'b0000000111100010110100001;
    rom[19926] = 25'b0000000111100011010010111;
    rom[19927] = 25'b0000000111100011110001101;
    rom[19928] = 25'b0000000111100100010000010;
    rom[19929] = 25'b0000000111100100101110111;
    rom[19930] = 25'b0000000111100101001101100;
    rom[19931] = 25'b0000000111100101101100001;
    rom[19932] = 25'b0000000111100110001010110;
    rom[19933] = 25'b0000000111100110101001011;
    rom[19934] = 25'b0000000111100111000111110;
    rom[19935] = 25'b0000000111100111100110011;
    rom[19936] = 25'b0000000111101000000100110;
    rom[19937] = 25'b0000000111101000100011010;
    rom[19938] = 25'b0000000111101001000001101;
    rom[19939] = 25'b0000000111101001100000000;
    rom[19940] = 25'b0000000111101001111110011;
    rom[19941] = 25'b0000000111101010011100110;
    rom[19942] = 25'b0000000111101010111011000;
    rom[19943] = 25'b0000000111101011011001010;
    rom[19944] = 25'b0000000111101011110111100;
    rom[19945] = 25'b0000000111101100010101110;
    rom[19946] = 25'b0000000111101100110011111;
    rom[19947] = 25'b0000000111101101010010001;
    rom[19948] = 25'b0000000111101101110000010;
    rom[19949] = 25'b0000000111101110001110010;
    rom[19950] = 25'b0000000111101110101100011;
    rom[19951] = 25'b0000000111101111001010011;
    rom[19952] = 25'b0000000111101111101000011;
    rom[19953] = 25'b0000000111110000000110011;
    rom[19954] = 25'b0000000111110000100100010;
    rom[19955] = 25'b0000000111110001000010010;
    rom[19956] = 25'b0000000111110001100000001;
    rom[19957] = 25'b0000000111110001111110000;
    rom[19958] = 25'b0000000111110010011011111;
    rom[19959] = 25'b0000000111110010111001101;
    rom[19960] = 25'b0000000111110011010111011;
    rom[19961] = 25'b0000000111110011110101010;
    rom[19962] = 25'b0000000111110100010010111;
    rom[19963] = 25'b0000000111110100110000101;
    rom[19964] = 25'b0000000111110101001110010;
    rom[19965] = 25'b0000000111110101101011110;
    rom[19966] = 25'b0000000111110110001001011;
    rom[19967] = 25'b0000000111110110100111000;
    rom[19968] = 25'b0000000111110111000100100;
    rom[19969] = 25'b0000000111110111100010000;
    rom[19970] = 25'b0000000111110111111111100;
    rom[19971] = 25'b0000000111111000011101000;
    rom[19972] = 25'b0000000111111000111010011;
    rom[19973] = 25'b0000000111111001010111110;
    rom[19974] = 25'b0000000111111001110101001;
    rom[19975] = 25'b0000000111111010010010011;
    rom[19976] = 25'b0000000111111010101111110;
    rom[19977] = 25'b0000000111111011001101000;
    rom[19978] = 25'b0000000111111011101010010;
    rom[19979] = 25'b0000000111111100000111100;
    rom[19980] = 25'b0000000111111100100100101;
    rom[19981] = 25'b0000000111111101000001110;
    rom[19982] = 25'b0000000111111101011110111;
    rom[19983] = 25'b0000000111111101111011111;
    rom[19984] = 25'b0000000111111110011001000;
    rom[19985] = 25'b0000000111111110110110000;
    rom[19986] = 25'b0000000111111111010010111;
    rom[19987] = 25'b0000000111111111101111111;
    rom[19988] = 25'b0000001000000000001100111;
    rom[19989] = 25'b0000001000000000101001110;
    rom[19990] = 25'b0000001000000001000110100;
    rom[19991] = 25'b0000001000000001100011011;
    rom[19992] = 25'b0000001000000010000000010;
    rom[19993] = 25'b0000001000000010011101000;
    rom[19994] = 25'b0000001000000010111001110;
    rom[19995] = 25'b0000001000000011010110100;
    rom[19996] = 25'b0000001000000011110011001;
    rom[19997] = 25'b0000001000000100001111110;
    rom[19998] = 25'b0000001000000100101100011;
    rom[19999] = 25'b0000001000000101001001000;
    rom[20000] = 25'b0000001000000101100101011;
    rom[20001] = 25'b0000001000000110000010000;
    rom[20002] = 25'b0000001000000110011110100;
    rom[20003] = 25'b0000001000000110111010111;
    rom[20004] = 25'b0000001000000111010111011;
    rom[20005] = 25'b0000001000000111110011110;
    rom[20006] = 25'b0000001000001000010000000;
    rom[20007] = 25'b0000001000001000101100011;
    rom[20008] = 25'b0000001000001001001000101;
    rom[20009] = 25'b0000001000001001100101000;
    rom[20010] = 25'b0000001000001010000001001;
    rom[20011] = 25'b0000001000001010011101011;
    rom[20012] = 25'b0000001000001010111001100;
    rom[20013] = 25'b0000001000001011010101101;
    rom[20014] = 25'b0000001000001011110001101;
    rom[20015] = 25'b0000001000001100001101110;
    rom[20016] = 25'b0000001000001100101001110;
    rom[20017] = 25'b0000001000001101000101111;
    rom[20018] = 25'b0000001000001101100001110;
    rom[20019] = 25'b0000001000001101111101101;
    rom[20020] = 25'b0000001000001110011001101;
    rom[20021] = 25'b0000001000001110110101011;
    rom[20022] = 25'b0000001000001111010001011;
    rom[20023] = 25'b0000001000001111101101001;
    rom[20024] = 25'b0000001000010000001000110;
    rom[20025] = 25'b0000001000010000100100100;
    rom[20026] = 25'b0000001000010001000000010;
    rom[20027] = 25'b0000001000010001011011111;
    rom[20028] = 25'b0000001000010001110111101;
    rom[20029] = 25'b0000001000010010010011010;
    rom[20030] = 25'b0000001000010010101110110;
    rom[20031] = 25'b0000001000010011001010010;
    rom[20032] = 25'b0000001000010011100101110;
    rom[20033] = 25'b0000001000010100000001010;
    rom[20034] = 25'b0000001000010100011100101;
    rom[20035] = 25'b0000001000010100111000000;
    rom[20036] = 25'b0000001000010101010011011;
    rom[20037] = 25'b0000001000010101101110110;
    rom[20038] = 25'b0000001000010110001010000;
    rom[20039] = 25'b0000001000010110100101010;
    rom[20040] = 25'b0000001000010111000000101;
    rom[20041] = 25'b0000001000010111011011110;
    rom[20042] = 25'b0000001000010111110110111;
    rom[20043] = 25'b0000001000011000010010000;
    rom[20044] = 25'b0000001000011000101101001;
    rom[20045] = 25'b0000001000011001001000001;
    rom[20046] = 25'b0000001000011001100011001;
    rom[20047] = 25'b0000001000011001111110001;
    rom[20048] = 25'b0000001000011010011001001;
    rom[20049] = 25'b0000001000011010110100000;
    rom[20050] = 25'b0000001000011011001110111;
    rom[20051] = 25'b0000001000011011101001111;
    rom[20052] = 25'b0000001000011100000100101;
    rom[20053] = 25'b0000001000011100011111011;
    rom[20054] = 25'b0000001000011100111010001;
    rom[20055] = 25'b0000001000011101010100111;
    rom[20056] = 25'b0000001000011101101111100;
    rom[20057] = 25'b0000001000011110001010001;
    rom[20058] = 25'b0000001000011110100100110;
    rom[20059] = 25'b0000001000011110111111010;
    rom[20060] = 25'b0000001000011111011001111;
    rom[20061] = 25'b0000001000011111110100011;
    rom[20062] = 25'b0000001000100000001110111;
    rom[20063] = 25'b0000001000100000101001010;
    rom[20064] = 25'b0000001000100001000011101;
    rom[20065] = 25'b0000001000100001011110000;
    rom[20066] = 25'b0000001000100001111000011;
    rom[20067] = 25'b0000001000100010010010101;
    rom[20068] = 25'b0000001000100010101100111;
    rom[20069] = 25'b0000001000100011000111001;
    rom[20070] = 25'b0000001000100011100001010;
    rom[20071] = 25'b0000001000100011111011011;
    rom[20072] = 25'b0000001000100100010101101;
    rom[20073] = 25'b0000001000100100101111101;
    rom[20074] = 25'b0000001000100101001001101;
    rom[20075] = 25'b0000001000100101100011101;
    rom[20076] = 25'b0000001000100101111101110;
    rom[20077] = 25'b0000001000100110010111100;
    rom[20078] = 25'b0000001000100110110001011;
    rom[20079] = 25'b0000001000100111001011010;
    rom[20080] = 25'b0000001000100111100101001;
    rom[20081] = 25'b0000001000100111111111000;
    rom[20082] = 25'b0000001000101000011000110;
    rom[20083] = 25'b0000001000101000110010011;
    rom[20084] = 25'b0000001000101001001100001;
    rom[20085] = 25'b0000001000101001100101110;
    rom[20086] = 25'b0000001000101001111111011;
    rom[20087] = 25'b0000001000101010011000111;
    rom[20088] = 25'b0000001000101010110010011;
    rom[20089] = 25'b0000001000101011001011111;
    rom[20090] = 25'b0000001000101011100101011;
    rom[20091] = 25'b0000001000101011111110111;
    rom[20092] = 25'b0000001000101100011000010;
    rom[20093] = 25'b0000001000101100110001100;
    rom[20094] = 25'b0000001000101101001010111;
    rom[20095] = 25'b0000001000101101100100001;
    rom[20096] = 25'b0000001000101101111101011;
    rom[20097] = 25'b0000001000101110010110101;
    rom[20098] = 25'b0000001000101110101111110;
    rom[20099] = 25'b0000001000101111001000111;
    rom[20100] = 25'b0000001000101111100001111;
    rom[20101] = 25'b0000001000101111111011000;
    rom[20102] = 25'b0000001000110000010100000;
    rom[20103] = 25'b0000001000110000101101000;
    rom[20104] = 25'b0000001000110001000110000;
    rom[20105] = 25'b0000001000110001011110111;
    rom[20106] = 25'b0000001000110001110111110;
    rom[20107] = 25'b0000001000110010010000101;
    rom[20108] = 25'b0000001000110010101001011;
    rom[20109] = 25'b0000001000110011000010001;
    rom[20110] = 25'b0000001000110011011010111;
    rom[20111] = 25'b0000001000110011110011100;
    rom[20112] = 25'b0000001000110100001100001;
    rom[20113] = 25'b0000001000110100100100101;
    rom[20114] = 25'b0000001000110100111101010;
    rom[20115] = 25'b0000001000110101010101110;
    rom[20116] = 25'b0000001000110101101110010;
    rom[20117] = 25'b0000001000110110000110110;
    rom[20118] = 25'b0000001000110110011111010;
    rom[20119] = 25'b0000001000110110110111101;
    rom[20120] = 25'b0000001000110111001111111;
    rom[20121] = 25'b0000001000110111101000001;
    rom[20122] = 25'b0000001000111000000000011;
    rom[20123] = 25'b0000001000111000011000101;
    rom[20124] = 25'b0000001000111000110000110;
    rom[20125] = 25'b0000001000111001001001000;
    rom[20126] = 25'b0000001000111001100001001;
    rom[20127] = 25'b0000001000111001111001001;
    rom[20128] = 25'b0000001000111010010001001;
    rom[20129] = 25'b0000001000111010101001001;
    rom[20130] = 25'b0000001000111011000001001;
    rom[20131] = 25'b0000001000111011011001000;
    rom[20132] = 25'b0000001000111011110000111;
    rom[20133] = 25'b0000001000111100001000110;
    rom[20134] = 25'b0000001000111100100000100;
    rom[20135] = 25'b0000001000111100111000010;
    rom[20136] = 25'b0000001000111101010000000;
    rom[20137] = 25'b0000001000111101100111101;
    rom[20138] = 25'b0000001000111101111111010;
    rom[20139] = 25'b0000001000111110010110111;
    rom[20140] = 25'b0000001000111110101110100;
    rom[20141] = 25'b0000001000111111000110000;
    rom[20142] = 25'b0000001000111111011101100;
    rom[20143] = 25'b0000001000111111110100111;
    rom[20144] = 25'b0000001001000000001100011;
    rom[20145] = 25'b0000001001000000100011101;
    rom[20146] = 25'b0000001001000000111011000;
    rom[20147] = 25'b0000001001000001010010010;
    rom[20148] = 25'b0000001001000001101001100;
    rom[20149] = 25'b0000001001000010000000101;
    rom[20150] = 25'b0000001001000010010111111;
    rom[20151] = 25'b0000001001000010101111000;
    rom[20152] = 25'b0000001001000011000110001;
    rom[20153] = 25'b0000001001000011011101001;
    rom[20154] = 25'b0000001001000011110100001;
    rom[20155] = 25'b0000001001000100001011001;
    rom[20156] = 25'b0000001001000100100010000;
    rom[20157] = 25'b0000001001000100111000111;
    rom[20158] = 25'b0000001001000101001111110;
    rom[20159] = 25'b0000001001000101100110100;
    rom[20160] = 25'b0000001001000101111101010;
    rom[20161] = 25'b0000001001000110010100000;
    rom[20162] = 25'b0000001001000110101010101;
    rom[20163] = 25'b0000001001000111000001011;
    rom[20164] = 25'b0000001001000111011000000;
    rom[20165] = 25'b0000001001000111101110100;
    rom[20166] = 25'b0000001001001000000101001;
    rom[20167] = 25'b0000001001001000011011100;
    rom[20168] = 25'b0000001001001000110001111;
    rom[20169] = 25'b0000001001001001001000011;
    rom[20170] = 25'b0000001001001001011110110;
    rom[20171] = 25'b0000001001001001110101000;
    rom[20172] = 25'b0000001001001010001011010;
    rom[20173] = 25'b0000001001001010100001100;
    rom[20174] = 25'b0000001001001010110111110;
    rom[20175] = 25'b0000001001001011001101111;
    rom[20176] = 25'b0000001001001011100100000;
    rom[20177] = 25'b0000001001001011111010000;
    rom[20178] = 25'b0000001001001100010000001;
    rom[20179] = 25'b0000001001001100100110001;
    rom[20180] = 25'b0000001001001100111100000;
    rom[20181] = 25'b0000001001001101010001111;
    rom[20182] = 25'b0000001001001101100111110;
    rom[20183] = 25'b0000001001001101111101101;
    rom[20184] = 25'b0000001001001110010011011;
    rom[20185] = 25'b0000001001001110101001001;
    rom[20186] = 25'b0000001001001110111110110;
    rom[20187] = 25'b0000001001001111010100100;
    rom[20188] = 25'b0000001001001111101010001;
    rom[20189] = 25'b0000001001001111111111110;
    rom[20190] = 25'b0000001001010000010101001;
    rom[20191] = 25'b0000001001010000101010101;
    rom[20192] = 25'b0000001001010001000000001;
    rom[20193] = 25'b0000001001010001010101100;
    rom[20194] = 25'b0000001001010001101010111;
    rom[20195] = 25'b0000001001010010000000010;
    rom[20196] = 25'b0000001001010010010101100;
    rom[20197] = 25'b0000001001010010101010110;
    rom[20198] = 25'b0000001001010010111111111;
    rom[20199] = 25'b0000001001010011010101001;
    rom[20200] = 25'b0000001001010011101010010;
    rom[20201] = 25'b0000001001010011111111010;
    rom[20202] = 25'b0000001001010100010100010;
    rom[20203] = 25'b0000001001010100101001010;
    rom[20204] = 25'b0000001001010100111110001;
    rom[20205] = 25'b0000001001010101010011001;
    rom[20206] = 25'b0000001001010101100111111;
    rom[20207] = 25'b0000001001010101111100110;
    rom[20208] = 25'b0000001001010110010001100;
    rom[20209] = 25'b0000001001010110100110010;
    rom[20210] = 25'b0000001001010110111010111;
    rom[20211] = 25'b0000001001010111001111100;
    rom[20212] = 25'b0000001001010111100100010;
    rom[20213] = 25'b0000001001010111111000110;
    rom[20214] = 25'b0000001001011000001101010;
    rom[20215] = 25'b0000001001011000100001101;
    rom[20216] = 25'b0000001001011000110110001;
    rom[20217] = 25'b0000001001011001001010100;
    rom[20218] = 25'b0000001001011001011110111;
    rom[20219] = 25'b0000001001011001110011001;
    rom[20220] = 25'b0000001001011010000111011;
    rom[20221] = 25'b0000001001011010011011101;
    rom[20222] = 25'b0000001001011010101111110;
    rom[20223] = 25'b0000001001011011000011111;
    rom[20224] = 25'b0000001001011011010111111;
    rom[20225] = 25'b0000001001011011101100000;
    rom[20226] = 25'b0000001001011100000000000;
    rom[20227] = 25'b0000001001011100010011111;
    rom[20228] = 25'b0000001001011100100111111;
    rom[20229] = 25'b0000001001011100111011101;
    rom[20230] = 25'b0000001001011101001111100;
    rom[20231] = 25'b0000001001011101100011010;
    rom[20232] = 25'b0000001001011101110111000;
    rom[20233] = 25'b0000001001011110001010101;
    rom[20234] = 25'b0000001001011110011110010;
    rom[20235] = 25'b0000001001011110110001111;
    rom[20236] = 25'b0000001001011111000101100;
    rom[20237] = 25'b0000001001011111011001000;
    rom[20238] = 25'b0000001001011111101100100;
    rom[20239] = 25'b0000001001011111111111111;
    rom[20240] = 25'b0000001001100000010011010;
    rom[20241] = 25'b0000001001100000100110100;
    rom[20242] = 25'b0000001001100000111001111;
    rom[20243] = 25'b0000001001100001001101001;
    rom[20244] = 25'b0000001001100001100000011;
    rom[20245] = 25'b0000001001100001110011100;
    rom[20246] = 25'b0000001001100010000110100;
    rom[20247] = 25'b0000001001100010011001101;
    rom[20248] = 25'b0000001001100010101100101;
    rom[20249] = 25'b0000001001100010111111101;
    rom[20250] = 25'b0000001001100011010010100;
    rom[20251] = 25'b0000001001100011100101011;
    rom[20252] = 25'b0000001001100011111000010;
    rom[20253] = 25'b0000001001100100001011000;
    rom[20254] = 25'b0000001001100100011101111;
    rom[20255] = 25'b0000001001100100110000100;
    rom[20256] = 25'b0000001001100101000011001;
    rom[20257] = 25'b0000001001100101010101110;
    rom[20258] = 25'b0000001001100101101000011;
    rom[20259] = 25'b0000001001100101111011000;
    rom[20260] = 25'b0000001001100110001101011;
    rom[20261] = 25'b0000001001100110011111111;
    rom[20262] = 25'b0000001001100110110010010;
    rom[20263] = 25'b0000001001100111000100100;
    rom[20264] = 25'b0000001001100111010110111;
    rom[20265] = 25'b0000001001100111101001001;
    rom[20266] = 25'b0000001001100111111011011;
    rom[20267] = 25'b0000001001101000001101100;
    rom[20268] = 25'b0000001001101000011111101;
    rom[20269] = 25'b0000001001101000110001110;
    rom[20270] = 25'b0000001001101001000011110;
    rom[20271] = 25'b0000001001101001010101101;
    rom[20272] = 25'b0000001001101001100111101;
    rom[20273] = 25'b0000001001101001111001100;
    rom[20274] = 25'b0000001001101010001011011;
    rom[20275] = 25'b0000001001101010011101001;
    rom[20276] = 25'b0000001001101010101110111;
    rom[20277] = 25'b0000001001101011000000101;
    rom[20278] = 25'b0000001001101011010010010;
    rom[20279] = 25'b0000001001101011100011111;
    rom[20280] = 25'b0000001001101011110101011;
    rom[20281] = 25'b0000001001101100000110111;
    rom[20282] = 25'b0000001001101100011000011;
    rom[20283] = 25'b0000001001101100101001111;
    rom[20284] = 25'b0000001001101100111011010;
    rom[20285] = 25'b0000001001101101001100101;
    rom[20286] = 25'b0000001001101101011101111;
    rom[20287] = 25'b0000001001101101101111000;
    rom[20288] = 25'b0000001001101110000000010;
    rom[20289] = 25'b0000001001101110010001011;
    rom[20290] = 25'b0000001001101110100010100;
    rom[20291] = 25'b0000001001101110110011101;
    rom[20292] = 25'b0000001001101111000100101;
    rom[20293] = 25'b0000001001101111010101101;
    rom[20294] = 25'b0000001001101111100110100;
    rom[20295] = 25'b0000001001101111110111010;
    rom[20296] = 25'b0000001001110000001000001;
    rom[20297] = 25'b0000001001110000011000111;
    rom[20298] = 25'b0000001001110000101001101;
    rom[20299] = 25'b0000001001110000111010011;
    rom[20300] = 25'b0000001001110001001011000;
    rom[20301] = 25'b0000001001110001011011100;
    rom[20302] = 25'b0000001001110001101100001;
    rom[20303] = 25'b0000001001110001111100100;
    rom[20304] = 25'b0000001001110010001101000;
    rom[20305] = 25'b0000001001110010011101011;
    rom[20306] = 25'b0000001001110010101101110;
    rom[20307] = 25'b0000001001110010111110000;
    rom[20308] = 25'b0000001001110011001110010;
    rom[20309] = 25'b0000001001110011011110100;
    rom[20310] = 25'b0000001001110011101110101;
    rom[20311] = 25'b0000001001110011111110111;
    rom[20312] = 25'b0000001001110100001110111;
    rom[20313] = 25'b0000001001110100011110111;
    rom[20314] = 25'b0000001001110100101110111;
    rom[20315] = 25'b0000001001110100111110110;
    rom[20316] = 25'b0000001001110101001110101;
    rom[20317] = 25'b0000001001110101011110100;
    rom[20318] = 25'b0000001001110101101110010;
    rom[20319] = 25'b0000001001110101111101111;
    rom[20320] = 25'b0000001001110110001101101;
    rom[20321] = 25'b0000001001110110011101010;
    rom[20322] = 25'b0000001001110110101100111;
    rom[20323] = 25'b0000001001110110111100011;
    rom[20324] = 25'b0000001001110111001011111;
    rom[20325] = 25'b0000001001110111011011010;
    rom[20326] = 25'b0000001001110111101010110;
    rom[20327] = 25'b0000001001110111111010000;
    rom[20328] = 25'b0000001001111000001001011;
    rom[20329] = 25'b0000001001111000011000101;
    rom[20330] = 25'b0000001001111000100111110;
    rom[20331] = 25'b0000001001111000110110111;
    rom[20332] = 25'b0000001001111001000110000;
    rom[20333] = 25'b0000001001111001010101001;
    rom[20334] = 25'b0000001001111001100100001;
    rom[20335] = 25'b0000001001111001110011000;
    rom[20336] = 25'b0000001001111010000010000;
    rom[20337] = 25'b0000001001111010010000111;
    rom[20338] = 25'b0000001001111010011111101;
    rom[20339] = 25'b0000001001111010101110011;
    rom[20340] = 25'b0000001001111010111101001;
    rom[20341] = 25'b0000001001111011001011110;
    rom[20342] = 25'b0000001001111011011010011;
    rom[20343] = 25'b0000001001111011101000111;
    rom[20344] = 25'b0000001001111011110111100;
    rom[20345] = 25'b0000001001111100000110000;
    rom[20346] = 25'b0000001001111100010100011;
    rom[20347] = 25'b0000001001111100100010110;
    rom[20348] = 25'b0000001001111100110001000;
    rom[20349] = 25'b0000001001111100111111010;
    rom[20350] = 25'b0000001001111101001101100;
    rom[20351] = 25'b0000001001111101011011101;
    rom[20352] = 25'b0000001001111101101001110;
    rom[20353] = 25'b0000001001111101110111111;
    rom[20354] = 25'b0000001001111110000101111;
    rom[20355] = 25'b0000001001111110010011111;
    rom[20356] = 25'b0000001001111110100001111;
    rom[20357] = 25'b0000001001111110101111101;
    rom[20358] = 25'b0000001001111110111101100;
    rom[20359] = 25'b0000001001111111001011010;
    rom[20360] = 25'b0000001001111111011001000;
    rom[20361] = 25'b0000001001111111100110101;
    rom[20362] = 25'b0000001001111111110100010;
    rom[20363] = 25'b0000001010000000000001111;
    rom[20364] = 25'b0000001010000000001111011;
    rom[20365] = 25'b0000001010000000011100111;
    rom[20366] = 25'b0000001010000000101010010;
    rom[20367] = 25'b0000001010000000110111110;
    rom[20368] = 25'b0000001010000001000101000;
    rom[20369] = 25'b0000001010000001010010011;
    rom[20370] = 25'b0000001010000001011111100;
    rom[20371] = 25'b0000001010000001101100101;
    rom[20372] = 25'b0000001010000001111001111;
    rom[20373] = 25'b0000001010000010000110111;
    rom[20374] = 25'b0000001010000010010011111;
    rom[20375] = 25'b0000001010000010100000111;
    rom[20376] = 25'b0000001010000010101101111;
    rom[20377] = 25'b0000001010000010111010101;
    rom[20378] = 25'b0000001010000011000111100;
    rom[20379] = 25'b0000001010000011010100010;
    rom[20380] = 25'b0000001010000011100001000;
    rom[20381] = 25'b0000001010000011101101101;
    rom[20382] = 25'b0000001010000011111010010;
    rom[20383] = 25'b0000001010000100000110111;
    rom[20384] = 25'b0000001010000100010011011;
    rom[20385] = 25'b0000001010000100011111111;
    rom[20386] = 25'b0000001010000100101100010;
    rom[20387] = 25'b0000001010000100111000101;
    rom[20388] = 25'b0000001010000101000101000;
    rom[20389] = 25'b0000001010000101010001001;
    rom[20390] = 25'b0000001010000101011101011;
    rom[20391] = 25'b0000001010000101101001100;
    rom[20392] = 25'b0000001010000101110101101;
    rom[20393] = 25'b0000001010000110000001110;
    rom[20394] = 25'b0000001010000110001101110;
    rom[20395] = 25'b0000001010000110011001110;
    rom[20396] = 25'b0000001010000110100101101;
    rom[20397] = 25'b0000001010000110110001100;
    rom[20398] = 25'b0000001010000110111101010;
    rom[20399] = 25'b0000001010000111001001000;
    rom[20400] = 25'b0000001010000111010100110;
    rom[20401] = 25'b0000001010000111100000011;
    rom[20402] = 25'b0000001010000111101011111;
    rom[20403] = 25'b0000001010000111110111100;
    rom[20404] = 25'b0000001010001000000011000;
    rom[20405] = 25'b0000001010001000001110100;
    rom[20406] = 25'b0000001010001000011001111;
    rom[20407] = 25'b0000001010001000100101001;
    rom[20408] = 25'b0000001010001000110000100;
    rom[20409] = 25'b0000001010001000111011101;
    rom[20410] = 25'b0000001010001001000110111;
    rom[20411] = 25'b0000001010001001010010000;
    rom[20412] = 25'b0000001010001001011101001;
    rom[20413] = 25'b0000001010001001101000001;
    rom[20414] = 25'b0000001010001001110011001;
    rom[20415] = 25'b0000001010001001111110001;
    rom[20416] = 25'b0000001010001010001000111;
    rom[20417] = 25'b0000001010001010010011110;
    rom[20418] = 25'b0000001010001010011110100;
    rom[20419] = 25'b0000001010001010101001010;
    rom[20420] = 25'b0000001010001010110011111;
    rom[20421] = 25'b0000001010001010111110100;
    rom[20422] = 25'b0000001010001011001001000;
    rom[20423] = 25'b0000001010001011010011100;
    rom[20424] = 25'b0000001010001011011110000;
    rom[20425] = 25'b0000001010001011101000011;
    rom[20426] = 25'b0000001010001011110010110;
    rom[20427] = 25'b0000001010001011111101001;
    rom[20428] = 25'b0000001010001100000111010;
    rom[20429] = 25'b0000001010001100010001100;
    rom[20430] = 25'b0000001010001100011011101;
    rom[20431] = 25'b0000001010001100100101110;
    rom[20432] = 25'b0000001010001100101111110;
    rom[20433] = 25'b0000001010001100111001101;
    rom[20434] = 25'b0000001010001101000011101;
    rom[20435] = 25'b0000001010001101001101101;
    rom[20436] = 25'b0000001010001101010111011;
    rom[20437] = 25'b0000001010001101100001001;
    rom[20438] = 25'b0000001010001101101010110;
    rom[20439] = 25'b0000001010001101110100100;
    rom[20440] = 25'b0000001010001101111110001;
    rom[20441] = 25'b0000001010001110000111101;
    rom[20442] = 25'b0000001010001110010001001;
    rom[20443] = 25'b0000001010001110011010101;
    rom[20444] = 25'b0000001010001110100100000;
    rom[20445] = 25'b0000001010001110101101011;
    rom[20446] = 25'b0000001010001110110110101;
    rom[20447] = 25'b0000001010001110111111111;
    rom[20448] = 25'b0000001010001111001001001;
    rom[20449] = 25'b0000001010001111010010001;
    rom[20450] = 25'b0000001010001111011011011;
    rom[20451] = 25'b0000001010001111100100010;
    rom[20452] = 25'b0000001010001111101101010;
    rom[20453] = 25'b0000001010001111110110010;
    rom[20454] = 25'b0000001010001111111111001;
    rom[20455] = 25'b0000001010010000000111111;
    rom[20456] = 25'b0000001010010000010000101;
    rom[20457] = 25'b0000001010010000011001011;
    rom[20458] = 25'b0000001010010000100010000;
    rom[20459] = 25'b0000001010010000101010101;
    rom[20460] = 25'b0000001010010000110011001;
    rom[20461] = 25'b0000001010010000111011101;
    rom[20462] = 25'b0000001010010001000100001;
    rom[20463] = 25'b0000001010010001001100011;
    rom[20464] = 25'b0000001010010001010100110;
    rom[20465] = 25'b0000001010010001011101000;
    rom[20466] = 25'b0000001010010001100101010;
    rom[20467] = 25'b0000001010010001101101011;
    rom[20468] = 25'b0000001010010001110101100;
    rom[20469] = 25'b0000001010010001111101101;
    rom[20470] = 25'b0000001010010010000101101;
    rom[20471] = 25'b0000001010010010001101100;
    rom[20472] = 25'b0000001010010010010101100;
    rom[20473] = 25'b0000001010010010011101010;
    rom[20474] = 25'b0000001010010010100101000;
    rom[20475] = 25'b0000001010010010101100110;
    rom[20476] = 25'b0000001010010010110100100;
    rom[20477] = 25'b0000001010010010111100001;
    rom[20478] = 25'b0000001010010011000011101;
    rom[20479] = 25'b0000001010010011001011001;
    rom[20480] = 25'b0000001010010011010010101;
    rom[20481] = 25'b0000001010010011011010001;
    rom[20482] = 25'b0000001010010011100001011;
    rom[20483] = 25'b0000001010010011101000101;
    rom[20484] = 25'b0000001010010011110000000;
    rom[20485] = 25'b0000001010010011110111001;
    rom[20486] = 25'b0000001010010011111110010;
    rom[20487] = 25'b0000001010010100000101011;
    rom[20488] = 25'b0000001010010100001100011;
    rom[20489] = 25'b0000001010010100010011011;
    rom[20490] = 25'b0000001010010100011010010;
    rom[20491] = 25'b0000001010010100100001001;
    rom[20492] = 25'b0000001010010100100111111;
    rom[20493] = 25'b0000001010010100101110110;
    rom[20494] = 25'b0000001010010100110101011;
    rom[20495] = 25'b0000001010010100111100000;
    rom[20496] = 25'b0000001010010101000010101;
    rom[20497] = 25'b0000001010010101001001001;
    rom[20498] = 25'b0000001010010101001111101;
    rom[20499] = 25'b0000001010010101010110000;
    rom[20500] = 25'b0000001010010101011100011;
    rom[20501] = 25'b0000001010010101100010101;
    rom[20502] = 25'b0000001010010101101000111;
    rom[20503] = 25'b0000001010010101101111001;
    rom[20504] = 25'b0000001010010101110101010;
    rom[20505] = 25'b0000001010010101111011011;
    rom[20506] = 25'b0000001010010110000001011;
    rom[20507] = 25'b0000001010010110000111011;
    rom[20508] = 25'b0000001010010110001101010;
    rom[20509] = 25'b0000001010010110010011001;
    rom[20510] = 25'b0000001010010110011001000;
    rom[20511] = 25'b0000001010010110011110101;
    rom[20512] = 25'b0000001010010110100100011;
    rom[20513] = 25'b0000001010010110101010001;
    rom[20514] = 25'b0000001010010110101111101;
    rom[20515] = 25'b0000001010010110110101001;
    rom[20516] = 25'b0000001010010110111010101;
    rom[20517] = 25'b0000001010010111000000000;
    rom[20518] = 25'b0000001010010111000101011;
    rom[20519] = 25'b0000001010010111001010101;
    rom[20520] = 25'b0000001010010111010000000;
    rom[20521] = 25'b0000001010010111010101001;
    rom[20522] = 25'b0000001010010111011010010;
    rom[20523] = 25'b0000001010010111011111011;
    rom[20524] = 25'b0000001010010111100100011;
    rom[20525] = 25'b0000001010010111101001011;
    rom[20526] = 25'b0000001010010111101110010;
    rom[20527] = 25'b0000001010010111110011001;
    rom[20528] = 25'b0000001010010111111000000;
    rom[20529] = 25'b0000001010010111111100110;
    rom[20530] = 25'b0000001010011000000001011;
    rom[20531] = 25'b0000001010011000000110000;
    rom[20532] = 25'b0000001010011000001010101;
    rom[20533] = 25'b0000001010011000001111001;
    rom[20534] = 25'b0000001010011000010011101;
    rom[20535] = 25'b0000001010011000011000000;
    rom[20536] = 25'b0000001010011000011100011;
    rom[20537] = 25'b0000001010011000100000101;
    rom[20538] = 25'b0000001010011000100100111;
    rom[20539] = 25'b0000001010011000101001001;
    rom[20540] = 25'b0000001010011000101101001;
    rom[20541] = 25'b0000001010011000110001010;
    rom[20542] = 25'b0000001010011000110101010;
    rom[20543] = 25'b0000001010011000111001010;
    rom[20544] = 25'b0000001010011000111101001;
    rom[20545] = 25'b0000001010011001000001000;
    rom[20546] = 25'b0000001010011001000100110;
    rom[20547] = 25'b0000001010011001001000100;
    rom[20548] = 25'b0000001010011001001100001;
    rom[20549] = 25'b0000001010011001001111110;
    rom[20550] = 25'b0000001010011001010011010;
    rom[20551] = 25'b0000001010011001010110111;
    rom[20552] = 25'b0000001010011001011010010;
    rom[20553] = 25'b0000001010011001011101101;
    rom[20554] = 25'b0000001010011001100001000;
    rom[20555] = 25'b0000001010011001100100010;
    rom[20556] = 25'b0000001010011001100111100;
    rom[20557] = 25'b0000001010011001101010101;
    rom[20558] = 25'b0000001010011001101101110;
    rom[20559] = 25'b0000001010011001110000110;
    rom[20560] = 25'b0000001010011001110011110;
    rom[20561] = 25'b0000001010011001110110101;
    rom[20562] = 25'b0000001010011001111001101;
    rom[20563] = 25'b0000001010011001111100011;
    rom[20564] = 25'b0000001010011001111111001;
    rom[20565] = 25'b0000001010011010000001111;
    rom[20566] = 25'b0000001010011010000100100;
    rom[20567] = 25'b0000001010011010000111001;
    rom[20568] = 25'b0000001010011010001001101;
    rom[20569] = 25'b0000001010011010001100000;
    rom[20570] = 25'b0000001010011010001110100;
    rom[20571] = 25'b0000001010011010010000111;
    rom[20572] = 25'b0000001010011010010011001;
    rom[20573] = 25'b0000001010011010010101011;
    rom[20574] = 25'b0000001010011010010111100;
    rom[20575] = 25'b0000001010011010011001110;
    rom[20576] = 25'b0000001010011010011011110;
    rom[20577] = 25'b0000001010011010011101110;
    rom[20578] = 25'b0000001010011010011111110;
    rom[20579] = 25'b0000001010011010100001101;
    rom[20580] = 25'b0000001010011010100011011;
    rom[20581] = 25'b0000001010011010100101010;
    rom[20582] = 25'b0000001010011010100111000;
    rom[20583] = 25'b0000001010011010101000101;
    rom[20584] = 25'b0000001010011010101010010;
    rom[20585] = 25'b0000001010011010101011111;
    rom[20586] = 25'b0000001010011010101101010;
    rom[20587] = 25'b0000001010011010101110110;
    rom[20588] = 25'b0000001010011010110000001;
    rom[20589] = 25'b0000001010011010110001011;
    rom[20590] = 25'b0000001010011010110010101;
    rom[20591] = 25'b0000001010011010110011111;
    rom[20592] = 25'b0000001010011010110101000;
    rom[20593] = 25'b0000001010011010110110001;
    rom[20594] = 25'b0000001010011010110111001;
    rom[20595] = 25'b0000001010011010111000000;
    rom[20596] = 25'b0000001010011010111001000;
    rom[20597] = 25'b0000001010011010111001111;
    rom[20598] = 25'b0000001010011010111010101;
    rom[20599] = 25'b0000001010011010111011011;
    rom[20600] = 25'b0000001010011010111100000;
    rom[20601] = 25'b0000001010011010111100101;
    rom[20602] = 25'b0000001010011010111101001;
    rom[20603] = 25'b0000001010011010111101101;
    rom[20604] = 25'b0000001010011010111110001;
    rom[20605] = 25'b0000001010011010111110100;
    rom[20606] = 25'b0000001010011010111110111;
    rom[20607] = 25'b0000001010011010111111000;
    rom[20608] = 25'b0000001010011010111111011;
    rom[20609] = 25'b0000001010011010111111011;
    rom[20610] = 25'b0000001010011010111111100;
    rom[20611] = 25'b0000001010011010111111100;
    rom[20612] = 25'b0000001010011010111111100;
    rom[20613] = 25'b0000001010011010111111011;
    rom[20614] = 25'b0000001010011010111111011;
    rom[20615] = 25'b0000001010011010111111000;
    rom[20616] = 25'b0000001010011010111110111;
    rom[20617] = 25'b0000001010011010111110100;
    rom[20618] = 25'b0000001010011010111110001;
    rom[20619] = 25'b0000001010011010111101101;
    rom[20620] = 25'b0000001010011010111101001;
    rom[20621] = 25'b0000001010011010111100101;
    rom[20622] = 25'b0000001010011010111100000;
    rom[20623] = 25'b0000001010011010111011011;
    rom[20624] = 25'b0000001010011010111010101;
    rom[20625] = 25'b0000001010011010111001111;
    rom[20626] = 25'b0000001010011010111001000;
    rom[20627] = 25'b0000001010011010111000000;
    rom[20628] = 25'b0000001010011010110111000;
    rom[20629] = 25'b0000001010011010110110000;
    rom[20630] = 25'b0000001010011010110101000;
    rom[20631] = 25'b0000001010011010110011110;
    rom[20632] = 25'b0000001010011010110010100;
    rom[20633] = 25'b0000001010011010110001011;
    rom[20634] = 25'b0000001010011010110000000;
    rom[20635] = 25'b0000001010011010101110101;
    rom[20636] = 25'b0000001010011010101101001;
    rom[20637] = 25'b0000001010011010101011101;
    rom[20638] = 25'b0000001010011010101010000;
    rom[20639] = 25'b0000001010011010101000100;
    rom[20640] = 25'b0000001010011010100110110;
    rom[20641] = 25'b0000001010011010100101000;
    rom[20642] = 25'b0000001010011010100011010;
    rom[20643] = 25'b0000001010011010100001011;
    rom[20644] = 25'b0000001010011010011111011;
    rom[20645] = 25'b0000001010011010011101011;
    rom[20646] = 25'b0000001010011010011011011;
    rom[20647] = 25'b0000001010011010011001011;
    rom[20648] = 25'b0000001010011010010111001;
    rom[20649] = 25'b0000001010011010010100111;
    rom[20650] = 25'b0000001010011010010010110;
    rom[20651] = 25'b0000001010011010010000010;
    rom[20652] = 25'b0000001010011010001101111;
    rom[20653] = 25'b0000001010011010001011011;
    rom[20654] = 25'b0000001010011010001000111;
    rom[20655] = 25'b0000001010011010000110011;
    rom[20656] = 25'b0000001010011010000011110;
    rom[20657] = 25'b0000001010011010000001000;
    rom[20658] = 25'b0000001010011001111110010;
    rom[20659] = 25'b0000001010011001111011100;
    rom[20660] = 25'b0000001010011001111000100;
    rom[20661] = 25'b0000001010011001110101101;
    rom[20662] = 25'b0000001010011001110010101;
    rom[20663] = 25'b0000001010011001101111101;
    rom[20664] = 25'b0000001010011001101100011;
    rom[20665] = 25'b0000001010011001101001010;
    rom[20666] = 25'b0000001010011001100110000;
    rom[20667] = 25'b0000001010011001100010110;
    rom[20668] = 25'b0000001010011001011111011;
    rom[20669] = 25'b0000001010011001011100000;
    rom[20670] = 25'b0000001010011001011000011;
    rom[20671] = 25'b0000001010011001010100111;
    rom[20672] = 25'b0000001010011001010001011;
    rom[20673] = 25'b0000001010011001001101101;
    rom[20674] = 25'b0000001010011001001010000;
    rom[20675] = 25'b0000001010011001000110001;
    rom[20676] = 25'b0000001010011001000010010;
    rom[20677] = 25'b0000001010011000111110011;
    rom[20678] = 25'b0000001010011000111010100;
    rom[20679] = 25'b0000001010011000110110011;
    rom[20680] = 25'b0000001010011000110010011;
    rom[20681] = 25'b0000001010011000101110010;
    rom[20682] = 25'b0000001010011000101010000;
    rom[20683] = 25'b0000001010011000100101110;
    rom[20684] = 25'b0000001010011000100001011;
    rom[20685] = 25'b0000001010011000011101000;
    rom[20686] = 25'b0000001010011000011000100;
    rom[20687] = 25'b0000001010011000010100000;
    rom[20688] = 25'b0000001010011000001111100;
    rom[20689] = 25'b0000001010011000001010111;
    rom[20690] = 25'b0000001010011000000110001;
    rom[20691] = 25'b0000001010011000000001011;
    rom[20692] = 25'b0000001010010111111100101;
    rom[20693] = 25'b0000001010010111110111101;
    rom[20694] = 25'b0000001010010111110010110;
    rom[20695] = 25'b0000001010010111101101110;
    rom[20696] = 25'b0000001010010111101000110;
    rom[20697] = 25'b0000001010010111100011101;
    rom[20698] = 25'b0000001010010111011110100;
    rom[20699] = 25'b0000001010010111011001010;
    rom[20700] = 25'b0000001010010111010011111;
    rom[20701] = 25'b0000001010010111001110100;
    rom[20702] = 25'b0000001010010111001001001;
    rom[20703] = 25'b0000001010010111000011101;
    rom[20704] = 25'b0000001010010110111110000;
    rom[20705] = 25'b0000001010010110111000100;
    rom[20706] = 25'b0000001010010110110010111;
    rom[20707] = 25'b0000001010010110101101000;
    rom[20708] = 25'b0000001010010110100111010;
    rom[20709] = 25'b0000001010010110100001100;
    rom[20710] = 25'b0000001010010110011011100;
    rom[20711] = 25'b0000001010010110010101101;
    rom[20712] = 25'b0000001010010110001111100;
    rom[20713] = 25'b0000001010010110001001100;
    rom[20714] = 25'b0000001010010110000011010;
    rom[20715] = 25'b0000001010010101111101000;
    rom[20716] = 25'b0000001010010101110110110;
    rom[20717] = 25'b0000001010010101110000100;
    rom[20718] = 25'b0000001010010101101010001;
    rom[20719] = 25'b0000001010010101100011101;
    rom[20720] = 25'b0000001010010101011101001;
    rom[20721] = 25'b0000001010010101010110100;
    rom[20722] = 25'b0000001010010101001111111;
    rom[20723] = 25'b0000001010010101001001001;
    rom[20724] = 25'b0000001010010101000010011;
    rom[20725] = 25'b0000001010010100111011101;
    rom[20726] = 25'b0000001010010100110100101;
    rom[20727] = 25'b0000001010010100101101101;
    rom[20728] = 25'b0000001010010100100110101;
    rom[20729] = 25'b0000001010010100011111101;
    rom[20730] = 25'b0000001010010100011000100;
    rom[20731] = 25'b0000001010010100010001010;
    rom[20732] = 25'b0000001010010100001010000;
    rom[20733] = 25'b0000001010010100000010110;
    rom[20734] = 25'b0000001010010011111011011;
    rom[20735] = 25'b0000001010010011110011111;
    rom[20736] = 25'b0000001010010011101100011;
    rom[20737] = 25'b0000001010010011100100111;
    rom[20738] = 25'b0000001010010011011101001;
    rom[20739] = 25'b0000001010010011010101100;
    rom[20740] = 25'b0000001010010011001101110;
    rom[20741] = 25'b0000001010010011000101111;
    rom[20742] = 25'b0000001010010010111110001;
    rom[20743] = 25'b0000001010010010110110001;
    rom[20744] = 25'b0000001010010010101110001;
    rom[20745] = 25'b0000001010010010100110001;
    rom[20746] = 25'b0000001010010010011110000;
    rom[20747] = 25'b0000001010010010010101110;
    rom[20748] = 25'b0000001010010010001101100;
    rom[20749] = 25'b0000001010010010000101010;
    rom[20750] = 25'b0000001010010001111100110;
    rom[20751] = 25'b0000001010010001110100011;
    rom[20752] = 25'b0000001010010001101011111;
    rom[20753] = 25'b0000001010010001100011010;
    rom[20754] = 25'b0000001010010001011010110;
    rom[20755] = 25'b0000001010010001010010000;
    rom[20756] = 25'b0000001010010001001001011;
    rom[20757] = 25'b0000001010010001000000100;
    rom[20758] = 25'b0000001010010000110111101;
    rom[20759] = 25'b0000001010010000101110110;
    rom[20760] = 25'b0000001010010000100101101;
    rom[20761] = 25'b0000001010010000011100101;
    rom[20762] = 25'b0000001010010000010011100;
    rom[20763] = 25'b0000001010010000001010011;
    rom[20764] = 25'b0000001010010000000001001;
    rom[20765] = 25'b0000001010001111110111111;
    rom[20766] = 25'b0000001010001111101110100;
    rom[20767] = 25'b0000001010001111100101000;
    rom[20768] = 25'b0000001010001111011011100;
    rom[20769] = 25'b0000001010001111010010000;
    rom[20770] = 25'b0000001010001111001000011;
    rom[20771] = 25'b0000001010001110111110110;
    rom[20772] = 25'b0000001010001110110101000;
    rom[20773] = 25'b0000001010001110101011001;
    rom[20774] = 25'b0000001010001110100001011;
    rom[20775] = 25'b0000001010001110010111011;
    rom[20776] = 25'b0000001010001110001101100;
    rom[20777] = 25'b0000001010001110000011011;
    rom[20778] = 25'b0000001010001101111001010;
    rom[20779] = 25'b0000001010001101101111001;
    rom[20780] = 25'b0000001010001101100100111;
    rom[20781] = 25'b0000001010001101011010100;
    rom[20782] = 25'b0000001010001101010000001;
    rom[20783] = 25'b0000001010001101000101110;
    rom[20784] = 25'b0000001010001100111011010;
    rom[20785] = 25'b0000001010001100110000110;
    rom[20786] = 25'b0000001010001100100110001;
    rom[20787] = 25'b0000001010001100011011011;
    rom[20788] = 25'b0000001010001100010000101;
    rom[20789] = 25'b0000001010001100000110000;
    rom[20790] = 25'b0000001010001011111011000;
    rom[20791] = 25'b0000001010001011110000001;
    rom[20792] = 25'b0000001010001011100101001;
    rom[20793] = 25'b0000001010001011011010001;
    rom[20794] = 25'b0000001010001011001111000;
    rom[20795] = 25'b0000001010001011000011111;
    rom[20796] = 25'b0000001010001010111000101;
    rom[20797] = 25'b0000001010001010101101011;
    rom[20798] = 25'b0000001010001010100001111;
    rom[20799] = 25'b0000001010001010010110100;
    rom[20800] = 25'b0000001010001010001011000;
    rom[20801] = 25'b0000001010001001111111100;
    rom[20802] = 25'b0000001010001001110011111;
    rom[20803] = 25'b0000001010001001101000010;
    rom[20804] = 25'b0000001010001001011100100;
    rom[20805] = 25'b0000001010001001010000101;
    rom[20806] = 25'b0000001010001001000100111;
    rom[20807] = 25'b0000001010001000111000111;
    rom[20808] = 25'b0000001010001000101100111;
    rom[20809] = 25'b0000001010001000100000110;
    rom[20810] = 25'b0000001010001000010100110;
    rom[20811] = 25'b0000001010001000001000100;
    rom[20812] = 25'b0000001010000111111100010;
    rom[20813] = 25'b0000001010000111110000000;
    rom[20814] = 25'b0000001010000111100011101;
    rom[20815] = 25'b0000001010000111010111001;
    rom[20816] = 25'b0000001010000111001010101;
    rom[20817] = 25'b0000001010000110111110001;
    rom[20818] = 25'b0000001010000110110001100;
    rom[20819] = 25'b0000001010000110100100111;
    rom[20820] = 25'b0000001010000110011000001;
    rom[20821] = 25'b0000001010000110001011010;
    rom[20822] = 25'b0000001010000101111110100;
    rom[20823] = 25'b0000001010000101110001100;
    rom[20824] = 25'b0000001010000101100100100;
    rom[20825] = 25'b0000001010000101010111011;
    rom[20826] = 25'b0000001010000101001010011;
    rom[20827] = 25'b0000001010000100111101001;
    rom[20828] = 25'b0000001010000100101111111;
    rom[20829] = 25'b0000001010000100100010101;
    rom[20830] = 25'b0000001010000100010101010;
    rom[20831] = 25'b0000001010000100000111110;
    rom[20832] = 25'b0000001010000011111010011;
    rom[20833] = 25'b0000001010000011101100101;
    rom[20834] = 25'b0000001010000011011111001;
    rom[20835] = 25'b0000001010000011010001011;
    rom[20836] = 25'b0000001010000011000011110;
    rom[20837] = 25'b0000001010000010110101111;
    rom[20838] = 25'b0000001010000010101000000;
    rom[20839] = 25'b0000001010000010011010000;
    rom[20840] = 25'b0000001010000010001100000;
    rom[20841] = 25'b0000001010000001111101111;
    rom[20842] = 25'b0000001010000001101111111;
    rom[20843] = 25'b0000001010000001100001101;
    rom[20844] = 25'b0000001010000001010011011;
    rom[20845] = 25'b0000001010000001000101000;
    rom[20846] = 25'b0000001010000000110110101;
    rom[20847] = 25'b0000001010000000101000010;
    rom[20848] = 25'b0000001010000000011001110;
    rom[20849] = 25'b0000001010000000001011001;
    rom[20850] = 25'b0000001001111111111100100;
    rom[20851] = 25'b0000001001111111101101111;
    rom[20852] = 25'b0000001001111111011111001;
    rom[20853] = 25'b0000001001111111010000010;
    rom[20854] = 25'b0000001001111111000001011;
    rom[20855] = 25'b0000001001111110110010011;
    rom[20856] = 25'b0000001001111110100011011;
    rom[20857] = 25'b0000001001111110010100010;
    rom[20858] = 25'b0000001001111110000101001;
    rom[20859] = 25'b0000001001111101110101111;
    rom[20860] = 25'b0000001001111101100110110;
    rom[20861] = 25'b0000001001111101010111011;
    rom[20862] = 25'b0000001001111101001000000;
    rom[20863] = 25'b0000001001111100111000100;
    rom[20864] = 25'b0000001001111100101001000;
    rom[20865] = 25'b0000001001111100011001011;
    rom[20866] = 25'b0000001001111100001001110;
    rom[20867] = 25'b0000001001111011111010000;
    rom[20868] = 25'b0000001001111011101010010;
    rom[20869] = 25'b0000001001111011011010011;
    rom[20870] = 25'b0000001001111011001010100;
    rom[20871] = 25'b0000001001111010111010100;
    rom[20872] = 25'b0000001001111010101010100;
    rom[20873] = 25'b0000001001111010011010011;
    rom[20874] = 25'b0000001001111010001010010;
    rom[20875] = 25'b0000001001111001111010000;
    rom[20876] = 25'b0000001001111001101001110;
    rom[20877] = 25'b0000001001111001011001011;
    rom[20878] = 25'b0000001001111001001001000;
    rom[20879] = 25'b0000001001111000111000100;
    rom[20880] = 25'b0000001001111000101000000;
    rom[20881] = 25'b0000001001111000010111011;
    rom[20882] = 25'b0000001001111000000110110;
    rom[20883] = 25'b0000001001110111110110000;
    rom[20884] = 25'b0000001001110111100101010;
    rom[20885] = 25'b0000001001110111010100011;
    rom[20886] = 25'b0000001001110111000011011;
    rom[20887] = 25'b0000001001110110110010100;
    rom[20888] = 25'b0000001001110110100001011;
    rom[20889] = 25'b0000001001110110010000010;
    rom[20890] = 25'b0000001001110101111111001;
    rom[20891] = 25'b0000001001110101101101111;
    rom[20892] = 25'b0000001001110101011100101;
    rom[20893] = 25'b0000001001110101001011010;
    rom[20894] = 25'b0000001001110100111001111;
    rom[20895] = 25'b0000001001110100101000010;
    rom[20896] = 25'b0000001001110100010110110;
    rom[20897] = 25'b0000001001110100000101001;
    rom[20898] = 25'b0000001001110011110011011;
    rom[20899] = 25'b0000001001110011100001101;
    rom[20900] = 25'b0000001001110011001111111;
    rom[20901] = 25'b0000001001110010111110000;
    rom[20902] = 25'b0000001001110010101100001;
    rom[20903] = 25'b0000001001110010011010000;
    rom[20904] = 25'b0000001001110010001000000;
    rom[20905] = 25'b0000001001110001110101111;
    rom[20906] = 25'b0000001001110001100011110;
    rom[20907] = 25'b0000001001110001010001100;
    rom[20908] = 25'b0000001001110000111111001;
    rom[20909] = 25'b0000001001110000101100110;
    rom[20910] = 25'b0000001001110000011010010;
    rom[20911] = 25'b0000001001110000000111110;
    rom[20912] = 25'b0000001001101111110101010;
    rom[20913] = 25'b0000001001101111100010100;
    rom[20914] = 25'b0000001001101111001111111;
    rom[20915] = 25'b0000001001101110111101001;
    rom[20916] = 25'b0000001001101110101010011;
    rom[20917] = 25'b0000001001101110010111011;
    rom[20918] = 25'b0000001001101110000100011;
    rom[20919] = 25'b0000001001101101110001100;
    rom[20920] = 25'b0000001001101101011110010;
    rom[20921] = 25'b0000001001101101001011001;
    rom[20922] = 25'b0000001001101100111000000;
    rom[20923] = 25'b0000001001101100100100110;
    rom[20924] = 25'b0000001001101100010001011;
    rom[20925] = 25'b0000001001101011111101111;
    rom[20926] = 25'b0000001001101011101010100;
    rom[20927] = 25'b0000001001101011010111000;
    rom[20928] = 25'b0000001001101011000011011;
    rom[20929] = 25'b0000001001101010101111110;
    rom[20930] = 25'b0000001001101010011100001;
    rom[20931] = 25'b0000001001101010001000010;
    rom[20932] = 25'b0000001001101001110100011;
    rom[20933] = 25'b0000001001101001100000100;
    rom[20934] = 25'b0000001001101001001100100;
    rom[20935] = 25'b0000001001101000111000011;
    rom[20936] = 25'b0000001001101000100100011;
    rom[20937] = 25'b0000001001101000010000001;
    rom[20938] = 25'b0000001001100111111100000;
    rom[20939] = 25'b0000001001100111100111101;
    rom[20940] = 25'b0000001001100111010011010;
    rom[20941] = 25'b0000001001100110111110111;
    rom[20942] = 25'b0000001001100110101010011;
    rom[20943] = 25'b0000001001100110010101111;
    rom[20944] = 25'b0000001001100110000001010;
    rom[20945] = 25'b0000001001100101101100100;
    rom[20946] = 25'b0000001001100101010111111;
    rom[20947] = 25'b0000001001100101000011000;
    rom[20948] = 25'b0000001001100100101110001;
    rom[20949] = 25'b0000001001100100011001010;
    rom[20950] = 25'b0000001001100100000100010;
    rom[20951] = 25'b0000001001100011101111001;
    rom[20952] = 25'b0000001001100011011010000;
    rom[20953] = 25'b0000001001100011000100111;
    rom[20954] = 25'b0000001001100010101111101;
    rom[20955] = 25'b0000001001100010011010011;
    rom[20956] = 25'b0000001001100010000101000;
    rom[20957] = 25'b0000001001100001101111100;
    rom[20958] = 25'b0000001001100001011010000;
    rom[20959] = 25'b0000001001100001000100011;
    rom[20960] = 25'b0000001001100000101110110;
    rom[20961] = 25'b0000001001100000011001001;
    rom[20962] = 25'b0000001001100000000011011;
    rom[20963] = 25'b0000001001011111101101100;
    rom[20964] = 25'b0000001001011111010111101;
    rom[20965] = 25'b0000001001011111000001101;
    rom[20966] = 25'b0000001001011110101011101;
    rom[20967] = 25'b0000001001011110010101100;
    rom[20968] = 25'b0000001001011101111111011;
    rom[20969] = 25'b0000001001011101101001010;
    rom[20970] = 25'b0000001001011101010010111;
    rom[20971] = 25'b0000001001011100111100101;
    rom[20972] = 25'b0000001001011100100110010;
    rom[20973] = 25'b0000001001011100001111110;
    rom[20974] = 25'b0000001001011011111001001;
    rom[20975] = 25'b0000001001011011100010101;
    rom[20976] = 25'b0000001001011011001100000;
    rom[20977] = 25'b0000001001011010110101010;
    rom[20978] = 25'b0000001001011010011110100;
    rom[20979] = 25'b0000001001011010000111101;
    rom[20980] = 25'b0000001001011001110000110;
    rom[20981] = 25'b0000001001011001011001110;
    rom[20982] = 25'b0000001001011001000010110;
    rom[20983] = 25'b0000001001011000101011101;
    rom[20984] = 25'b0000001001011000010100100;
    rom[20985] = 25'b0000001001010111111101010;
    rom[20986] = 25'b0000001001010111100101111;
    rom[20987] = 25'b0000001001010111001110100;
    rom[20988] = 25'b0000001001010110110111001;
    rom[20989] = 25'b0000001001010110011111101;
    rom[20990] = 25'b0000001001010110001000001;
    rom[20991] = 25'b0000001001010101110000100;
    rom[20992] = 25'b0000001001010101011000111;
    rom[20993] = 25'b0000001001010101000001001;
    rom[20994] = 25'b0000001001010100101001011;
    rom[20995] = 25'b0000001001010100010001011;
    rom[20996] = 25'b0000001001010011111001100;
    rom[20997] = 25'b0000001001010011100001100;
    rom[20998] = 25'b0000001001010011001001011;
    rom[20999] = 25'b0000001001010010110001011;
    rom[21000] = 25'b0000001001010010011001001;
    rom[21001] = 25'b0000001001010010000000111;
    rom[21002] = 25'b0000001001010001101000101;
    rom[21003] = 25'b0000001001010001010000010;
    rom[21004] = 25'b0000001001010000110111110;
    rom[21005] = 25'b0000001001010000011111010;
    rom[21006] = 25'b0000001001010000000110110;
    rom[21007] = 25'b0000001001001111101110000;
    rom[21008] = 25'b0000001001001111010101011;
    rom[21009] = 25'b0000001001001110111100101;
    rom[21010] = 25'b0000001001001110100011110;
    rom[21011] = 25'b0000001001001110001011000;
    rom[21012] = 25'b0000001001001101110010000;
    rom[21013] = 25'b0000001001001101011001000;
    rom[21014] = 25'b0000001001001100111111111;
    rom[21015] = 25'b0000001001001100100110110;
    rom[21016] = 25'b0000001001001100001101100;
    rom[21017] = 25'b0000001001001011110100010;
    rom[21018] = 25'b0000001001001011011010111;
    rom[21019] = 25'b0000001001001011000001100;
    rom[21020] = 25'b0000001001001010101000001;
    rom[21021] = 25'b0000001001001010001110100;
    rom[21022] = 25'b0000001001001001110101000;
    rom[21023] = 25'b0000001001001001011011011;
    rom[21024] = 25'b0000001001001001000001101;
    rom[21025] = 25'b0000001001001000100111111;
    rom[21026] = 25'b0000001001001000001110000;
    rom[21027] = 25'b0000001001000111110100001;
    rom[21028] = 25'b0000001001000111011010001;
    rom[21029] = 25'b0000001001000111000000001;
    rom[21030] = 25'b0000001001000110100110000;
    rom[21031] = 25'b0000001001000110001011111;
    rom[21032] = 25'b0000001001000101110001101;
    rom[21033] = 25'b0000001001000101010111011;
    rom[21034] = 25'b0000001001000100111101000;
    rom[21035] = 25'b0000001001000100100010101;
    rom[21036] = 25'b0000001001000100001000001;
    rom[21037] = 25'b0000001001000011101101101;
    rom[21038] = 25'b0000001001000011010011000;
    rom[21039] = 25'b0000001001000010111000011;
    rom[21040] = 25'b0000001001000010011101101;
    rom[21041] = 25'b0000001001000010000010111;
    rom[21042] = 25'b0000001001000001100111111;
    rom[21043] = 25'b0000001001000001001101000;
    rom[21044] = 25'b0000001001000000110010000;
    rom[21045] = 25'b0000001001000000010111000;
    rom[21046] = 25'b0000001000111111111011111;
    rom[21047] = 25'b0000001000111111100000110;
    rom[21048] = 25'b0000001000111111000101100;
    rom[21049] = 25'b0000001000111110101010001;
    rom[21050] = 25'b0000001000111110001110110;
    rom[21051] = 25'b0000001000111101110011011;
    rom[21052] = 25'b0000001000111101010111111;
    rom[21053] = 25'b0000001000111100111100011;
    rom[21054] = 25'b0000001000111100100000110;
    rom[21055] = 25'b0000001000111100000101001;
    rom[21056] = 25'b0000001000111011101001011;
    rom[21057] = 25'b0000001000111011001101100;
    rom[21058] = 25'b0000001000111010110001101;
    rom[21059] = 25'b0000001000111010010101110;
    rom[21060] = 25'b0000001000111001111001110;
    rom[21061] = 25'b0000001000111001011101101;
    rom[21062] = 25'b0000001000111001000001100;
    rom[21063] = 25'b0000001000111000100101010;
    rom[21064] = 25'b0000001000111000001001001;
    rom[21065] = 25'b0000001000110111101100110;
    rom[21066] = 25'b0000001000110111010000011;
    rom[21067] = 25'b0000001000110110110100000;
    rom[21068] = 25'b0000001000110110010111100;
    rom[21069] = 25'b0000001000110101111010111;
    rom[21070] = 25'b0000001000110101011110010;
    rom[21071] = 25'b0000001000110101000001100;
    rom[21072] = 25'b0000001000110100100100110;
    rom[21073] = 25'b0000001000110100001000000;
    rom[21074] = 25'b0000001000110011101011001;
    rom[21075] = 25'b0000001000110011001110001;
    rom[21076] = 25'b0000001000110010110001001;
    rom[21077] = 25'b0000001000110010010100001;
    rom[21078] = 25'b0000001000110001110111000;
    rom[21079] = 25'b0000001000110001011001110;
    rom[21080] = 25'b0000001000110000111100100;
    rom[21081] = 25'b0000001000110000011111010;
    rom[21082] = 25'b0000001000110000000001110;
    rom[21083] = 25'b0000001000101111100100010;
    rom[21084] = 25'b0000001000101111000110110;
    rom[21085] = 25'b0000001000101110101001010;
    rom[21086] = 25'b0000001000101110001011100;
    rom[21087] = 25'b0000001000101101101101111;
    rom[21088] = 25'b0000001000101101010000001;
    rom[21089] = 25'b0000001000101100110010010;
    rom[21090] = 25'b0000001000101100010100011;
    rom[21091] = 25'b0000001000101011110110011;
    rom[21092] = 25'b0000001000101011011000100;
    rom[21093] = 25'b0000001000101010111010011;
    rom[21094] = 25'b0000001000101010011100010;
    rom[21095] = 25'b0000001000101001111110000;
    rom[21096] = 25'b0000001000101001011111110;
    rom[21097] = 25'b0000001000101001000001011;
    rom[21098] = 25'b0000001000101000100011000;
    rom[21099] = 25'b0000001000101000000100100;
    rom[21100] = 25'b0000001000100111100110000;
    rom[21101] = 25'b0000001000100111000111011;
    rom[21102] = 25'b0000001000100110101000110;
    rom[21103] = 25'b0000001000100110001010000;
    rom[21104] = 25'b0000001000100101101011010;
    rom[21105] = 25'b0000001000100101001100100;
    rom[21106] = 25'b0000001000100100101101101;
    rom[21107] = 25'b0000001000100100001110100;
    rom[21108] = 25'b0000001000100011101111100;
    rom[21109] = 25'b0000001000100011010000100;
    rom[21110] = 25'b0000001000100010110001011;
    rom[21111] = 25'b0000001000100010010010001;
    rom[21112] = 25'b0000001000100001110010110;
    rom[21113] = 25'b0000001000100001010011100;
    rom[21114] = 25'b0000001000100000110100001;
    rom[21115] = 25'b0000001000100000010100101;
    rom[21116] = 25'b0000001000011111110101001;
    rom[21117] = 25'b0000001000011111010101100;
    rom[21118] = 25'b0000001000011110110101111;
    rom[21119] = 25'b0000001000011110010110001;
    rom[21120] = 25'b0000001000011101110110011;
    rom[21121] = 25'b0000001000011101010110100;
    rom[21122] = 25'b0000001000011100110110101;
    rom[21123] = 25'b0000001000011100010110101;
    rom[21124] = 25'b0000001000011011110110101;
    rom[21125] = 25'b0000001000011011010110101;
    rom[21126] = 25'b0000001000011010110110011;
    rom[21127] = 25'b0000001000011010010110001;
    rom[21128] = 25'b0000001000011001110101111;
    rom[21129] = 25'b0000001000011001010101100;
    rom[21130] = 25'b0000001000011000110101001;
    rom[21131] = 25'b0000001000011000010100110;
    rom[21132] = 25'b0000001000010111110100001;
    rom[21133] = 25'b0000001000010111010011100;
    rom[21134] = 25'b0000001000010110110010111;
    rom[21135] = 25'b0000001000010110010010001;
    rom[21136] = 25'b0000001000010101110001011;
    rom[21137] = 25'b0000001000010101010000101;
    rom[21138] = 25'b0000001000010100101111101;
    rom[21139] = 25'b0000001000010100001110101;
    rom[21140] = 25'b0000001000010011101101110;
    rom[21141] = 25'b0000001000010011001100101;
    rom[21142] = 25'b0000001000010010101011100;
    rom[21143] = 25'b0000001000010010001010010;
    rom[21144] = 25'b0000001000010001101001000;
    rom[21145] = 25'b0000001000010001000111101;
    rom[21146] = 25'b0000001000010000100110010;
    rom[21147] = 25'b0000001000010000000100110;
    rom[21148] = 25'b0000001000001111100011010;
    rom[21149] = 25'b0000001000001111000001101;
    rom[21150] = 25'b0000001000001110100000000;
    rom[21151] = 25'b0000001000001101111110011;
    rom[21152] = 25'b0000001000001101011100100;
    rom[21153] = 25'b0000001000001100111010110;
    rom[21154] = 25'b0000001000001100011000110;
    rom[21155] = 25'b0000001000001011110110110;
    rom[21156] = 25'b0000001000001011010100111;
    rom[21157] = 25'b0000001000001010110010110;
    rom[21158] = 25'b0000001000001010010000100;
    rom[21159] = 25'b0000001000001001101110011;
    rom[21160] = 25'b0000001000001001001100001;
    rom[21161] = 25'b0000001000001000101001110;
    rom[21162] = 25'b0000001000001000000111011;
    rom[21163] = 25'b0000001000000111100100111;
    rom[21164] = 25'b0000001000000111000010011;
    rom[21165] = 25'b0000001000000110011111110;
    rom[21166] = 25'b0000001000000101111101001;
    rom[21167] = 25'b0000001000000101011010100;
    rom[21168] = 25'b0000001000000100110111101;
    rom[21169] = 25'b0000001000000100010100111;
    rom[21170] = 25'b0000001000000011110010000;
    rom[21171] = 25'b0000001000000011001111000;
    rom[21172] = 25'b0000001000000010101100000;
    rom[21173] = 25'b0000001000000010001001000;
    rom[21174] = 25'b0000001000000001100101111;
    rom[21175] = 25'b0000001000000001000010101;
    rom[21176] = 25'b0000001000000000011111011;
    rom[21177] = 25'b0000000111111111111100000;
    rom[21178] = 25'b0000000111111111011000101;
    rom[21179] = 25'b0000000111111110110101010;
    rom[21180] = 25'b0000000111111110010001101;
    rom[21181] = 25'b0000000111111101101110001;
    rom[21182] = 25'b0000000111111101001010100;
    rom[21183] = 25'b0000000111111100100110111;
    rom[21184] = 25'b0000000111111100000011000;
    rom[21185] = 25'b0000000111111011011111010;
    rom[21186] = 25'b0000000111111010111011011;
    rom[21187] = 25'b0000000111111010010111100;
    rom[21188] = 25'b0000000111111001110011011;
    rom[21189] = 25'b0000000111111001001111011;
    rom[21190] = 25'b0000000111111000101011010;
    rom[21191] = 25'b0000000111111000000111001;
    rom[21192] = 25'b0000000111110111100010111;
    rom[21193] = 25'b0000000111110110111110100;
    rom[21194] = 25'b0000000111110110011010010;
    rom[21195] = 25'b0000000111110101110101110;
    rom[21196] = 25'b0000000111110101010001010;
    rom[21197] = 25'b0000000111110100101100110;
    rom[21198] = 25'b0000000111110100001000000;
    rom[21199] = 25'b0000000111110011100011100;
    rom[21200] = 25'b0000000111110010111110101;
    rom[21201] = 25'b0000000111110010011001111;
    rom[21202] = 25'b0000000111110001110101001;
    rom[21203] = 25'b0000000111110001010000001;
    rom[21204] = 25'b0000000111110000101011010;
    rom[21205] = 25'b0000000111110000000110001;
    rom[21206] = 25'b0000000111101111100001000;
    rom[21207] = 25'b0000000111101110111011111;
    rom[21208] = 25'b0000000111101110010110101;
    rom[21209] = 25'b0000000111101101110001011;
    rom[21210] = 25'b0000000111101101001100000;
    rom[21211] = 25'b0000000111101100100110101;
    rom[21212] = 25'b0000000111101100000001001;
    rom[21213] = 25'b0000000111101011011011101;
    rom[21214] = 25'b0000000111101010110110000;
    rom[21215] = 25'b0000000111101010010000011;
    rom[21216] = 25'b0000000111101001101010101;
    rom[21217] = 25'b0000000111101001000100111;
    rom[21218] = 25'b0000000111101000011111001;
    rom[21219] = 25'b0000000111100111111001010;
    rom[21220] = 25'b0000000111100111010011010;
    rom[21221] = 25'b0000000111100110101101010;
    rom[21222] = 25'b0000000111100110000111001;
    rom[21223] = 25'b0000000111100101100001001;
    rom[21224] = 25'b0000000111100100111010111;
    rom[21225] = 25'b0000000111100100010100101;
    rom[21226] = 25'b0000000111100011101110010;
    rom[21227] = 25'b0000000111100011000111111;
    rom[21228] = 25'b0000000111100010100001011;
    rom[21229] = 25'b0000000111100001111011000;
    rom[21230] = 25'b0000000111100001010100011;
    rom[21231] = 25'b0000000111100000101101111;
    rom[21232] = 25'b0000000111100000000111001;
    rom[21233] = 25'b0000000111011111100000011;
    rom[21234] = 25'b0000000111011110111001100;
    rom[21235] = 25'b0000000111011110010010110;
    rom[21236] = 25'b0000000111011101101011110;
    rom[21237] = 25'b0000000111011101000100111;
    rom[21238] = 25'b0000000111011100011101110;
    rom[21239] = 25'b0000000111011011110110101;
    rom[21240] = 25'b0000000111011011001111100;
    rom[21241] = 25'b0000000111011010101000010;
    rom[21242] = 25'b0000000111011010000001000;
    rom[21243] = 25'b0000000111011001011001101;
    rom[21244] = 25'b0000000111011000110010010;
    rom[21245] = 25'b0000000111011000001010111;
    rom[21246] = 25'b0000000111010111100011010;
    rom[21247] = 25'b0000000111010110111011110;
    rom[21248] = 25'b0000000111010110010100001;
    rom[21249] = 25'b0000000111010101101100011;
    rom[21250] = 25'b0000000111010101000100101;
    rom[21251] = 25'b0000000111010100011100111;
    rom[21252] = 25'b0000000111010011110100111;
    rom[21253] = 25'b0000000111010011001101000;
    rom[21254] = 25'b0000000111010010100101000;
    rom[21255] = 25'b0000000111010001111100111;
    rom[21256] = 25'b0000000111010001010100110;
    rom[21257] = 25'b0000000111010000101100101;
    rom[21258] = 25'b0000000111010000000100011;
    rom[21259] = 25'b0000000111001111011100001;
    rom[21260] = 25'b0000000111001110110011101;
    rom[21261] = 25'b0000000111001110001011011;
    rom[21262] = 25'b0000000111001101100010110;
    rom[21263] = 25'b0000000111001100111010010;
    rom[21264] = 25'b0000000111001100010001101;
    rom[21265] = 25'b0000000111001011101001000;
    rom[21266] = 25'b0000000111001011000000011;
    rom[21267] = 25'b0000000111001010010111101;
    rom[21268] = 25'b0000000111001001101110110;
    rom[21269] = 25'b0000000111001001000101110;
    rom[21270] = 25'b0000000111001000011100111;
    rom[21271] = 25'b0000000111000111110011111;
    rom[21272] = 25'b0000000111000111001010110;
    rom[21273] = 25'b0000000111000110100001101;
    rom[21274] = 25'b0000000111000101111000011;
    rom[21275] = 25'b0000000111000101001111010;
    rom[21276] = 25'b0000000111000100100101111;
    rom[21277] = 25'b0000000111000011111100100;
    rom[21278] = 25'b0000000111000011010011001;
    rom[21279] = 25'b0000000111000010101001101;
    rom[21280] = 25'b0000000111000010000000001;
    rom[21281] = 25'b0000000111000001010110100;
    rom[21282] = 25'b0000000111000000101100111;
    rom[21283] = 25'b0000000111000000000011001;
    rom[21284] = 25'b0000000110111111011001011;
    rom[21285] = 25'b0000000110111110101111100;
    rom[21286] = 25'b0000000110111110000101101;
    rom[21287] = 25'b0000000110111101011011101;
    rom[21288] = 25'b0000000110111100110001101;
    rom[21289] = 25'b0000000110111100000111100;
    rom[21290] = 25'b0000000110111011011101011;
    rom[21291] = 25'b0000000110111010110011001;
    rom[21292] = 25'b0000000110111010001001000;
    rom[21293] = 25'b0000000110111001011110101;
    rom[21294] = 25'b0000000110111000110100010;
    rom[21295] = 25'b0000000110111000001001111;
    rom[21296] = 25'b0000000110110111011111011;
    rom[21297] = 25'b0000000110110110110100110;
    rom[21298] = 25'b0000000110110110001010010;
    rom[21299] = 25'b0000000110110101011111100;
    rom[21300] = 25'b0000000110110100110100111;
    rom[21301] = 25'b0000000110110100001010001;
    rom[21302] = 25'b0000000110110011011111010;
    rom[21303] = 25'b0000000110110010110100011;
    rom[21304] = 25'b0000000110110010001001011;
    rom[21305] = 25'b0000000110110001011110011;
    rom[21306] = 25'b0000000110110000110011010;
    rom[21307] = 25'b0000000110110000001000001;
    rom[21308] = 25'b0000000110101111011101000;
    rom[21309] = 25'b0000000110101110110001110;
    rom[21310] = 25'b0000000110101110000110011;
    rom[21311] = 25'b0000000110101101011011001;
    rom[21312] = 25'b0000000110101100101111101;
    rom[21313] = 25'b0000000110101100000100001;
    rom[21314] = 25'b0000000110101011011000101;
    rom[21315] = 25'b0000000110101010101101000;
    rom[21316] = 25'b0000000110101010000001011;
    rom[21317] = 25'b0000000110101001010101110;
    rom[21318] = 25'b0000000110101000101001111;
    rom[21319] = 25'b0000000110100111111110001;
    rom[21320] = 25'b0000000110100111010010010;
    rom[21321] = 25'b0000000110100110100110010;
    rom[21322] = 25'b0000000110100101111010010;
    rom[21323] = 25'b0000000110100101001110010;
    rom[21324] = 25'b0000000110100100100010001;
    rom[21325] = 25'b0000000110100011110101111;
    rom[21326] = 25'b0000000110100011001001110;
    rom[21327] = 25'b0000000110100010011101100;
    rom[21328] = 25'b0000000110100001110001001;
    rom[21329] = 25'b0000000110100001000100101;
    rom[21330] = 25'b0000000110100000011000010;
    rom[21331] = 25'b0000000110011111101011101;
    rom[21332] = 25'b0000000110011110111111001;
    rom[21333] = 25'b0000000110011110010010100;
    rom[21334] = 25'b0000000110011101100101111;
    rom[21335] = 25'b0000000110011100111001001;
    rom[21336] = 25'b0000000110011100001100010;
    rom[21337] = 25'b0000000110011011011111100;
    rom[21338] = 25'b0000000110011010110010100;
    rom[21339] = 25'b0000000110011010000101100;
    rom[21340] = 25'b0000000110011001011000100;
    rom[21341] = 25'b0000000110011000101011011;
    rom[21342] = 25'b0000000110010111111110010;
    rom[21343] = 25'b0000000110010111010001000;
    rom[21344] = 25'b0000000110010110100011110;
    rom[21345] = 25'b0000000110010101110110100;
    rom[21346] = 25'b0000000110010101001001001;
    rom[21347] = 25'b0000000110010100011011101;
    rom[21348] = 25'b0000000110010011101110001;
    rom[21349] = 25'b0000000110010011000000101;
    rom[21350] = 25'b0000000110010010010011000;
    rom[21351] = 25'b0000000110010001100101011;
    rom[21352] = 25'b0000000110010000110111101;
    rom[21353] = 25'b0000000110010000001001111;
    rom[21354] = 25'b0000000110001111011100001;
    rom[21355] = 25'b0000000110001110101110010;
    rom[21356] = 25'b0000000110001110000000010;
    rom[21357] = 25'b0000000110001101010010010;
    rom[21358] = 25'b0000000110001100100100010;
    rom[21359] = 25'b0000000110001011110110000;
    rom[21360] = 25'b0000000110001011000111111;
    rom[21361] = 25'b0000000110001010011001110;
    rom[21362] = 25'b0000000110001001101011011;
    rom[21363] = 25'b0000000110001000111101000;
    rom[21364] = 25'b0000000110001000001110110;
    rom[21365] = 25'b0000000110000111100000010;
    rom[21366] = 25'b0000000110000110110001110;
    rom[21367] = 25'b0000000110000110000011010;
    rom[21368] = 25'b0000000110000101010100101;
    rom[21369] = 25'b0000000110000100100101111;
    rom[21370] = 25'b0000000110000011110111001;
    rom[21371] = 25'b0000000110000011001000011;
    rom[21372] = 25'b0000000110000010011001101;
    rom[21373] = 25'b0000000110000001101010101;
    rom[21374] = 25'b0000000110000000111011110;
    rom[21375] = 25'b0000000110000000001100110;
    rom[21376] = 25'b0000000101111111011101101;
    rom[21377] = 25'b0000000101111110101110100;
    rom[21378] = 25'b0000000101111101111111011;
    rom[21379] = 25'b0000000101111101010000001;
    rom[21380] = 25'b0000000101111100100000111;
    rom[21381] = 25'b0000000101111011110001100;
    rom[21382] = 25'b0000000101111011000010000;
    rom[21383] = 25'b0000000101111010010010101;
    rom[21384] = 25'b0000000101111001100011001;
    rom[21385] = 25'b0000000101111000110011100;
    rom[21386] = 25'b0000000101111000000011111;
    rom[21387] = 25'b0000000101110111010100010;
    rom[21388] = 25'b0000000101110110100100101;
    rom[21389] = 25'b0000000101110101110100110;
    rom[21390] = 25'b0000000101110101000101000;
    rom[21391] = 25'b0000000101110100010101000;
    rom[21392] = 25'b0000000101110011100101001;
    rom[21393] = 25'b0000000101110010110101001;
    rom[21394] = 25'b0000000101110010000101000;
    rom[21395] = 25'b0000000101110001010101000;
    rom[21396] = 25'b0000000101110000100100110;
    rom[21397] = 25'b0000000101101111110100100;
    rom[21398] = 25'b0000000101101111000100010;
    rom[21399] = 25'b0000000101101110010011111;
    rom[21400] = 25'b0000000101101101100011100;
    rom[21401] = 25'b0000000101101100110011001;
    rom[21402] = 25'b0000000101101100000010101;
    rom[21403] = 25'b0000000101101011010010000;
    rom[21404] = 25'b0000000101101010100001011;
    rom[21405] = 25'b0000000101101001110000110;
    rom[21406] = 25'b0000000101101001000000001;
    rom[21407] = 25'b0000000101101000001111010;
    rom[21408] = 25'b0000000101100111011110011;
    rom[21409] = 25'b0000000101100110101101100;
    rom[21410] = 25'b0000000101100101111100101;
    rom[21411] = 25'b0000000101100101001011101;
    rom[21412] = 25'b0000000101100100011010100;
    rom[21413] = 25'b0000000101100011101001100;
    rom[21414] = 25'b0000000101100010111000011;
    rom[21415] = 25'b0000000101100010000111001;
    rom[21416] = 25'b0000000101100001010101111;
    rom[21417] = 25'b0000000101100000100100101;
    rom[21418] = 25'b0000000101011111110011001;
    rom[21419] = 25'b0000000101011111000001110;
    rom[21420] = 25'b0000000101011110010000010;
    rom[21421] = 25'b0000000101011101011110110;
    rom[21422] = 25'b0000000101011100101101010;
    rom[21423] = 25'b0000000101011011111011100;
    rom[21424] = 25'b0000000101011011001001111;
    rom[21425] = 25'b0000000101011010011000001;
    rom[21426] = 25'b0000000101011001100110010;
    rom[21427] = 25'b0000000101011000110100011;
    rom[21428] = 25'b0000000101011000000010100;
    rom[21429] = 25'b0000000101010111010000101;
    rom[21430] = 25'b0000000101010110011110101;
    rom[21431] = 25'b0000000101010101101100100;
    rom[21432] = 25'b0000000101010100111010011;
    rom[21433] = 25'b0000000101010100001000001;
    rom[21434] = 25'b0000000101010011010110000;
    rom[21435] = 25'b0000000101010010100011101;
    rom[21436] = 25'b0000000101010001110001011;
    rom[21437] = 25'b0000000101010000111111000;
    rom[21438] = 25'b0000000101010000001100101;
    rom[21439] = 25'b0000000101001111011010001;
    rom[21440] = 25'b0000000101001110100111100;
    rom[21441] = 25'b0000000101001101110100111;
    rom[21442] = 25'b0000000101001101000010010;
    rom[21443] = 25'b0000000101001100001111101;
    rom[21444] = 25'b0000000101001011011100110;
    rom[21445] = 25'b0000000101001010101010000;
    rom[21446] = 25'b0000000101001001110111001;
    rom[21447] = 25'b0000000101001001000100010;
    rom[21448] = 25'b0000000101001000010001010;
    rom[21449] = 25'b0000000101000111011110010;
    rom[21450] = 25'b0000000101000110101011001;
    rom[21451] = 25'b0000000101000101111000000;
    rom[21452] = 25'b0000000101000101000100111;
    rom[21453] = 25'b0000000101000100010001101;
    rom[21454] = 25'b0000000101000011011110011;
    rom[21455] = 25'b0000000101000010101011000;
    rom[21456] = 25'b0000000101000001110111101;
    rom[21457] = 25'b0000000101000001000100001;
    rom[21458] = 25'b0000000101000000010000110;
    rom[21459] = 25'b0000000100111111011101001;
    rom[21460] = 25'b0000000100111110101001100;
    rom[21461] = 25'b0000000100111101110101111;
    rom[21462] = 25'b0000000100111101000010001;
    rom[21463] = 25'b0000000100111100001110011;
    rom[21464] = 25'b0000000100111011011010101;
    rom[21465] = 25'b0000000100111010100110110;
    rom[21466] = 25'b0000000100111001110010111;
    rom[21467] = 25'b0000000100111000111110111;
    rom[21468] = 25'b0000000100111000001010111;
    rom[21469] = 25'b0000000100110111010110110;
    rom[21470] = 25'b0000000100110110100010101;
    rom[21471] = 25'b0000000100110101101110100;
    rom[21472] = 25'b0000000100110100111010011;
    rom[21473] = 25'b0000000100110100000110000;
    rom[21474] = 25'b0000000100110011010001110;
    rom[21475] = 25'b0000000100110010011101011;
    rom[21476] = 25'b0000000100110001101000111;
    rom[21477] = 25'b0000000100110000110100011;
    rom[21478] = 25'b0000000100101111111111111;
    rom[21479] = 25'b0000000100101111001011011;
    rom[21480] = 25'b0000000100101110010110101;
    rom[21481] = 25'b0000000100101101100010000;
    rom[21482] = 25'b0000000100101100101101011;
    rom[21483] = 25'b0000000100101011111000100;
    rom[21484] = 25'b0000000100101011000011110;
    rom[21485] = 25'b0000000100101010001110110;
    rom[21486] = 25'b0000000100101001011001110;
    rom[21487] = 25'b0000000100101000100100111;
    rom[21488] = 25'b0000000100100111101111110;
    rom[21489] = 25'b0000000100100110111010110;
    rom[21490] = 25'b0000000100100110000101101;
    rom[21491] = 25'b0000000100100101010000011;
    rom[21492] = 25'b0000000100100100011011001;
    rom[21493] = 25'b0000000100100011100101111;
    rom[21494] = 25'b0000000100100010110000100;
    rom[21495] = 25'b0000000100100001111011001;
    rom[21496] = 25'b0000000100100001000101101;
    rom[21497] = 25'b0000000100100000010000001;
    rom[21498] = 25'b0000000100011111011010101;
    rom[21499] = 25'b0000000100011110100101000;
    rom[21500] = 25'b0000000100011101101111100;
    rom[21501] = 25'b0000000100011100111001110;
    rom[21502] = 25'b0000000100011100000100000;
    rom[21503] = 25'b0000000100011011001110001;
    rom[21504] = 25'b0000000100011010011000011;
    rom[21505] = 25'b0000000100011001100010011;
    rom[21506] = 25'b0000000100011000101100100;
    rom[21507] = 25'b0000000100010111110110100;
    rom[21508] = 25'b0000000100010111000000100;
    rom[21509] = 25'b0000000100010110001010011;
    rom[21510] = 25'b0000000100010101010100010;
    rom[21511] = 25'b0000000100010100011110001;
    rom[21512] = 25'b0000000100010011100111110;
    rom[21513] = 25'b0000000100010010110001100;
    rom[21514] = 25'b0000000100010001111011010;
    rom[21515] = 25'b0000000100010001000100110;
    rom[21516] = 25'b0000000100010000001110011;
    rom[21517] = 25'b0000000100001111010111111;
    rom[21518] = 25'b0000000100001110100001011;
    rom[21519] = 25'b0000000100001101101010110;
    rom[21520] = 25'b0000000100001100110100001;
    rom[21521] = 25'b0000000100001011111101011;
    rom[21522] = 25'b0000000100001011000110101;
    rom[21523] = 25'b0000000100001010001111111;
    rom[21524] = 25'b0000000100001001011001001;
    rom[21525] = 25'b0000000100001000100010001;
    rom[21526] = 25'b0000000100000111101011010;
    rom[21527] = 25'b0000000100000110110100010;
    rom[21528] = 25'b0000000100000101111101010;
    rom[21529] = 25'b0000000100000101000110001;
    rom[21530] = 25'b0000000100000100001111000;
    rom[21531] = 25'b0000000100000011010111111;
    rom[21532] = 25'b0000000100000010100000101;
    rom[21533] = 25'b0000000100000001101001011;
    rom[21534] = 25'b0000000100000000110010000;
    rom[21535] = 25'b0000000011111111111010101;
    rom[21536] = 25'b0000000011111111000011010;
    rom[21537] = 25'b0000000011111110001011110;
    rom[21538] = 25'b0000000011111101010100010;
    rom[21539] = 25'b0000000011111100011100110;
    rom[21540] = 25'b0000000011111011100101001;
    rom[21541] = 25'b0000000011111010101101011;
    rom[21542] = 25'b0000000011111001110101110;
    rom[21543] = 25'b0000000011111000111110000;
    rom[21544] = 25'b0000000011111000000110001;
    rom[21545] = 25'b0000000011110111001110011;
    rom[21546] = 25'b0000000011110110010110100;
    rom[21547] = 25'b0000000011110101011110100;
    rom[21548] = 25'b0000000011110100100110100;
    rom[21549] = 25'b0000000011110011101110100;
    rom[21550] = 25'b0000000011110010110110011;
    rom[21551] = 25'b0000000011110001111110010;
    rom[21552] = 25'b0000000011110001000110001;
    rom[21553] = 25'b0000000011110000001101111;
    rom[21554] = 25'b0000000011101111010101100;
    rom[21555] = 25'b0000000011101110011101010;
    rom[21556] = 25'b0000000011101101100100111;
    rom[21557] = 25'b0000000011101100101100011;
    rom[21558] = 25'b0000000011101011110100000;
    rom[21559] = 25'b0000000011101010111011011;
    rom[21560] = 25'b0000000011101010000010111;
    rom[21561] = 25'b0000000011101001001010011;
    rom[21562] = 25'b0000000011101000010001101;
    rom[21563] = 25'b0000000011100111011001000;
    rom[21564] = 25'b0000000011100110100000010;
    rom[21565] = 25'b0000000011100101100111011;
    rom[21566] = 25'b0000000011100100101110100;
    rom[21567] = 25'b0000000011100011110101101;
    rom[21568] = 25'b0000000011100010111100110;
    rom[21569] = 25'b0000000011100010000011111;
    rom[21570] = 25'b0000000011100001001010110;
    rom[21571] = 25'b0000000011100000010001110;
    rom[21572] = 25'b0000000011011111011000100;
    rom[21573] = 25'b0000000011011110011111011;
    rom[21574] = 25'b0000000011011101100110001;
    rom[21575] = 25'b0000000011011100101100111;
    rom[21576] = 25'b0000000011011011110011101;
    rom[21577] = 25'b0000000011011010111010011;
    rom[21578] = 25'b0000000011011010000000111;
    rom[21579] = 25'b0000000011011001000111100;
    rom[21580] = 25'b0000000011011000001101111;
    rom[21581] = 25'b0000000011010111010100011;
    rom[21582] = 25'b0000000011010110011010111;
    rom[21583] = 25'b0000000011010101100001010;
    rom[21584] = 25'b0000000011010100100111100;
    rom[21585] = 25'b0000000011010011101101111;
    rom[21586] = 25'b0000000011010010110100001;
    rom[21587] = 25'b0000000011010001111010011;
    rom[21588] = 25'b0000000011010001000000011;
    rom[21589] = 25'b0000000011010000000110100;
    rom[21590] = 25'b0000000011001111001100101;
    rom[21591] = 25'b0000000011001110010010101;
    rom[21592] = 25'b0000000011001101011000100;
    rom[21593] = 25'b0000000011001100011110100;
    rom[21594] = 25'b0000000011001011100100011;
    rom[21595] = 25'b0000000011001010101010001;
    rom[21596] = 25'b0000000011001001110000000;
    rom[21597] = 25'b0000000011001000110101110;
    rom[21598] = 25'b0000000011000111111011100;
    rom[21599] = 25'b0000000011000111000001001;
    rom[21600] = 25'b0000000011000110000110110;
    rom[21601] = 25'b0000000011000101001100010;
    rom[21602] = 25'b0000000011000100010001110;
    rom[21603] = 25'b0000000011000011010111010;
    rom[21604] = 25'b0000000011000010011100110;
    rom[21605] = 25'b0000000011000001100010000;
    rom[21606] = 25'b0000000011000000100111011;
    rom[21607] = 25'b0000000010111111101100110;
    rom[21608] = 25'b0000000010111110110010000;
    rom[21609] = 25'b0000000010111101110111001;
    rom[21610] = 25'b0000000010111100111100011;
    rom[21611] = 25'b0000000010111100000001100;
    rom[21612] = 25'b0000000010111011000110101;
    rom[21613] = 25'b0000000010111010001011100;
    rom[21614] = 25'b0000000010111001010000100;
    rom[21615] = 25'b0000000010111000010101100;
    rom[21616] = 25'b0000000010110111011010011;
    rom[21617] = 25'b0000000010110110011111010;
    rom[21618] = 25'b0000000010110101100100001;
    rom[21619] = 25'b0000000010110100101000111;
    rom[21620] = 25'b0000000010110011101101101;
    rom[21621] = 25'b0000000010110010110010010;
    rom[21622] = 25'b0000000010110001110111000;
    rom[21623] = 25'b0000000010110000111011101;
    rom[21624] = 25'b0000000010110000000000001;
    rom[21625] = 25'b0000000010101111000100101;
    rom[21626] = 25'b0000000010101110001001001;
    rom[21627] = 25'b0000000010101101001101100;
    rom[21628] = 25'b0000000010101100010001111;
    rom[21629] = 25'b0000000010101011010110010;
    rom[21630] = 25'b0000000010101010011010100;
    rom[21631] = 25'b0000000010101001011110110;
    rom[21632] = 25'b0000000010101000100011000;
    rom[21633] = 25'b0000000010100111100111010;
    rom[21634] = 25'b0000000010100110101011010;
    rom[21635] = 25'b0000000010100101101111011;
    rom[21636] = 25'b0000000010100100110011100;
    rom[21637] = 25'b0000000010100011110111011;
    rom[21638] = 25'b0000000010100010111011011;
    rom[21639] = 25'b0000000010100001111111010;
    rom[21640] = 25'b0000000010100001000011001;
    rom[21641] = 25'b0000000010100000000111000;
    rom[21642] = 25'b0000000010011111001010110;
    rom[21643] = 25'b0000000010011110001110100;
    rom[21644] = 25'b0000000010011101010010010;
    rom[21645] = 25'b0000000010011100010101111;
    rom[21646] = 25'b0000000010011011011001100;
    rom[21647] = 25'b0000000010011010011101001;
    rom[21648] = 25'b0000000010011001100000101;
    rom[21649] = 25'b0000000010011000100100001;
    rom[21650] = 25'b0000000010010111100111101;
    rom[21651] = 25'b0000000010010110101011000;
    rom[21652] = 25'b0000000010010101101110011;
    rom[21653] = 25'b0000000010010100110001101;
    rom[21654] = 25'b0000000010010011110101000;
    rom[21655] = 25'b0000000010010010111000010;
    rom[21656] = 25'b0000000010010001111011100;
    rom[21657] = 25'b0000000010010000111110101;
    rom[21658] = 25'b0000000010010000000001110;
    rom[21659] = 25'b0000000010001111000100111;
    rom[21660] = 25'b0000000010001110000111111;
    rom[21661] = 25'b0000000010001101001010111;
    rom[21662] = 25'b0000000010001100001101111;
    rom[21663] = 25'b0000000010001011010000110;
    rom[21664] = 25'b0000000010001010010011101;
    rom[21665] = 25'b0000000010001001010110100;
    rom[21666] = 25'b0000000010001000011001010;
    rom[21667] = 25'b0000000010000111011100000;
    rom[21668] = 25'b0000000010000110011110110;
    rom[21669] = 25'b0000000010000101100001011;
    rom[21670] = 25'b0000000010000100100100000;
    rom[21671] = 25'b0000000010000011100110110;
    rom[21672] = 25'b0000000010000010101001010;
    rom[21673] = 25'b0000000010000001101011110;
    rom[21674] = 25'b0000000010000000101110010;
    rom[21675] = 25'b0000000001111111110000101;
    rom[21676] = 25'b0000000001111110110011001;
    rom[21677] = 25'b0000000001111101110101100;
    rom[21678] = 25'b0000000001111100110111110;
    rom[21679] = 25'b0000000001111011111010000;
    rom[21680] = 25'b0000000001111010111100010;
    rom[21681] = 25'b0000000001111001111110100;
    rom[21682] = 25'b0000000001111001000000101;
    rom[21683] = 25'b0000000001111000000010110;
    rom[21684] = 25'b0000000001110111000100110;
    rom[21685] = 25'b0000000001110110000110111;
    rom[21686] = 25'b0000000001110101001000111;
    rom[21687] = 25'b0000000001110100001010111;
    rom[21688] = 25'b0000000001110011001100110;
    rom[21689] = 25'b0000000001110010001110101;
    rom[21690] = 25'b0000000001110001010000100;
    rom[21691] = 25'b0000000001110000010010011;
    rom[21692] = 25'b0000000001101111010100000;
    rom[21693] = 25'b0000000001101110010101110;
    rom[21694] = 25'b0000000001101101010111100;
    rom[21695] = 25'b0000000001101100011001010;
    rom[21696] = 25'b0000000001101011011010110;
    rom[21697] = 25'b0000000001101010011100011;
    rom[21698] = 25'b0000000001101001011101111;
    rom[21699] = 25'b0000000001101000011111011;
    rom[21700] = 25'b0000000001100111100000111;
    rom[21701] = 25'b0000000001100110100010010;
    rom[21702] = 25'b0000000001100101100011101;
    rom[21703] = 25'b0000000001100100100101000;
    rom[21704] = 25'b0000000001100011100110011;
    rom[21705] = 25'b0000000001100010100111101;
    rom[21706] = 25'b0000000001100001101000111;
    rom[21707] = 25'b0000000001100000101010000;
    rom[21708] = 25'b0000000001011111101011001;
    rom[21709] = 25'b0000000001011110101100010;
    rom[21710] = 25'b0000000001011101101101011;
    rom[21711] = 25'b0000000001011100101110011;
    rom[21712] = 25'b0000000001011011101111100;
    rom[21713] = 25'b0000000001011010110000011;
    rom[21714] = 25'b0000000001011001110001010;
    rom[21715] = 25'b0000000001011000110010010;
    rom[21716] = 25'b0000000001010111110011001;
    rom[21717] = 25'b0000000001010110110011111;
    rom[21718] = 25'b0000000001010101110100101;
    rom[21719] = 25'b0000000001010100110101100;
    rom[21720] = 25'b0000000001010011110110001;
    rom[21721] = 25'b0000000001010010110110111;
    rom[21722] = 25'b0000000001010001110111100;
    rom[21723] = 25'b0000000001010000111000001;
    rom[21724] = 25'b0000000001001111111000110;
    rom[21725] = 25'b0000000001001110111001001;
    rom[21726] = 25'b0000000001001101111001101;
    rom[21727] = 25'b0000000001001100111010001;
    rom[21728] = 25'b0000000001001011111010101;
    rom[21729] = 25'b0000000001001010111010111;
    rom[21730] = 25'b0000000001001001111011010;
    rom[21731] = 25'b0000000001001000111011101;
    rom[21732] = 25'b0000000001000111111011111;
    rom[21733] = 25'b0000000001000110111100001;
    rom[21734] = 25'b0000000001000101111100011;
    rom[21735] = 25'b0000000001000100111100100;
    rom[21736] = 25'b0000000001000011111100101;
    rom[21737] = 25'b0000000001000010111100110;
    rom[21738] = 25'b0000000001000001111100110;
    rom[21739] = 25'b0000000001000000111100110;
    rom[21740] = 25'b0000000000111111111100110;
    rom[21741] = 25'b0000000000111110111100110;
    rom[21742] = 25'b0000000000111101111100101;
    rom[21743] = 25'b0000000000111100111100100;
    rom[21744] = 25'b0000000000111011111100011;
    rom[21745] = 25'b0000000000111010111100010;
    rom[21746] = 25'b0000000000111001111100000;
    rom[21747] = 25'b0000000000111000111011110;
    rom[21748] = 25'b0000000000110111111011100;
    rom[21749] = 25'b0000000000110110111011001;
    rom[21750] = 25'b0000000000110101111010110;
    rom[21751] = 25'b0000000000110100111010011;
    rom[21752] = 25'b0000000000110011111001111;
    rom[21753] = 25'b0000000000110010111001100;
    rom[21754] = 25'b0000000000110001111000111;
    rom[21755] = 25'b0000000000110000111000011;
    rom[21756] = 25'b0000000000101111110111111;
    rom[21757] = 25'b0000000000101110110111010;
    rom[21758] = 25'b0000000000101101110110101;
    rom[21759] = 25'b0000000000101100110110000;
    rom[21760] = 25'b0000000000101011110101010;
    rom[21761] = 25'b0000000000101010110100101;
    rom[21762] = 25'b0000000000101001110011110;
    rom[21763] = 25'b0000000000101000110011000;
    rom[21764] = 25'b0000000000100111110010001;
    rom[21765] = 25'b0000000000100110110001010;
    rom[21766] = 25'b0000000000100101110000011;
    rom[21767] = 25'b0000000000100100101111011;
    rom[21768] = 25'b0000000000100011101110011;
    rom[21769] = 25'b0000000000100010101101011;
    rom[21770] = 25'b0000000000100001101100011;
    rom[21771] = 25'b0000000000100000101011011;
    rom[21772] = 25'b0000000000011111101010010;
    rom[21773] = 25'b0000000000011110101001001;
    rom[21774] = 25'b0000000000011101100111111;
    rom[21775] = 25'b0000000000011100100110110;
    rom[21776] = 25'b0000000000011011100101100;
    rom[21777] = 25'b0000000000011010100100010;
    rom[21778] = 25'b0000000000011001100010111;
    rom[21779] = 25'b0000000000011000100001101;
    rom[21780] = 25'b0000000000010111100000010;
    rom[21781] = 25'b0000000000010110011110111;
    rom[21782] = 25'b0000000000010101011101011;
    rom[21783] = 25'b0000000000010100011011111;
    rom[21784] = 25'b0000000000010011011010100;
    rom[21785] = 25'b0000000000010010011000111;
    rom[21786] = 25'b0000000000010001010111011;
    rom[21787] = 25'b0000000000010000010101110;
    rom[21788] = 25'b0000000000001111010100001;
    rom[21789] = 25'b0000000000001110010010100;
    rom[21790] = 25'b0000000000001101010000110;
    rom[21791] = 25'b0000000000001100001111001;
    rom[21792] = 25'b0000000000001011001101011;
    rom[21793] = 25'b0000000000001010001011100;
    rom[21794] = 25'b0000000000001001001001110;
    rom[21795] = 25'b0000000000001000000111111;
    rom[21796] = 25'b0000000000000111000110000;
    rom[21797] = 25'b0000000000000110000100000;
    rom[21798] = 25'b0000000000000101000010001;
    rom[21799] = 25'b0000000000000100000000010;
    rom[21800] = 25'b0000000000000010111110001;
    rom[21801] = 25'b0000000000000001111100001;
    rom[21802] = 25'b0000000000000000111010001;
    rom[21803] = 25'b1111111111111111111000001;
    rom[21804] = 25'b1111111111111110110110000;
    rom[21805] = 25'b1111111111111101110011111;
    rom[21806] = 25'b1111111111111100110001101;
    rom[21807] = 25'b1111111111111011101111011;
    rom[21808] = 25'b1111111111111010101101010;
    rom[21809] = 25'b1111111111111001101010111;
    rom[21810] = 25'b1111111111111000101000101;
    rom[21811] = 25'b1111111111110111100110010;
    rom[21812] = 25'b1111111111110110100011111;
    rom[21813] = 25'b1111111111110101100001100;
    rom[21814] = 25'b1111111111110100011111001;
    rom[21815] = 25'b1111111111110011011100101;
    rom[21816] = 25'b1111111111110010011010001;
    rom[21817] = 25'b1111111111110001010111101;
    rom[21818] = 25'b1111111111110000010101000;
    rom[21819] = 25'b1111111111101111010010101;
    rom[21820] = 25'b1111111111101110001111111;
    rom[21821] = 25'b1111111111101101001101010;
    rom[21822] = 25'b1111111111101100001010101;
    rom[21823] = 25'b1111111111101011001000000;
    rom[21824] = 25'b1111111111101010000101010;
    rom[21825] = 25'b1111111111101001000010100;
    rom[21826] = 25'b1111111111100111111111110;
    rom[21827] = 25'b1111111111100110111100111;
    rom[21828] = 25'b1111111111100101111010001;
    rom[21829] = 25'b1111111111100100110111010;
    rom[21830] = 25'b1111111111100011110100010;
    rom[21831] = 25'b1111111111100010110001011;
    rom[21832] = 25'b1111111111100001101110011;
    rom[21833] = 25'b1111111111100000101011100;
    rom[21834] = 25'b1111111111011111101000011;
    rom[21835] = 25'b1111111111011110100101011;
    rom[21836] = 25'b1111111111011101100010011;
    rom[21837] = 25'b1111111111011100011111010;
    rom[21838] = 25'b1111111111011011011100001;
    rom[21839] = 25'b1111111111011010011001000;
    rom[21840] = 25'b1111111111011001010101111;
    rom[21841] = 25'b1111111111011000010010101;
    rom[21842] = 25'b1111111111010111001111011;
    rom[21843] = 25'b1111111111010110001100001;
    rom[21844] = 25'b1111111111010101001000111;
    rom[21845] = 25'b1111111111010100000101100;
    rom[21846] = 25'b1111111111010011000010010;
    rom[21847] = 25'b1111111111010001111110111;
    rom[21848] = 25'b1111111111010000111011100;
    rom[21849] = 25'b1111111111001111111000000;
    rom[21850] = 25'b1111111111001110110100101;
    rom[21851] = 25'b1111111111001101110001001;
    rom[21852] = 25'b1111111111001100101101101;
    rom[21853] = 25'b1111111111001011101010000;
    rom[21854] = 25'b1111111111001010100110100;
    rom[21855] = 25'b1111111111001001100010111;
    rom[21856] = 25'b1111111111001000011111010;
    rom[21857] = 25'b1111111111000111011011110;
    rom[21858] = 25'b1111111111000110011000001;
    rom[21859] = 25'b1111111111000101010100011;
    rom[21860] = 25'b1111111111000100010000101;
    rom[21861] = 25'b1111111111000011001100111;
    rom[21862] = 25'b1111111111000010001001001;
    rom[21863] = 25'b1111111111000001000101011;
    rom[21864] = 25'b1111111111000000000001101;
    rom[21865] = 25'b1111111110111110111101101;
    rom[21866] = 25'b1111111110111101111001110;
    rom[21867] = 25'b1111111110111100110101111;
    rom[21868] = 25'b1111111110111011110010000;
    rom[21869] = 25'b1111111110111010101110001;
    rom[21870] = 25'b1111111110111001101010001;
    rom[21871] = 25'b1111111110111000100110001;
    rom[21872] = 25'b1111111110110111100010000;
    rom[21873] = 25'b1111111110110110011110001;
    rom[21874] = 25'b1111111110110101011010000;
    rom[21875] = 25'b1111111110110100010101111;
    rom[21876] = 25'b1111111110110011010001110;
    rom[21877] = 25'b1111111110110010001101101;
    rom[21878] = 25'b1111111110110001001001011;
    rom[21879] = 25'b1111111110110000000101010;
    rom[21880] = 25'b1111111110101111000001000;
    rom[21881] = 25'b1111111110101101111100110;
    rom[21882] = 25'b1111111110101100111000100;
    rom[21883] = 25'b1111111110101011110100010;
    rom[21884] = 25'b1111111110101010101111111;
    rom[21885] = 25'b1111111110101001101011100;
    rom[21886] = 25'b1111111110101000100111001;
    rom[21887] = 25'b1111111110100111100010111;
    rom[21888] = 25'b1111111110100110011110011;
    rom[21889] = 25'b1111111110100101011010000;
    rom[21890] = 25'b1111111110100100010101100;
    rom[21891] = 25'b1111111110100011010001000;
    rom[21892] = 25'b1111111110100010001100100;
    rom[21893] = 25'b1111111110100001001000000;
    rom[21894] = 25'b1111111110100000000011100;
    rom[21895] = 25'b1111111110011110111110111;
    rom[21896] = 25'b1111111110011101111010010;
    rom[21897] = 25'b1111111110011100110101101;
    rom[21898] = 25'b1111111110011011110001000;
    rom[21899] = 25'b1111111110011010101100010;
    rom[21900] = 25'b1111111110011001100111101;
    rom[21901] = 25'b1111111110011000100010111;
    rom[21902] = 25'b1111111110010111011110001;
    rom[21903] = 25'b1111111110010110011001011;
    rom[21904] = 25'b1111111110010101010100101;
    rom[21905] = 25'b1111111110010100001111110;
    rom[21906] = 25'b1111111110010011001011000;
    rom[21907] = 25'b1111111110010010000110001;
    rom[21908] = 25'b1111111110010001000001010;
    rom[21909] = 25'b1111111110001111111100011;
    rom[21910] = 25'b1111111110001110110111100;
    rom[21911] = 25'b1111111110001101110010100;
    rom[21912] = 25'b1111111110001100101101100;
    rom[21913] = 25'b1111111110001011101000100;
    rom[21914] = 25'b1111111110001010100011101;
    rom[21915] = 25'b1111111110001001011110100;
    rom[21916] = 25'b1111111110001000011001100;
    rom[21917] = 25'b1111111110000111010100011;
    rom[21918] = 25'b1111111110000110001111011;
    rom[21919] = 25'b1111111110000101001010010;
    rom[21920] = 25'b1111111110000100000101000;
    rom[21921] = 25'b1111111110000011000000000;
    rom[21922] = 25'b1111111110000001111010110;
    rom[21923] = 25'b1111111110000000110101100;
    rom[21924] = 25'b1111111101111111110000011;
    rom[21925] = 25'b1111111101111110101011000;
    rom[21926] = 25'b1111111101111101100101111;
    rom[21927] = 25'b1111111101111100100000100;
    rom[21928] = 25'b1111111101111011011011010;
    rom[21929] = 25'b1111111101111010010110000;
    rom[21930] = 25'b1111111101111001010000101;
    rom[21931] = 25'b1111111101111000001011010;
    rom[21932] = 25'b1111111101110111000101110;
    rom[21933] = 25'b1111111101110110000000011;
    rom[21934] = 25'b1111111101110100111011000;
    rom[21935] = 25'b1111111101110011110101100;
    rom[21936] = 25'b1111111101110010110000001;
    rom[21937] = 25'b1111111101110001101010110;
    rom[21938] = 25'b1111111101110000100101001;
    rom[21939] = 25'b1111111101101111011111101;
    rom[21940] = 25'b1111111101101110011010000;
    rom[21941] = 25'b1111111101101101010100100;
    rom[21942] = 25'b1111111101101100001110111;
    rom[21943] = 25'b1111111101101011001001011;
    rom[21944] = 25'b1111111101101010000011110;
    rom[21945] = 25'b1111111101101000111110001;
    rom[21946] = 25'b1111111101100111111000011;
    rom[21947] = 25'b1111111101100110110010110;
    rom[21948] = 25'b1111111101100101101101001;
    rom[21949] = 25'b1111111101100100100111011;
    rom[21950] = 25'b1111111101100011100001101;
    rom[21951] = 25'b1111111101100010011011111;
    rom[21952] = 25'b1111111101100001010110001;
    rom[21953] = 25'b1111111101100000010000011;
    rom[21954] = 25'b1111111101011111001010100;
    rom[21955] = 25'b1111111101011110000100101;
    rom[21956] = 25'b1111111101011100111110111;
    rom[21957] = 25'b1111111101011011111001001;
    rom[21958] = 25'b1111111101011010110011001;
    rom[21959] = 25'b1111111101011001101101010;
    rom[21960] = 25'b1111111101011000100111011;
    rom[21961] = 25'b1111111101010111100001100;
    rom[21962] = 25'b1111111101010110011011100;
    rom[21963] = 25'b1111111101010101010101100;
    rom[21964] = 25'b1111111101010100001111100;
    rom[21965] = 25'b1111111101010011001001101;
    rom[21966] = 25'b1111111101010010000011100;
    rom[21967] = 25'b1111111101010000111101100;
    rom[21968] = 25'b1111111101001111110111100;
    rom[21969] = 25'b1111111101001110110001011;
    rom[21970] = 25'b1111111101001101101011010;
    rom[21971] = 25'b1111111101001100100101001;
    rom[21972] = 25'b1111111101001011011111001;
    rom[21973] = 25'b1111111101001010011001000;
    rom[21974] = 25'b1111111101001001010010111;
    rom[21975] = 25'b1111111101001000001100101;
    rom[21976] = 25'b1111111101000111000110100;
    rom[21977] = 25'b1111111101000110000000010;
    rom[21978] = 25'b1111111101000100111010000;
    rom[21979] = 25'b1111111101000011110011111;
    rom[21980] = 25'b1111111101000010101101101;
    rom[21981] = 25'b1111111101000001100111011;
    rom[21982] = 25'b1111111101000000100001000;
    rom[21983] = 25'b1111111100111111011010110;
    rom[21984] = 25'b1111111100111110010100011;
    rom[21985] = 25'b1111111100111101001110001;
    rom[21986] = 25'b1111111100111100000111110;
    rom[21987] = 25'b1111111100111011000001011;
    rom[21988] = 25'b1111111100111001111011000;
    rom[21989] = 25'b1111111100111000110100110;
    rom[21990] = 25'b1111111100110111101110010;
    rom[21991] = 25'b1111111100110110100111111;
    rom[21992] = 25'b1111111100110101100001100;
    rom[21993] = 25'b1111111100110100011011000;
    rom[21994] = 25'b1111111100110011010100100;
    rom[21995] = 25'b1111111100110010001110000;
    rom[21996] = 25'b1111111100110001000111100;
    rom[21997] = 25'b1111111100110000000001000;
    rom[21998] = 25'b1111111100101110111010100;
    rom[21999] = 25'b1111111100101101110100000;
    rom[22000] = 25'b1111111100101100101101100;
    rom[22001] = 25'b1111111100101011100110111;
    rom[22002] = 25'b1111111100101010100000010;
    rom[22003] = 25'b1111111100101001011001110;
    rom[22004] = 25'b1111111100101000010011001;
    rom[22005] = 25'b1111111100100111001100100;
    rom[22006] = 25'b1111111100100110000101111;
    rom[22007] = 25'b1111111100100100111111010;
    rom[22008] = 25'b1111111100100011111000101;
    rom[22009] = 25'b1111111100100010110001111;
    rom[22010] = 25'b1111111100100001101011010;
    rom[22011] = 25'b1111111100100000100100100;
    rom[22012] = 25'b1111111100011111011101111;
    rom[22013] = 25'b1111111100011110010111001;
    rom[22014] = 25'b1111111100011101010000011;
    rom[22015] = 25'b1111111100011100001001101;
    rom[22016] = 25'b1111111100011011000010111;
    rom[22017] = 25'b1111111100011001111100001;
    rom[22018] = 25'b1111111100011000110101010;
    rom[22019] = 25'b1111111100010111101110100;
    rom[22020] = 25'b1111111100010110100111110;
    rom[22021] = 25'b1111111100010101100000111;
    rom[22022] = 25'b1111111100010100011010000;
    rom[22023] = 25'b1111111100010011010011010;
    rom[22024] = 25'b1111111100010010001100011;
    rom[22025] = 25'b1111111100010001000101100;
    rom[22026] = 25'b1111111100001111111110101;
    rom[22027] = 25'b1111111100001110110111110;
    rom[22028] = 25'b1111111100001101110000111;
    rom[22029] = 25'b1111111100001100101001111;
    rom[22030] = 25'b1111111100001011100011000;
    rom[22031] = 25'b1111111100001010011100000;
    rom[22032] = 25'b1111111100001001010101000;
    rom[22033] = 25'b1111111100001000001110001;
    rom[22034] = 25'b1111111100000111000111001;
    rom[22035] = 25'b1111111100000110000000001;
    rom[22036] = 25'b1111111100000100111001001;
    rom[22037] = 25'b1111111100000011110010001;
    rom[22038] = 25'b1111111100000010101011001;
    rom[22039] = 25'b1111111100000001100100001;
    rom[22040] = 25'b1111111100000000011101001;
    rom[22041] = 25'b1111111011111111010110000;
    rom[22042] = 25'b1111111011111110001110111;
    rom[22043] = 25'b1111111011111101000111111;
    rom[22044] = 25'b1111111011111100000000110;
    rom[22045] = 25'b1111111011111010111001110;
    rom[22046] = 25'b1111111011111001110010101;
    rom[22047] = 25'b1111111011111000101011100;
    rom[22048] = 25'b1111111011110111100100011;
    rom[22049] = 25'b1111111011110110011101010;
    rom[22050] = 25'b1111111011110101010110010;
    rom[22051] = 25'b1111111011110100001111000;
    rom[22052] = 25'b1111111011110011000111111;
    rom[22053] = 25'b1111111011110010000000110;
    rom[22054] = 25'b1111111011110000111001101;
    rom[22055] = 25'b1111111011101111110010010;
    rom[22056] = 25'b1111111011101110101011001;
    rom[22057] = 25'b1111111011101101100100000;
    rom[22058] = 25'b1111111011101100011100110;
    rom[22059] = 25'b1111111011101011010101101;
    rom[22060] = 25'b1111111011101010001110011;
    rom[22061] = 25'b1111111011101001000111001;
    rom[22062] = 25'b1111111011100111111111110;
    rom[22063] = 25'b1111111011100110111000100;
    rom[22064] = 25'b1111111011100101110001010;
    rom[22065] = 25'b1111111011100100101010000;
    rom[22066] = 25'b1111111011100011100010110;
    rom[22067] = 25'b1111111011100010011011100;
    rom[22068] = 25'b1111111011100001010100010;
    rom[22069] = 25'b1111111011100000001100111;
    rom[22070] = 25'b1111111011011111000101101;
    rom[22071] = 25'b1111111011011101111110010;
    rom[22072] = 25'b1111111011011100110111000;
    rom[22073] = 25'b1111111011011011101111101;
    rom[22074] = 25'b1111111011011010101000010;
    rom[22075] = 25'b1111111011011001100001000;
    rom[22076] = 25'b1111111011011000011001101;
    rom[22077] = 25'b1111111011010111010010010;
    rom[22078] = 25'b1111111011010110001010111;
    rom[22079] = 25'b1111111011010101000011100;
    rom[22080] = 25'b1111111011010011111100001;
    rom[22081] = 25'b1111111011010010110100110;
    rom[22082] = 25'b1111111011010001101101011;
    rom[22083] = 25'b1111111011010000100110000;
    rom[22084] = 25'b1111111011001111011110100;
    rom[22085] = 25'b1111111011001110010111001;
    rom[22086] = 25'b1111111011001101001111110;
    rom[22087] = 25'b1111111011001100001000010;
    rom[22088] = 25'b1111111011001011000000111;
    rom[22089] = 25'b1111111011001001111001011;
    rom[22090] = 25'b1111111011001000110010000;
    rom[22091] = 25'b1111111011000111101010100;
    rom[22092] = 25'b1111111011000110100011001;
    rom[22093] = 25'b1111111011000101011011101;
    rom[22094] = 25'b1111111011000100010100010;
    rom[22095] = 25'b1111111011000011001100101;
    rom[22096] = 25'b1111111011000010000101010;
    rom[22097] = 25'b1111111011000000111101110;
    rom[22098] = 25'b1111111010111111110110010;
    rom[22099] = 25'b1111111010111110101110111;
    rom[22100] = 25'b1111111010111101100111010;
    rom[22101] = 25'b1111111010111100011111111;
    rom[22102] = 25'b1111111010111011011000011;
    rom[22103] = 25'b1111111010111010010000110;
    rom[22104] = 25'b1111111010111001001001011;
    rom[22105] = 25'b1111111010111000000001110;
    rom[22106] = 25'b1111111010110110111010010;
    rom[22107] = 25'b1111111010110101110010110;
    rom[22108] = 25'b1111111010110100101011010;
    rom[22109] = 25'b1111111010110011100011101;
    rom[22110] = 25'b1111111010110010011100001;
    rom[22111] = 25'b1111111010110001010100101;
    rom[22112] = 25'b1111111010110000001101001;
    rom[22113] = 25'b1111111010101111000101100;
    rom[22114] = 25'b1111111010101101111110000;
    rom[22115] = 25'b1111111010101100110110100;
    rom[22116] = 25'b1111111010101011101110111;
    rom[22117] = 25'b1111111010101010100111010;
    rom[22118] = 25'b1111111010101001011111110;
    rom[22119] = 25'b1111111010101000011000010;
    rom[22120] = 25'b1111111010100111010000101;
    rom[22121] = 25'b1111111010100110001001001;
    rom[22122] = 25'b1111111010100101000001100;
    rom[22123] = 25'b1111111010100011111001111;
    rom[22124] = 25'b1111111010100010110010011;
    rom[22125] = 25'b1111111010100001101010110;
    rom[22126] = 25'b1111111010100000100011010;
    rom[22127] = 25'b1111111010011111011011101;
    rom[22128] = 25'b1111111010011110010100000;
    rom[22129] = 25'b1111111010011101001100011;
    rom[22130] = 25'b1111111010011100000100110;
    rom[22131] = 25'b1111111010011010111101010;
    rom[22132] = 25'b1111111010011001110101101;
    rom[22133] = 25'b1111111010011000101110001;
    rom[22134] = 25'b1111111010010111100110100;
    rom[22135] = 25'b1111111010010110011110111;
    rom[22136] = 25'b1111111010010101010111010;
    rom[22137] = 25'b1111111010010100001111101;
    rom[22138] = 25'b1111111010010011001000000;
    rom[22139] = 25'b1111111010010010000000011;
    rom[22140] = 25'b1111111010010000111000111;
    rom[22141] = 25'b1111111010001111110001010;
    rom[22142] = 25'b1111111010001110101001101;
    rom[22143] = 25'b1111111010001101100010000;
    rom[22144] = 25'b1111111010001100011010100;
    rom[22145] = 25'b1111111010001011010010111;
    rom[22146] = 25'b1111111010001010001011010;
    rom[22147] = 25'b1111111010001001000011101;
    rom[22148] = 25'b1111111010000111111100000;
    rom[22149] = 25'b1111111010000110110100011;
    rom[22150] = 25'b1111111010000101101100110;
    rom[22151] = 25'b1111111010000100100101001;
    rom[22152] = 25'b1111111010000011011101100;
    rom[22153] = 25'b1111111010000010010110000;
    rom[22154] = 25'b1111111010000001001110011;
    rom[22155] = 25'b1111111010000000000110110;
    rom[22156] = 25'b1111111001111110111111001;
    rom[22157] = 25'b1111111001111101110111101;
    rom[22158] = 25'b1111111001111100110000000;
    rom[22159] = 25'b1111111001111011101000011;
    rom[22160] = 25'b1111111001111010100000110;
    rom[22161] = 25'b1111111001111001011001001;
    rom[22162] = 25'b1111111001111000010001100;
    rom[22163] = 25'b1111111001110111001001111;
    rom[22164] = 25'b1111111001110110000010011;
    rom[22165] = 25'b1111111001110100111010110;
    rom[22166] = 25'b1111111001110011110011010;
    rom[22167] = 25'b1111111001110010101011101;
    rom[22168] = 25'b1111111001110001100100000;
    rom[22169] = 25'b1111111001110000011100011;
    rom[22170] = 25'b1111111001101111010100110;
    rom[22171] = 25'b1111111001101110001101010;
    rom[22172] = 25'b1111111001101101000101101;
    rom[22173] = 25'b1111111001101011111110001;
    rom[22174] = 25'b1111111001101010110110100;
    rom[22175] = 25'b1111111001101001101110111;
    rom[22176] = 25'b1111111001101000100111011;
    rom[22177] = 25'b1111111001100111011111110;
    rom[22178] = 25'b1111111001100110011000010;
    rom[22179] = 25'b1111111001100101010000110;
    rom[22180] = 25'b1111111001100100001001001;
    rom[22181] = 25'b1111111001100011000001100;
    rom[22182] = 25'b1111111001100001111010000;
    rom[22183] = 25'b1111111001100000110010100;
    rom[22184] = 25'b1111111001011111101011000;
    rom[22185] = 25'b1111111001011110100011011;
    rom[22186] = 25'b1111111001011101011011111;
    rom[22187] = 25'b1111111001011100010100011;
    rom[22188] = 25'b1111111001011011001100110;
    rom[22189] = 25'b1111111001011010000101010;
    rom[22190] = 25'b1111111001011000111101110;
    rom[22191] = 25'b1111111001010111110110010;
    rom[22192] = 25'b1111111001010110101110101;
    rom[22193] = 25'b1111111001010101100111010;
    rom[22194] = 25'b1111111001010100011111110;
    rom[22195] = 25'b1111111001010011011000001;
    rom[22196] = 25'b1111111001010010010000110;
    rom[22197] = 25'b1111111001010001001001001;
    rom[22198] = 25'b1111111001010000000001110;
    rom[22199] = 25'b1111111001001110111010010;
    rom[22200] = 25'b1111111001001101110010110;
    rom[22201] = 25'b1111111001001100101011011;
    rom[22202] = 25'b1111111001001011100011110;
    rom[22203] = 25'b1111111001001010011100011;
    rom[22204] = 25'b1111111001001001010100111;
    rom[22205] = 25'b1111111001001000001101100;
    rom[22206] = 25'b1111111001000111000110000;
    rom[22207] = 25'b1111111001000101111110101;
    rom[22208] = 25'b1111111001000100110111001;
    rom[22209] = 25'b1111111001000011101111110;
    rom[22210] = 25'b1111111001000010101000011;
    rom[22211] = 25'b1111111001000001100000111;
    rom[22212] = 25'b1111111001000000011001100;
    rom[22213] = 25'b1111111000111111010010001;
    rom[22214] = 25'b1111111000111110001010101;
    rom[22215] = 25'b1111111000111101000011011;
    rom[22216] = 25'b1111111000111011111011111;
    rom[22217] = 25'b1111111000111010110100100;
    rom[22218] = 25'b1111111000111001101101010;
    rom[22219] = 25'b1111111000111000100101111;
    rom[22220] = 25'b1111111000110111011110100;
    rom[22221] = 25'b1111111000110110010111001;
    rom[22222] = 25'b1111111000110101001111110;
    rom[22223] = 25'b1111111000110100001000100;
    rom[22224] = 25'b1111111000110011000001001;
    rom[22225] = 25'b1111111000110001111001111;
    rom[22226] = 25'b1111111000110000110010100;
    rom[22227] = 25'b1111111000101111101011010;
    rom[22228] = 25'b1111111000101110100011111;
    rom[22229] = 25'b1111111000101101011100101;
    rom[22230] = 25'b1111111000101100010101011;
    rom[22231] = 25'b1111111000101011001110001;
    rom[22232] = 25'b1111111000101010000110110;
    rom[22233] = 25'b1111111000101000111111100;
    rom[22234] = 25'b1111111000100111111000011;
    rom[22235] = 25'b1111111000100110110001001;
    rom[22236] = 25'b1111111000100101101001111;
    rom[22237] = 25'b1111111000100100100010110;
    rom[22238] = 25'b1111111000100011011011100;
    rom[22239] = 25'b1111111000100010010100010;
    rom[22240] = 25'b1111111000100001001101000;
    rom[22241] = 25'b1111111000100000000101111;
    rom[22242] = 25'b1111111000011110111110110;
    rom[22243] = 25'b1111111000011101110111100;
    rom[22244] = 25'b1111111000011100110000011;
    rom[22245] = 25'b1111111000011011101001010;
    rom[22246] = 25'b1111111000011010100010001;
    rom[22247] = 25'b1111111000011001011011000;
    rom[22248] = 25'b1111111000011000010100000;
    rom[22249] = 25'b1111111000010111001100110;
    rom[22250] = 25'b1111111000010110000101110;
    rom[22251] = 25'b1111111000010100111110101;
    rom[22252] = 25'b1111111000010011110111101;
    rom[22253] = 25'b1111111000010010110000100;
    rom[22254] = 25'b1111111000010001101001100;
    rom[22255] = 25'b1111111000010000100010011;
    rom[22256] = 25'b1111111000001111011011011;
    rom[22257] = 25'b1111111000001110010100011;
    rom[22258] = 25'b1111111000001101001101011;
    rom[22259] = 25'b1111111000001100000110011;
    rom[22260] = 25'b1111111000001010111111011;
    rom[22261] = 25'b1111111000001001111000011;
    rom[22262] = 25'b1111111000001000110001100;
    rom[22263] = 25'b1111111000000111101010100;
    rom[22264] = 25'b1111111000000110100011100;
    rom[22265] = 25'b1111111000000101011100101;
    rom[22266] = 25'b1111111000000100010101101;
    rom[22267] = 25'b1111111000000011001110110;
    rom[22268] = 25'b1111111000000010000111111;
    rom[22269] = 25'b1111111000000001000001000;
    rom[22270] = 25'b1111110111111111111010001;
    rom[22271] = 25'b1111110111111110110011011;
    rom[22272] = 25'b1111110111111101101100100;
    rom[22273] = 25'b1111110111111100100101101;
    rom[22274] = 25'b1111110111111011011110110;
    rom[22275] = 25'b1111110111111010011000000;
    rom[22276] = 25'b1111110111111001010001010;
    rom[22277] = 25'b1111110111111000001010100;
    rom[22278] = 25'b1111110111110111000011101;
    rom[22279] = 25'b1111110111110101111101000;
    rom[22280] = 25'b1111110111110100110110001;
    rom[22281] = 25'b1111110111110011101111100;
    rom[22282] = 25'b1111110111110010101000110;
    rom[22283] = 25'b1111110111110001100010001;
    rom[22284] = 25'b1111110111110000011011011;
    rom[22285] = 25'b1111110111101111010100110;
    rom[22286] = 25'b1111110111101110001110000;
    rom[22287] = 25'b1111110111101101000111011;
    rom[22288] = 25'b1111110111101100000000110;
    rom[22289] = 25'b1111110111101010111010001;
    rom[22290] = 25'b1111110111101001110011100;
    rom[22291] = 25'b1111110111101000101100111;
    rom[22292] = 25'b1111110111100111100110011;
    rom[22293] = 25'b1111110111100110011111110;
    rom[22294] = 25'b1111110111100101011001010;
    rom[22295] = 25'b1111110111100100010010110;
    rom[22296] = 25'b1111110111100011001100010;
    rom[22297] = 25'b1111110111100010000101110;
    rom[22298] = 25'b1111110111100000111111010;
    rom[22299] = 25'b1111110111011111111000110;
    rom[22300] = 25'b1111110111011110110010011;
    rom[22301] = 25'b1111110111011101101011111;
    rom[22302] = 25'b1111110111011100100101100;
    rom[22303] = 25'b1111110111011011011111001;
    rom[22304] = 25'b1111110111011010011000110;
    rom[22305] = 25'b1111110111011001010010010;
    rom[22306] = 25'b1111110111011000001100000;
    rom[22307] = 25'b1111110111010111000101101;
    rom[22308] = 25'b1111110111010101111111011;
    rom[22309] = 25'b1111110111010100111001000;
    rom[22310] = 25'b1111110111010011110010101;
    rom[22311] = 25'b1111110111010010101100011;
    rom[22312] = 25'b1111110111010001100110001;
    rom[22313] = 25'b1111110111010000011111111;
    rom[22314] = 25'b1111110111001111011001101;
    rom[22315] = 25'b1111110111001110010011100;
    rom[22316] = 25'b1111110111001101001101010;
    rom[22317] = 25'b1111110111001100000111001;
    rom[22318] = 25'b1111110111001011000001000;
    rom[22319] = 25'b1111110111001001111010111;
    rom[22320] = 25'b1111110111001000110100101;
    rom[22321] = 25'b1111110111000111101110100;
    rom[22322] = 25'b1111110111000110101000100;
    rom[22323] = 25'b1111110111000101100010011;
    rom[22324] = 25'b1111110111000100011100011;
    rom[22325] = 25'b1111110111000011010110010;
    rom[22326] = 25'b1111110111000010010000010;
    rom[22327] = 25'b1111110111000001001010010;
    rom[22328] = 25'b1111110111000000000100010;
    rom[22329] = 25'b1111110110111110111110011;
    rom[22330] = 25'b1111110110111101111000011;
    rom[22331] = 25'b1111110110111100110010100;
    rom[22332] = 25'b1111110110111011101100101;
    rom[22333] = 25'b1111110110111010100110110;
    rom[22334] = 25'b1111110110111001100000110;
    rom[22335] = 25'b1111110110111000011010111;
    rom[22336] = 25'b1111110110110111010101001;
    rom[22337] = 25'b1111110110110110001111010;
    rom[22338] = 25'b1111110110110101001001100;
    rom[22339] = 25'b1111110110110100000011110;
    rom[22340] = 25'b1111110110110010111110000;
    rom[22341] = 25'b1111110110110001111000010;
    rom[22342] = 25'b1111110110110000110010100;
    rom[22343] = 25'b1111110110101111101100111;
    rom[22344] = 25'b1111110110101110100111001;
    rom[22345] = 25'b1111110110101101100001100;
    rom[22346] = 25'b1111110110101100011011111;
    rom[22347] = 25'b1111110110101011010110010;
    rom[22348] = 25'b1111110110101010010000110;
    rom[22349] = 25'b1111110110101001001011001;
    rom[22350] = 25'b1111110110101000000101100;
    rom[22351] = 25'b1111110110100111000000000;
    rom[22352] = 25'b1111110110100101111010100;
    rom[22353] = 25'b1111110110100100110101000;
    rom[22354] = 25'b1111110110100011101111100;
    rom[22355] = 25'b1111110110100010101010000;
    rom[22356] = 25'b1111110110100001100100101;
    rom[22357] = 25'b1111110110100000011111010;
    rom[22358] = 25'b1111110110011111011001111;
    rom[22359] = 25'b1111110110011110010100100;
    rom[22360] = 25'b1111110110011101001111010;
    rom[22361] = 25'b1111110110011100001001111;
    rom[22362] = 25'b1111110110011011000100100;
    rom[22363] = 25'b1111110110011001111111010;
    rom[22364] = 25'b1111110110011000111010000;
    rom[22365] = 25'b1111110110010111110100110;
    rom[22366] = 25'b1111110110010110101111100;
    rom[22367] = 25'b1111110110010101101010011;
    rom[22368] = 25'b1111110110010100100101010;
    rom[22369] = 25'b1111110110010011100000000;
    rom[22370] = 25'b1111110110010010011010111;
    rom[22371] = 25'b1111110110010001010101111;
    rom[22372] = 25'b1111110110010000010000111;
    rom[22373] = 25'b1111110110001111001011110;
    rom[22374] = 25'b1111110110001110000110110;
    rom[22375] = 25'b1111110110001101000001101;
    rom[22376] = 25'b1111110110001011111100110;
    rom[22377] = 25'b1111110110001010110111110;
    rom[22378] = 25'b1111110110001001110010111;
    rom[22379] = 25'b1111110110001000101101111;
    rom[22380] = 25'b1111110110000111101001000;
    rom[22381] = 25'b1111110110000110100100001;
    rom[22382] = 25'b1111110110000101011111011;
    rom[22383] = 25'b1111110110000100011010100;
    rom[22384] = 25'b1111110110000011010101101;
    rom[22385] = 25'b1111110110000010010001000;
    rom[22386] = 25'b1111110110000001001100010;
    rom[22387] = 25'b1111110110000000000111100;
    rom[22388] = 25'b1111110101111111000010110;
    rom[22389] = 25'b1111110101111101111110001;
    rom[22390] = 25'b1111110101111100111001100;
    rom[22391] = 25'b1111110101111011110100111;
    rom[22392] = 25'b1111110101111010110000010;
    rom[22393] = 25'b1111110101111001101011110;
    rom[22394] = 25'b1111110101111000100111010;
    rom[22395] = 25'b1111110101110111100010101;
    rom[22396] = 25'b1111110101110110011110001;
    rom[22397] = 25'b1111110101110101011001101;
    rom[22398] = 25'b1111110101110100010101010;
    rom[22399] = 25'b1111110101110011010000111;
    rom[22400] = 25'b1111110101110010001100011;
    rom[22401] = 25'b1111110101110001001000000;
    rom[22402] = 25'b1111110101110000000011110;
    rom[22403] = 25'b1111110101101110111111011;
    rom[22404] = 25'b1111110101101101111011001;
    rom[22405] = 25'b1111110101101100110110111;
    rom[22406] = 25'b1111110101101011110010101;
    rom[22407] = 25'b1111110101101010101110011;
    rom[22408] = 25'b1111110101101001101010010;
    rom[22409] = 25'b1111110101101000100110001;
    rom[22410] = 25'b1111110101100111100001111;
    rom[22411] = 25'b1111110101100110011101111;
    rom[22412] = 25'b1111110101100101011001110;
    rom[22413] = 25'b1111110101100100010101110;
    rom[22414] = 25'b1111110101100011010001110;
    rom[22415] = 25'b1111110101100010001101110;
    rom[22416] = 25'b1111110101100001001001110;
    rom[22417] = 25'b1111110101100000000101111;
    rom[22418] = 25'b1111110101011111000010000;
    rom[22419] = 25'b1111110101011101111110000;
    rom[22420] = 25'b1111110101011100111010001;
    rom[22421] = 25'b1111110101011011110110011;
    rom[22422] = 25'b1111110101011010110010100;
    rom[22423] = 25'b1111110101011001101110110;
    rom[22424] = 25'b1111110101011000101011000;
    rom[22425] = 25'b1111110101010111100111011;
    rom[22426] = 25'b1111110101010110100011101;
    rom[22427] = 25'b1111110101010101100000000;
    rom[22428] = 25'b1111110101010100011100011;
    rom[22429] = 25'b1111110101010011011000110;
    rom[22430] = 25'b1111110101010010010101010;
    rom[22431] = 25'b1111110101010001010001101;
    rom[22432] = 25'b1111110101010000001110001;
    rom[22433] = 25'b1111110101001111001010110;
    rom[22434] = 25'b1111110101001110000111010;
    rom[22435] = 25'b1111110101001101000011110;
    rom[22436] = 25'b1111110101001100000000100;
    rom[22437] = 25'b1111110101001010111101001;
    rom[22438] = 25'b1111110101001001111001110;
    rom[22439] = 25'b1111110101001000110110100;
    rom[22440] = 25'b1111110101000111110011010;
    rom[22441] = 25'b1111110101000110110000000;
    rom[22442] = 25'b1111110101000101101100110;
    rom[22443] = 25'b1111110101000100101001100;
    rom[22444] = 25'b1111110101000011100110011;
    rom[22445] = 25'b1111110101000010100011010;
    rom[22446] = 25'b1111110101000001100000001;
    rom[22447] = 25'b1111110101000000011101001;
    rom[22448] = 25'b1111110100111111011010000;
    rom[22449] = 25'b1111110100111110010111001;
    rom[22450] = 25'b1111110100111101010100001;
    rom[22451] = 25'b1111110100111100010001001;
    rom[22452] = 25'b1111110100111011001110011;
    rom[22453] = 25'b1111110100111010001011100;
    rom[22454] = 25'b1111110100111001001000101;
    rom[22455] = 25'b1111110100111000000101110;
    rom[22456] = 25'b1111110100110111000011000;
    rom[22457] = 25'b1111110100110110000000010;
    rom[22458] = 25'b1111110100110100111101101;
    rom[22459] = 25'b1111110100110011111010111;
    rom[22460] = 25'b1111110100110010111000010;
    rom[22461] = 25'b1111110100110001110101101;
    rom[22462] = 25'b1111110100110000110011001;
    rom[22463] = 25'b1111110100101111110000100;
    rom[22464] = 25'b1111110100101110101110000;
    rom[22465] = 25'b1111110100101101101011100;
    rom[22466] = 25'b1111110100101100101001000;
    rom[22467] = 25'b1111110100101011100110101;
    rom[22468] = 25'b1111110100101010100100010;
    rom[22469] = 25'b1111110100101001100001111;
    rom[22470] = 25'b1111110100101000011111100;
    rom[22471] = 25'b1111110100100111011101010;
    rom[22472] = 25'b1111110100100110011011000;
    rom[22473] = 25'b1111110100100101011000110;
    rom[22474] = 25'b1111110100100100010110101;
    rom[22475] = 25'b1111110100100011010100100;
    rom[22476] = 25'b1111110100100010010010011;
    rom[22477] = 25'b1111110100100001010000010;
    rom[22478] = 25'b1111110100100000001110001;
    rom[22479] = 25'b1111110100011111001100001;
    rom[22480] = 25'b1111110100011110001010010;
    rom[22481] = 25'b1111110100011101001000010;
    rom[22482] = 25'b1111110100011100000110011;
    rom[22483] = 25'b1111110100011011000100011;
    rom[22484] = 25'b1111110100011010000010101;
    rom[22485] = 25'b1111110100011001000000111;
    rom[22486] = 25'b1111110100010111111111000;
    rom[22487] = 25'b1111110100010110111101010;
    rom[22488] = 25'b1111110100010101111011101;
    rom[22489] = 25'b1111110100010100111010000;
    rom[22490] = 25'b1111110100010011111000011;
    rom[22491] = 25'b1111110100010010110110101;
    rom[22492] = 25'b1111110100010001110101001;
    rom[22493] = 25'b1111110100010000110011101;
    rom[22494] = 25'b1111110100001111110010001;
    rom[22495] = 25'b1111110100001110110000110;
    rom[22496] = 25'b1111110100001101101111010;
    rom[22497] = 25'b1111110100001100101101111;
    rom[22498] = 25'b1111110100001011101100100;
    rom[22499] = 25'b1111110100001010101011010;
    rom[22500] = 25'b1111110100001001101010000;
    rom[22501] = 25'b1111110100001000101000101;
    rom[22502] = 25'b1111110100000111100111100;
    rom[22503] = 25'b1111110100000110100110011;
    rom[22504] = 25'b1111110100000101100101010;
    rom[22505] = 25'b1111110100000100100100001;
    rom[22506] = 25'b1111110100000011100011001;
    rom[22507] = 25'b1111110100000010100010000;
    rom[22508] = 25'b1111110100000001100001001;
    rom[22509] = 25'b1111110100000000100000001;
    rom[22510] = 25'b1111110011111111011111010;
    rom[22511] = 25'b1111110011111110011110011;
    rom[22512] = 25'b1111110011111101011101101;
    rom[22513] = 25'b1111110011111100011100110;
    rom[22514] = 25'b1111110011111011011100000;
    rom[22515] = 25'b1111110011111010011011011;
    rom[22516] = 25'b1111110011111001011010101;
    rom[22517] = 25'b1111110011111000011010000;
    rom[22518] = 25'b1111110011110111011001011;
    rom[22519] = 25'b1111110011110110011000111;
    rom[22520] = 25'b1111110011110101011000011;
    rom[22521] = 25'b1111110011110100010111111;
    rom[22522] = 25'b1111110011110011010111011;
    rom[22523] = 25'b1111110011110010010111000;
    rom[22524] = 25'b1111110011110001010110101;
    rom[22525] = 25'b1111110011110000010110011;
    rom[22526] = 25'b1111110011101111010110000;
    rom[22527] = 25'b1111110011101110010101110;
    rom[22528] = 25'b1111110011101101010101101;
    rom[22529] = 25'b1111110011101100010101100;
    rom[22530] = 25'b1111110011101011010101010;
    rom[22531] = 25'b1111110011101010010101010;
    rom[22532] = 25'b1111110011101001010101001;
    rom[22533] = 25'b1111110011101000010101001;
    rom[22534] = 25'b1111110011100111010101001;
    rom[22535] = 25'b1111110011100110010101010;
    rom[22536] = 25'b1111110011100101010101011;
    rom[22537] = 25'b1111110011100100010101100;
    rom[22538] = 25'b1111110011100011010101110;
    rom[22539] = 25'b1111110011100010010101111;
    rom[22540] = 25'b1111110011100001010110001;
    rom[22541] = 25'b1111110011100000010110100;
    rom[22542] = 25'b1111110011011111010110111;
    rom[22543] = 25'b1111110011011110010111010;
    rom[22544] = 25'b1111110011011101010111101;
    rom[22545] = 25'b1111110011011100011000001;
    rom[22546] = 25'b1111110011011011011000101;
    rom[22547] = 25'b1111110011011010011001010;
    rom[22548] = 25'b1111110011011001011001111;
    rom[22549] = 25'b1111110011011000011010100;
    rom[22550] = 25'b1111110011010111011011010;
    rom[22551] = 25'b1111110011010110011011111;
    rom[22552] = 25'b1111110011010101011100101;
    rom[22553] = 25'b1111110011010100011101100;
    rom[22554] = 25'b1111110011010011011110010;
    rom[22555] = 25'b1111110011010010011111010;
    rom[22556] = 25'b1111110011010001100000001;
    rom[22557] = 25'b1111110011010000100001010;
    rom[22558] = 25'b1111110011001111100010001;
    rom[22559] = 25'b1111110011001110100011010;
    rom[22560] = 25'b1111110011001101100100011;
    rom[22561] = 25'b1111110011001100100101100;
    rom[22562] = 25'b1111110011001011100110101;
    rom[22563] = 25'b1111110011001010100111111;
    rom[22564] = 25'b1111110011001001101001010;
    rom[22565] = 25'b1111110011001000101010101;
    rom[22566] = 25'b1111110011000111101011111;
    rom[22567] = 25'b1111110011000110101101011;
    rom[22568] = 25'b1111110011000101101110110;
    rom[22569] = 25'b1111110011000100110000011;
    rom[22570] = 25'b1111110011000011110001111;
    rom[22571] = 25'b1111110011000010110011100;
    rom[22572] = 25'b1111110011000001110101001;
    rom[22573] = 25'b1111110011000000110110110;
    rom[22574] = 25'b1111110010111111111000100;
    rom[22575] = 25'b1111110010111110111010010;
    rom[22576] = 25'b1111110010111101111100000;
    rom[22577] = 25'b1111110010111100111101111;
    rom[22578] = 25'b1111110010111011111111110;
    rom[22579] = 25'b1111110010111011000001110;
    rom[22580] = 25'b1111110010111010000011110;
    rom[22581] = 25'b1111110010111001000101110;
    rom[22582] = 25'b1111110010111000000111111;
    rom[22583] = 25'b1111110010110111001010000;
    rom[22584] = 25'b1111110010110110001100001;
    rom[22585] = 25'b1111110010110101001110010;
    rom[22586] = 25'b1111110010110100010000101;
    rom[22587] = 25'b1111110010110011010010111;
    rom[22588] = 25'b1111110010110010010101010;
    rom[22589] = 25'b1111110010110001010111101;
    rom[22590] = 25'b1111110010110000011010001;
    rom[22591] = 25'b1111110010101111011100101;
    rom[22592] = 25'b1111110010101110011111001;
    rom[22593] = 25'b1111110010101101100001101;
    rom[22594] = 25'b1111110010101100100100011;
    rom[22595] = 25'b1111110010101011100111000;
    rom[22596] = 25'b1111110010101010101001110;
    rom[22597] = 25'b1111110010101001101100100;
    rom[22598] = 25'b1111110010101000101111010;
    rom[22599] = 25'b1111110010100111110010010;
    rom[22600] = 25'b1111110010100110110101000;
    rom[22601] = 25'b1111110010100101111000000;
    rom[22602] = 25'b1111110010100100111011001;
    rom[22603] = 25'b1111110010100011111110001;
    rom[22604] = 25'b1111110010100011000001010;
    rom[22605] = 25'b1111110010100010000100011;
    rom[22606] = 25'b1111110010100001000111100;
    rom[22607] = 25'b1111110010100000001010110;
    rom[22608] = 25'b1111110010011111001110000;
    rom[22609] = 25'b1111110010011110010001011;
    rom[22610] = 25'b1111110010011101010100110;
    rom[22611] = 25'b1111110010011100011000010;
    rom[22612] = 25'b1111110010011011011011110;
    rom[22613] = 25'b1111110010011010011111010;
    rom[22614] = 25'b1111110010011001100010111;
    rom[22615] = 25'b1111110010011000100110011;
    rom[22616] = 25'b1111110010010111101010001;
    rom[22617] = 25'b1111110010010110101101111;
    rom[22618] = 25'b1111110010010101110001101;
    rom[22619] = 25'b1111110010010100110101011;
    rom[22620] = 25'b1111110010010011111001011;
    rom[22621] = 25'b1111110010010010111101010;
    rom[22622] = 25'b1111110010010010000001001;
    rom[22623] = 25'b1111110010010001000101010;
    rom[22624] = 25'b1111110010010000001001010;
    rom[22625] = 25'b1111110010001111001101011;
    rom[22626] = 25'b1111110010001110010001101;
    rom[22627] = 25'b1111110010001101010101110;
    rom[22628] = 25'b1111110010001100011010001;
    rom[22629] = 25'b1111110010001011011110011;
    rom[22630] = 25'b1111110010001010100010110;
    rom[22631] = 25'b1111110010001001100111001;
    rom[22632] = 25'b1111110010001000101011101;
    rom[22633] = 25'b1111110010000111110000001;
    rom[22634] = 25'b1111110010000110110100110;
    rom[22635] = 25'b1111110010000101111001011;
    rom[22636] = 25'b1111110010000100111110000;
    rom[22637] = 25'b1111110010000100000010110;
    rom[22638] = 25'b1111110010000011000111100;
    rom[22639] = 25'b1111110010000010001100011;
    rom[22640] = 25'b1111110010000001010001010;
    rom[22641] = 25'b1111110010000000010110001;
    rom[22642] = 25'b1111110001111111011011001;
    rom[22643] = 25'b1111110001111110100000010;
    rom[22644] = 25'b1111110001111101100101010;
    rom[22645] = 25'b1111110001111100101010011;
    rom[22646] = 25'b1111110001111011101111101;
    rom[22647] = 25'b1111110001111010110100111;
    rom[22648] = 25'b1111110001111001111010001;
    rom[22649] = 25'b1111110001111000111111100;
    rom[22650] = 25'b1111110001111000000100111;
    rom[22651] = 25'b1111110001110111001010010;
    rom[22652] = 25'b1111110001110110001111111;
    rom[22653] = 25'b1111110001110101010101011;
    rom[22654] = 25'b1111110001110100011011000;
    rom[22655] = 25'b1111110001110011100000101;
    rom[22656] = 25'b1111110001110010100110011;
    rom[22657] = 25'b1111110001110001101100001;
    rom[22658] = 25'b1111110001110000110001111;
    rom[22659] = 25'b1111110001101111110111110;
    rom[22660] = 25'b1111110001101110111101110;
    rom[22661] = 25'b1111110001101110000011110;
    rom[22662] = 25'b1111110001101101001001110;
    rom[22663] = 25'b1111110001101100001111111;
    rom[22664] = 25'b1111110001101011010101111;
    rom[22665] = 25'b1111110001101010011100001;
    rom[22666] = 25'b1111110001101001100010011;
    rom[22667] = 25'b1111110001101000101000110;
    rom[22668] = 25'b1111110001100111101111001;
    rom[22669] = 25'b1111110001100110110101100;
    rom[22670] = 25'b1111110001100101111011111;
    rom[22671] = 25'b1111110001100101000010011;
    rom[22672] = 25'b1111110001100100001001000;
    rom[22673] = 25'b1111110001100011001111101;
    rom[22674] = 25'b1111110001100010010110010;
    rom[22675] = 25'b1111110001100001011101000;
    rom[22676] = 25'b1111110001100000100011110;
    rom[22677] = 25'b1111110001011111101010101;
    rom[22678] = 25'b1111110001011110110001101;
    rom[22679] = 25'b1111110001011101111000100;
    rom[22680] = 25'b1111110001011100111111101;
    rom[22681] = 25'b1111110001011100000110101;
    rom[22682] = 25'b1111110001011011001101110;
    rom[22683] = 25'b1111110001011010010101000;
    rom[22684] = 25'b1111110001011001011100001;
    rom[22685] = 25'b1111110001011000100011100;
    rom[22686] = 25'b1111110001010111101010110;
    rom[22687] = 25'b1111110001010110110010010;
    rom[22688] = 25'b1111110001010101111001110;
    rom[22689] = 25'b1111110001010101000001010;
    rom[22690] = 25'b1111110001010100001000110;
    rom[22691] = 25'b1111110001010011010000011;
    rom[22692] = 25'b1111110001010010011000001;
    rom[22693] = 25'b1111110001010001011111111;
    rom[22694] = 25'b1111110001010000100111101;
    rom[22695] = 25'b1111110001001111101111100;
    rom[22696] = 25'b1111110001001110110111011;
    rom[22697] = 25'b1111110001001101111111011;
    rom[22698] = 25'b1111110001001101000111011;
    rom[22699] = 25'b1111110001001100001111100;
    rom[22700] = 25'b1111110001001011010111101;
    rom[22701] = 25'b1111110001001010011111110;
    rom[22702] = 25'b1111110001001001101000000;
    rom[22703] = 25'b1111110001001000110000011;
    rom[22704] = 25'b1111110001000111111000111;
    rom[22705] = 25'b1111110001000111000001010;
    rom[22706] = 25'b1111110001000110001001101;
    rom[22707] = 25'b1111110001000101010010010;
    rom[22708] = 25'b1111110001000100011010111;
    rom[22709] = 25'b1111110001000011100011100;
    rom[22710] = 25'b1111110001000010101100010;
    rom[22711] = 25'b1111110001000001110101000;
    rom[22712] = 25'b1111110001000000111101111;
    rom[22713] = 25'b1111110001000000000110110;
    rom[22714] = 25'b1111110000111111001111101;
    rom[22715] = 25'b1111110000111110011000110;
    rom[22716] = 25'b1111110000111101100001111;
    rom[22717] = 25'b1111110000111100101011000;
    rom[22718] = 25'b1111110000111011110100001;
    rom[22719] = 25'b1111110000111010111101011;
    rom[22720] = 25'b1111110000111010000110101;
    rom[22721] = 25'b1111110000111001010000000;
    rom[22722] = 25'b1111110000111000011001100;
    rom[22723] = 25'b1111110000110111100011000;
    rom[22724] = 25'b1111110000110110101100100;
    rom[22725] = 25'b1111110000110101110110001;
    rom[22726] = 25'b1111110000110100111111111;
    rom[22727] = 25'b1111110000110100001001101;
    rom[22728] = 25'b1111110000110011010011011;
    rom[22729] = 25'b1111110000110010011101010;
    rom[22730] = 25'b1111110000110001100111001;
    rom[22731] = 25'b1111110000110000110001001;
    rom[22732] = 25'b1111110000101111111011010;
    rom[22733] = 25'b1111110000101111000101010;
    rom[22734] = 25'b1111110000101110001111100;
    rom[22735] = 25'b1111110000101101011001101;
    rom[22736] = 25'b1111110000101100100100000;
    rom[22737] = 25'b1111110000101011101110010;
    rom[22738] = 25'b1111110000101010111000101;
    rom[22739] = 25'b1111110000101010000011001;
    rom[22740] = 25'b1111110000101001001101101;
    rom[22741] = 25'b1111110000101000011000010;
    rom[22742] = 25'b1111110000100111100010111;
    rom[22743] = 25'b1111110000100110101101101;
    rom[22744] = 25'b1111110000100101111000011;
    rom[22745] = 25'b1111110000100101000011010;
    rom[22746] = 25'b1111110000100100001110001;
    rom[22747] = 25'b1111110000100011011001001;
    rom[22748] = 25'b1111110000100010100100001;
    rom[22749] = 25'b1111110000100001101111010;
    rom[22750] = 25'b1111110000100000111010011;
    rom[22751] = 25'b1111110000100000000101100;
    rom[22752] = 25'b1111110000011111010000111;
    rom[22753] = 25'b1111110000011110011100001;
    rom[22754] = 25'b1111110000011101100111101;
    rom[22755] = 25'b1111110000011100110011000;
    rom[22756] = 25'b1111110000011011111110100;
    rom[22757] = 25'b1111110000011011001010001;
    rom[22758] = 25'b1111110000011010010101110;
    rom[22759] = 25'b1111110000011001100001100;
    rom[22760] = 25'b1111110000011000101101010;
    rom[22761] = 25'b1111110000010111111001001;
    rom[22762] = 25'b1111110000010111000101000;
    rom[22763] = 25'b1111110000010110010001000;
    rom[22764] = 25'b1111110000010101011101000;
    rom[22765] = 25'b1111110000010100101001001;
    rom[22766] = 25'b1111110000010011110101011;
    rom[22767] = 25'b1111110000010011000001100;
    rom[22768] = 25'b1111110000010010001101110;
    rom[22769] = 25'b1111110000010001011010001;
    rom[22770] = 25'b1111110000010000100110101;
    rom[22771] = 25'b1111110000001111110011001;
    rom[22772] = 25'b1111110000001110111111101;
    rom[22773] = 25'b1111110000001110001100010;
    rom[22774] = 25'b1111110000001101011000111;
    rom[22775] = 25'b1111110000001100100101101;
    rom[22776] = 25'b1111110000001011110010100;
    rom[22777] = 25'b1111110000001010111111010;
    rom[22778] = 25'b1111110000001010001100011;
    rom[22779] = 25'b1111110000001001011001011;
    rom[22780] = 25'b1111110000001000100110011;
    rom[22781] = 25'b1111110000000111110011100;
    rom[22782] = 25'b1111110000000111000000110;
    rom[22783] = 25'b1111110000000110001101111;
    rom[22784] = 25'b1111110000000101011011011;
    rom[22785] = 25'b1111110000000100101000110;
    rom[22786] = 25'b1111110000000011110110001;
    rom[22787] = 25'b1111110000000011000011110;
    rom[22788] = 25'b1111110000000010010001011;
    rom[22789] = 25'b1111110000000001011111000;
    rom[22790] = 25'b1111110000000000101100110;
    rom[22791] = 25'b1111101111111111111010100;
    rom[22792] = 25'b1111101111111111001000011;
    rom[22793] = 25'b1111101111111110010110010;
    rom[22794] = 25'b1111101111111101100100011;
    rom[22795] = 25'b1111101111111100110010011;
    rom[22796] = 25'b1111101111111100000000100;
    rom[22797] = 25'b1111101111111011001110110;
    rom[22798] = 25'b1111101111111010011101000;
    rom[22799] = 25'b1111101111111001101011010;
    rom[22800] = 25'b1111101111111000111001101;
    rom[22801] = 25'b1111101111111000001000001;
    rom[22802] = 25'b1111101111110111010110110;
    rom[22803] = 25'b1111101111110110100101011;
    rom[22804] = 25'b1111101111110101110100000;
    rom[22805] = 25'b1111101111110101000010110;
    rom[22806] = 25'b1111101111110100010001100;
    rom[22807] = 25'b1111101111110011100000011;
    rom[22808] = 25'b1111101111110010101111011;
    rom[22809] = 25'b1111101111110001111110011;
    rom[22810] = 25'b1111101111110001001101100;
    rom[22811] = 25'b1111101111110000011100110;
    rom[22812] = 25'b1111101111101111101011111;
    rom[22813] = 25'b1111101111101110111011010;
    rom[22814] = 25'b1111101111101110001010100;
    rom[22815] = 25'b1111101111101101011010000;
    rom[22816] = 25'b1111101111101100101001011;
    rom[22817] = 25'b1111101111101011111001000;
    rom[22818] = 25'b1111101111101011001000101;
    rom[22819] = 25'b1111101111101010011000011;
    rom[22820] = 25'b1111101111101001101000001;
    rom[22821] = 25'b1111101111101000111000000;
    rom[22822] = 25'b1111101111101000000111111;
    rom[22823] = 25'b1111101111100111010111111;
    rom[22824] = 25'b1111101111100110100111111;
    rom[22825] = 25'b1111101111100101111000001;
    rom[22826] = 25'b1111101111100101001000010;
    rom[22827] = 25'b1111101111100100011000101;
    rom[22828] = 25'b1111101111100011101000111;
    rom[22829] = 25'b1111101111100010111001010;
    rom[22830] = 25'b1111101111100010001001110;
    rom[22831] = 25'b1111101111100001011010011;
    rom[22832] = 25'b1111101111100000101010111;
    rom[22833] = 25'b1111101111011111111011101;
    rom[22834] = 25'b1111101111011111001100011;
    rom[22835] = 25'b1111101111011110011101010;
    rom[22836] = 25'b1111101111011101101110001;
    rom[22837] = 25'b1111101111011100111111001;
    rom[22838] = 25'b1111101111011100010000001;
    rom[22839] = 25'b1111101111011011100001010;
    rom[22840] = 25'b1111101111011010110010100;
    rom[22841] = 25'b1111101111011010000011101;
    rom[22842] = 25'b1111101111011001010101001;
    rom[22843] = 25'b1111101111011000100110100;
    rom[22844] = 25'b1111101111010111110111111;
    rom[22845] = 25'b1111101111010111001001100;
    rom[22846] = 25'b1111101111010110011011000;
    rom[22847] = 25'b1111101111010101101100110;
    rom[22848] = 25'b1111101111010100111110100;
    rom[22849] = 25'b1111101111010100010000011;
    rom[22850] = 25'b1111101111010011100010010;
    rom[22851] = 25'b1111101111010010110100010;
    rom[22852] = 25'b1111101111010010000110011;
    rom[22853] = 25'b1111101111010001011000011;
    rom[22854] = 25'b1111101111010000101010101;
    rom[22855] = 25'b1111101111001111111100111;
    rom[22856] = 25'b1111101111001111001111010;
    rom[22857] = 25'b1111101111001110100001101;
    rom[22858] = 25'b1111101111001101110100001;
    rom[22859] = 25'b1111101111001101000110101;
    rom[22860] = 25'b1111101111001100011001011;
    rom[22861] = 25'b1111101111001011101100001;
    rom[22862] = 25'b1111101111001010111110111;
    rom[22863] = 25'b1111101111001010010001101;
    rom[22864] = 25'b1111101111001001100100101;
    rom[22865] = 25'b1111101111001000110111101;
    rom[22866] = 25'b1111101111001000001010110;
    rom[22867] = 25'b1111101111000111011101111;
    rom[22868] = 25'b1111101111000110110001001;
    rom[22869] = 25'b1111101111000110000100100;
    rom[22870] = 25'b1111101111000101010111110;
    rom[22871] = 25'b1111101111000100101011010;
    rom[22872] = 25'b1111101111000011111110110;
    rom[22873] = 25'b1111101111000011010010011;
    rom[22874] = 25'b1111101111000010100110000;
    rom[22875] = 25'b1111101111000001111001111;
    rom[22876] = 25'b1111101111000001001101101;
    rom[22877] = 25'b1111101111000000100001100;
    rom[22878] = 25'b1111101110111111110101100;
    rom[22879] = 25'b1111101110111111001001100;
    rom[22880] = 25'b1111101110111110011101101;
    rom[22881] = 25'b1111101110111101110001111;
    rom[22882] = 25'b1111101110111101000110001;
    rom[22883] = 25'b1111101110111100011010100;
    rom[22884] = 25'b1111101110111011101110111;
    rom[22885] = 25'b1111101110111011000011011;
    rom[22886] = 25'b1111101110111010011000000;
    rom[22887] = 25'b1111101110111001101100101;
    rom[22888] = 25'b1111101110111001000001011;
    rom[22889] = 25'b1111101110111000010110010;
    rom[22890] = 25'b1111101110110111101011001;
    rom[22891] = 25'b1111101110110111000000000;
    rom[22892] = 25'b1111101110110110010101001;
    rom[22893] = 25'b1111101110110101101010010;
    rom[22894] = 25'b1111101110110100111111011;
    rom[22895] = 25'b1111101110110100010100101;
    rom[22896] = 25'b1111101110110011101010000;
    rom[22897] = 25'b1111101110110010111111011;
    rom[22898] = 25'b1111101110110010010100111;
    rom[22899] = 25'b1111101110110001101010100;
    rom[22900] = 25'b1111101110110001000000001;
    rom[22901] = 25'b1111101110110000010101111;
    rom[22902] = 25'b1111101110101111101011110;
    rom[22903] = 25'b1111101110101111000001101;
    rom[22904] = 25'b1111101110101110010111101;
    rom[22905] = 25'b1111101110101101101101100;
    rom[22906] = 25'b1111101110101101000011110;
    rom[22907] = 25'b1111101110101100011001111;
    rom[22908] = 25'b1111101110101011110000001;
    rom[22909] = 25'b1111101110101011000110100;
    rom[22910] = 25'b1111101110101010011100111;
    rom[22911] = 25'b1111101110101001110011100;
    rom[22912] = 25'b1111101110101001001010000;
    rom[22913] = 25'b1111101110101000100000110;
    rom[22914] = 25'b1111101110100111110111011;
    rom[22915] = 25'b1111101110100111001110010;
    rom[22916] = 25'b1111101110100110100101001;
    rom[22917] = 25'b1111101110100101111100001;
    rom[22918] = 25'b1111101110100101010011001;
    rom[22919] = 25'b1111101110100100101010011;
    rom[22920] = 25'b1111101110100100000001100;
    rom[22921] = 25'b1111101110100011011000111;
    rom[22922] = 25'b1111101110100010110000010;
    rom[22923] = 25'b1111101110100010000111101;
    rom[22924] = 25'b1111101110100001011111001;
    rom[22925] = 25'b1111101110100000110110110;
    rom[22926] = 25'b1111101110100000001110100;
    rom[22927] = 25'b1111101110011111100110010;
    rom[22928] = 25'b1111101110011110111110001;
    rom[22929] = 25'b1111101110011110010110001;
    rom[22930] = 25'b1111101110011101101110000;
    rom[22931] = 25'b1111101110011101000110001;
    rom[22932] = 25'b1111101110011100011110010;
    rom[22933] = 25'b1111101110011011110110101;
    rom[22934] = 25'b1111101110011011001110111;
    rom[22935] = 25'b1111101110011010100111010;
    rom[22936] = 25'b1111101110011001111111110;
    rom[22937] = 25'b1111101110011001011000011;
    rom[22938] = 25'b1111101110011000110001001;
    rom[22939] = 25'b1111101110011000001001110;
    rom[22940] = 25'b1111101110010111100010100;
    rom[22941] = 25'b1111101110010110111011100;
    rom[22942] = 25'b1111101110010110010100100;
    rom[22943] = 25'b1111101110010101101101100;
    rom[22944] = 25'b1111101110010101000110101;
    rom[22945] = 25'b1111101110010100011111111;
    rom[22946] = 25'b1111101110010011111001001;
    rom[22947] = 25'b1111101110010011010010101;
    rom[22948] = 25'b1111101110010010101100000;
    rom[22949] = 25'b1111101110010010000101100;
    rom[22950] = 25'b1111101110010001011111001;
    rom[22951] = 25'b1111101110010000111000111;
    rom[22952] = 25'b1111101110010000010010101;
    rom[22953] = 25'b1111101110001111101100101;
    rom[22954] = 25'b1111101110001111000110100;
    rom[22955] = 25'b1111101110001110100000100;
    rom[22956] = 25'b1111101110001101111010101;
    rom[22957] = 25'b1111101110001101010100111;
    rom[22958] = 25'b1111101110001100101111001;
    rom[22959] = 25'b1111101110001100001001100;
    rom[22960] = 25'b1111101110001011100100000;
    rom[22961] = 25'b1111101110001010111110100;
    rom[22962] = 25'b1111101110001010011001001;
    rom[22963] = 25'b1111101110001001110011111;
    rom[22964] = 25'b1111101110001001001110101;
    rom[22965] = 25'b1111101110001000101001100;
    rom[22966] = 25'b1111101110001000000100011;
    rom[22967] = 25'b1111101110000111011111100;
    rom[22968] = 25'b1111101110000110111010101;
    rom[22969] = 25'b1111101110000110010101110;
    rom[22970] = 25'b1111101110000101110001001;
    rom[22971] = 25'b1111101110000101001100100;
    rom[22972] = 25'b1111101110000100100111111;
    rom[22973] = 25'b1111101110000100000011011;
    rom[22974] = 25'b1111101110000011011111000;
    rom[22975] = 25'b1111101110000010111010101;
    rom[22976] = 25'b1111101110000010010110100;
    rom[22977] = 25'b1111101110000001110010011;
    rom[22978] = 25'b1111101110000001001110011;
    rom[22979] = 25'b1111101110000000101010011;
    rom[22980] = 25'b1111101110000000000110100;
    rom[22981] = 25'b1111101101111111100010101;
    rom[22982] = 25'b1111101101111110111111000;
    rom[22983] = 25'b1111101101111110011011011;
    rom[22984] = 25'b1111101101111101110111111;
    rom[22985] = 25'b1111101101111101010100011;
    rom[22986] = 25'b1111101101111100110001000;
    rom[22987] = 25'b1111101101111100001101110;
    rom[22988] = 25'b1111101101111011101010100;
    rom[22989] = 25'b1111101101111011000111100;
    rom[22990] = 25'b1111101101111010100100011;
    rom[22991] = 25'b1111101101111010000001011;
    rom[22992] = 25'b1111101101111001011110101;
    rom[22993] = 25'b1111101101111000111011111;
    rom[22994] = 25'b1111101101111000011001001;
    rom[22995] = 25'b1111101101110111110110100;
    rom[22996] = 25'b1111101101110111010100000;
    rom[22997] = 25'b1111101101110110110001101;
    rom[22998] = 25'b1111101101110110001111010;
    rom[22999] = 25'b1111101101110101101101000;
    rom[23000] = 25'b1111101101110101001010110;
    rom[23001] = 25'b1111101101110100101000110;
    rom[23002] = 25'b1111101101110100000110110;
    rom[23003] = 25'b1111101101110011100100111;
    rom[23004] = 25'b1111101101110011000011000;
    rom[23005] = 25'b1111101101110010100001010;
    rom[23006] = 25'b1111101101110001111111101;
    rom[23007] = 25'b1111101101110001011110000;
    rom[23008] = 25'b1111101101110000111100100;
    rom[23009] = 25'b1111101101110000011011010;
    rom[23010] = 25'b1111101101101111111001111;
    rom[23011] = 25'b1111101101101111011000101;
    rom[23012] = 25'b1111101101101110110111100;
    rom[23013] = 25'b1111101101101110010110100;
    rom[23014] = 25'b1111101101101101110101100;
    rom[23015] = 25'b1111101101101101010100101;
    rom[23016] = 25'b1111101101101100110011111;
    rom[23017] = 25'b1111101101101100010011010;
    rom[23018] = 25'b1111101101101011110010101;
    rom[23019] = 25'b1111101101101011010010000;
    rom[23020] = 25'b1111101101101010110001101;
    rom[23021] = 25'b1111101101101010010001010;
    rom[23022] = 25'b1111101101101001110001000;
    rom[23023] = 25'b1111101101101001010000111;
    rom[23024] = 25'b1111101101101000110000111;
    rom[23025] = 25'b1111101101101000010000110;
    rom[23026] = 25'b1111101101100111110000111;
    rom[23027] = 25'b1111101101100111010001001;
    rom[23028] = 25'b1111101101100110110001011;
    rom[23029] = 25'b1111101101100110010001101;
    rom[23030] = 25'b1111101101100101110010001;
    rom[23031] = 25'b1111101101100101010010110;
    rom[23032] = 25'b1111101101100100110011011;
    rom[23033] = 25'b1111101101100100010100001;
    rom[23034] = 25'b1111101101100011110100111;
    rom[23035] = 25'b1111101101100011010101110;
    rom[23036] = 25'b1111101101100010110110110;
    rom[23037] = 25'b1111101101100010010111111;
    rom[23038] = 25'b1111101101100001111001000;
    rom[23039] = 25'b1111101101100001011010010;
    rom[23040] = 25'b1111101101100000111011101;
    rom[23041] = 25'b1111101101100000011101001;
    rom[23042] = 25'b1111101101011111111110100;
    rom[23043] = 25'b1111101101011111100000001;
    rom[23044] = 25'b1111101101011111000001111;
    rom[23045] = 25'b1111101101011110100011101;
    rom[23046] = 25'b1111101101011110000101100;
    rom[23047] = 25'b1111101101011101100111100;
    rom[23048] = 25'b1111101101011101001001100;
    rom[23049] = 25'b1111101101011100101011110;
    rom[23050] = 25'b1111101101011100001110000;
    rom[23051] = 25'b1111101101011011110000011;
    rom[23052] = 25'b1111101101011011010010110;
    rom[23053] = 25'b1111101101011010110101010;
    rom[23054] = 25'b1111101101011010010111111;
    rom[23055] = 25'b1111101101011001111010101;
    rom[23056] = 25'b1111101101011001011101011;
    rom[23057] = 25'b1111101101011001000000010;
    rom[23058] = 25'b1111101101011000100011010;
    rom[23059] = 25'b1111101101011000000110010;
    rom[23060] = 25'b1111101101010111101001011;
    rom[23061] = 25'b1111101101010111001100101;
    rom[23062] = 25'b1111101101010110110000000;
    rom[23063] = 25'b1111101101010110010011011;
    rom[23064] = 25'b1111101101010101110110111;
    rom[23065] = 25'b1111101101010101011010100;
    rom[23066] = 25'b1111101101010100111110010;
    rom[23067] = 25'b1111101101010100100010000;
    rom[23068] = 25'b1111101101010100000101111;
    rom[23069] = 25'b1111101101010011101001111;
    rom[23070] = 25'b1111101101010011001110000;
    rom[23071] = 25'b1111101101010010110010001;
    rom[23072] = 25'b1111101101010010010110011;
    rom[23073] = 25'b1111101101010001111010110;
    rom[23074] = 25'b1111101101010001011111010;
    rom[23075] = 25'b1111101101010001000011110;
    rom[23076] = 25'b1111101101010000101000010;
    rom[23077] = 25'b1111101101010000001101000;
    rom[23078] = 25'b1111101101001111110001111;
    rom[23079] = 25'b1111101101001111010110110;
    rom[23080] = 25'b1111101101001110111011110;
    rom[23081] = 25'b1111101101001110100000110;
    rom[23082] = 25'b1111101101001110000110000;
    rom[23083] = 25'b1111101101001101101011010;
    rom[23084] = 25'b1111101101001101010000101;
    rom[23085] = 25'b1111101101001100110110001;
    rom[23086] = 25'b1111101101001100011011101;
    rom[23087] = 25'b1111101101001100000001010;
    rom[23088] = 25'b1111101101001011100111000;
    rom[23089] = 25'b1111101101001011001100111;
    rom[23090] = 25'b1111101101001010110010110;
    rom[23091] = 25'b1111101101001010011000110;
    rom[23092] = 25'b1111101101001001111110111;
    rom[23093] = 25'b1111101101001001100101001;
    rom[23094] = 25'b1111101101001001001011100;
    rom[23095] = 25'b1111101101001000110001110;
    rom[23096] = 25'b1111101101001000011000010;
    rom[23097] = 25'b1111101101000111111110111;
    rom[23098] = 25'b1111101101000111100101101;
    rom[23099] = 25'b1111101101000111001100011;
    rom[23100] = 25'b1111101101000110110011001;
    rom[23101] = 25'b1111101101000110011010001;
    rom[23102] = 25'b1111101101000110000001001;
    rom[23103] = 25'b1111101101000101101000011;
    rom[23104] = 25'b1111101101000101001111101;
    rom[23105] = 25'b1111101101000100110111000;
    rom[23106] = 25'b1111101101000100011110011;
    rom[23107] = 25'b1111101101000100000101111;
    rom[23108] = 25'b1111101101000011101101100;
    rom[23109] = 25'b1111101101000011010101010;
    rom[23110] = 25'b1111101101000010111101001;
    rom[23111] = 25'b1111101101000010100101000;
    rom[23112] = 25'b1111101101000010001101000;
    rom[23113] = 25'b1111101101000001110101001;
    rom[23114] = 25'b1111101101000001011101010;
    rom[23115] = 25'b1111101101000001000101100;
    rom[23116] = 25'b1111101101000000101101111;
    rom[23117] = 25'b1111101101000000010110011;
    rom[23118] = 25'b1111101100111111111110111;
    rom[23119] = 25'b1111101100111111100111101;
    rom[23120] = 25'b1111101100111111010000011;
    rom[23121] = 25'b1111101100111110111001010;
    rom[23122] = 25'b1111101100111110100010010;
    rom[23123] = 25'b1111101100111110001011010;
    rom[23124] = 25'b1111101100111101110100100;
    rom[23125] = 25'b1111101100111101011101101;
    rom[23126] = 25'b1111101100111101000111000;
    rom[23127] = 25'b1111101100111100110000100;
    rom[23128] = 25'b1111101100111100011010000;
    rom[23129] = 25'b1111101100111100000011101;
    rom[23130] = 25'b1111101100111011101101010;
    rom[23131] = 25'b1111101100111011010111001;
    rom[23132] = 25'b1111101100111011000001001;
    rom[23133] = 25'b1111101100111010101011001;
    rom[23134] = 25'b1111101100111010010101010;
    rom[23135] = 25'b1111101100111001111111100;
    rom[23136] = 25'b1111101100111001101001110;
    rom[23137] = 25'b1111101100111001010100001;
    rom[23138] = 25'b1111101100111000111110101;
    rom[23139] = 25'b1111101100111000101001010;
    rom[23140] = 25'b1111101100111000010100000;
    rom[23141] = 25'b1111101100110111111110110;
    rom[23142] = 25'b1111101100110111101001110;
    rom[23143] = 25'b1111101100110111010100101;
    rom[23144] = 25'b1111101100110110111111110;
    rom[23145] = 25'b1111101100110110101010111;
    rom[23146] = 25'b1111101100110110010110010;
    rom[23147] = 25'b1111101100110110000001101;
    rom[23148] = 25'b1111101100110101101101001;
    rom[23149] = 25'b1111101100110101011000101;
    rom[23150] = 25'b1111101100110101000100010;
    rom[23151] = 25'b1111101100110100110000001;
    rom[23152] = 25'b1111101100110100011100000;
    rom[23153] = 25'b1111101100110100001000000;
    rom[23154] = 25'b1111101100110011110100000;
    rom[23155] = 25'b1111101100110011100000010;
    rom[23156] = 25'b1111101100110011001100100;
    rom[23157] = 25'b1111101100110010111000110;
    rom[23158] = 25'b1111101100110010100101010;
    rom[23159] = 25'b1111101100110010010001111;
    rom[23160] = 25'b1111101100110001111110100;
    rom[23161] = 25'b1111101100110001101011010;
    rom[23162] = 25'b1111101100110001011000001;
    rom[23163] = 25'b1111101100110001000101001;
    rom[23164] = 25'b1111101100110000110010001;
    rom[23165] = 25'b1111101100110000011111010;
    rom[23166] = 25'b1111101100110000001100101;
    rom[23167] = 25'b1111101100101111111001111;
    rom[23168] = 25'b1111101100101111100111011;
    rom[23169] = 25'b1111101100101111010100111;
    rom[23170] = 25'b1111101100101111000010100;
    rom[23171] = 25'b1111101100101110110000010;
    rom[23172] = 25'b1111101100101110011110010;
    rom[23173] = 25'b1111101100101110001100001;
    rom[23174] = 25'b1111101100101101111010001;
    rom[23175] = 25'b1111101100101101101000010;
    rom[23176] = 25'b1111101100101101010110101;
    rom[23177] = 25'b1111101100101101000100111;
    rom[23178] = 25'b1111101100101100110011011;
    rom[23179] = 25'b1111101100101100100001111;
    rom[23180] = 25'b1111101100101100010000101;
    rom[23181] = 25'b1111101100101011111111011;
    rom[23182] = 25'b1111101100101011101110001;
    rom[23183] = 25'b1111101100101011011101001;
    rom[23184] = 25'b1111101100101011001100001;
    rom[23185] = 25'b1111101100101010111011011;
    rom[23186] = 25'b1111101100101010101010100;
    rom[23187] = 25'b1111101100101010011001111;
    rom[23188] = 25'b1111101100101010001001011;
    rom[23189] = 25'b1111101100101001111001000;
    rom[23190] = 25'b1111101100101001101000101;
    rom[23191] = 25'b1111101100101001011000011;
    rom[23192] = 25'b1111101100101001001000010;
    rom[23193] = 25'b1111101100101000111000001;
    rom[23194] = 25'b1111101100101000101000010;
    rom[23195] = 25'b1111101100101000011000011;
    rom[23196] = 25'b1111101100101000001000110;
    rom[23197] = 25'b1111101100100111111001000;
    rom[23198] = 25'b1111101100100111101001100;
    rom[23199] = 25'b1111101100100111011010001;
    rom[23200] = 25'b1111101100100111001010110;
    rom[23201] = 25'b1111101100100110111011100;
    rom[23202] = 25'b1111101100100110101100011;
    rom[23203] = 25'b1111101100100110011101011;
    rom[23204] = 25'b1111101100100110001110100;
    rom[23205] = 25'b1111101100100101111111101;
    rom[23206] = 25'b1111101100100101110000111;
    rom[23207] = 25'b1111101100100101100010010;
    rom[23208] = 25'b1111101100100101010011110;
    rom[23209] = 25'b1111101100100101000101011;
    rom[23210] = 25'b1111101100100100110111000;
    rom[23211] = 25'b1111101100100100101000111;
    rom[23212] = 25'b1111101100100100011010110;
    rom[23213] = 25'b1111101100100100001100110;
    rom[23214] = 25'b1111101100100011111110111;
    rom[23215] = 25'b1111101100100011110001000;
    rom[23216] = 25'b1111101100100011100011010;
    rom[23217] = 25'b1111101100100011010101110;
    rom[23218] = 25'b1111101100100011001000010;
    rom[23219] = 25'b1111101100100010111010111;
    rom[23220] = 25'b1111101100100010101101101;
    rom[23221] = 25'b1111101100100010100000011;
    rom[23222] = 25'b1111101100100010010011010;
    rom[23223] = 25'b1111101100100010000110010;
    rom[23224] = 25'b1111101100100001111001100;
    rom[23225] = 25'b1111101100100001101100101;
    rom[23226] = 25'b1111101100100001100000000;
    rom[23227] = 25'b1111101100100001010011100;
    rom[23228] = 25'b1111101100100001000111000;
    rom[23229] = 25'b1111101100100000111010101;
    rom[23230] = 25'b1111101100100000101110011;
    rom[23231] = 25'b1111101100100000100010010;
    rom[23232] = 25'b1111101100100000010110010;
    rom[23233] = 25'b1111101100100000001010010;
    rom[23234] = 25'b1111101100011111111110011;
    rom[23235] = 25'b1111101100011111110010101;
    rom[23236] = 25'b1111101100011111100111000;
    rom[23237] = 25'b1111101100011111011011100;
    rom[23238] = 25'b1111101100011111010000001;
    rom[23239] = 25'b1111101100011111000100110;
    rom[23240] = 25'b1111101100011110111001101;
    rom[23241] = 25'b1111101100011110101110100;
    rom[23242] = 25'b1111101100011110100011011;
    rom[23243] = 25'b1111101100011110011000100;
    rom[23244] = 25'b1111101100011110001101101;
    rom[23245] = 25'b1111101100011110000011000;
    rom[23246] = 25'b1111101100011101111000100;
    rom[23247] = 25'b1111101100011101101101111;
    rom[23248] = 25'b1111101100011101100011100;
    rom[23249] = 25'b1111101100011101011001010;
    rom[23250] = 25'b1111101100011101001111001;
    rom[23251] = 25'b1111101100011101000101000;
    rom[23252] = 25'b1111101100011100111011001;
    rom[23253] = 25'b1111101100011100110001010;
    rom[23254] = 25'b1111101100011100100111100;
    rom[23255] = 25'b1111101100011100011101110;
    rom[23256] = 25'b1111101100011100010100010;
    rom[23257] = 25'b1111101100011100001010111;
    rom[23258] = 25'b1111101100011100000001100;
    rom[23259] = 25'b1111101100011011111000011;
    rom[23260] = 25'b1111101100011011101111010;
    rom[23261] = 25'b1111101100011011100110001;
    rom[23262] = 25'b1111101100011011011101010;
    rom[23263] = 25'b1111101100011011010100100;
    rom[23264] = 25'b1111101100011011001011110;
    rom[23265] = 25'b1111101100011011000011010;
    rom[23266] = 25'b1111101100011010111010110;
    rom[23267] = 25'b1111101100011010110010010;
    rom[23268] = 25'b1111101100011010101010000;
    rom[23269] = 25'b1111101100011010100001111;
    rom[23270] = 25'b1111101100011010011001111;
    rom[23271] = 25'b1111101100011010010001110;
    rom[23272] = 25'b1111101100011010001010000;
    rom[23273] = 25'b1111101100011010000010010;
    rom[23274] = 25'b1111101100011001111010101;
    rom[23275] = 25'b1111101100011001110011001;
    rom[23276] = 25'b1111101100011001101011101;
    rom[23277] = 25'b1111101100011001100100011;
    rom[23278] = 25'b1111101100011001011101001;
    rom[23279] = 25'b1111101100011001010110000;
    rom[23280] = 25'b1111101100011001001111000;
    rom[23281] = 25'b1111101100011001001000001;
    rom[23282] = 25'b1111101100011001000001010;
    rom[23283] = 25'b1111101100011000111010101;
    rom[23284] = 25'b1111101100011000110100000;
    rom[23285] = 25'b1111101100011000101101101;
    rom[23286] = 25'b1111101100011000100111010;
    rom[23287] = 25'b1111101100011000100001000;
    rom[23288] = 25'b1111101100011000011010111;
    rom[23289] = 25'b1111101100011000010100110;
    rom[23290] = 25'b1111101100011000001110111;
    rom[23291] = 25'b1111101100011000001001001;
    rom[23292] = 25'b1111101100011000000011010;
    rom[23293] = 25'b1111101100010111111101110;
    rom[23294] = 25'b1111101100010111111000010;
    rom[23295] = 25'b1111101100010111110010111;
    rom[23296] = 25'b1111101100010111101101100;
    rom[23297] = 25'b1111101100010111101000011;
    rom[23298] = 25'b1111101100010111100011010;
    rom[23299] = 25'b1111101100010111011110011;
    rom[23300] = 25'b1111101100010111011001100;
    rom[23301] = 25'b1111101100010111010100110;
    rom[23302] = 25'b1111101100010111010000000;
    rom[23303] = 25'b1111101100010111001011100;
    rom[23304] = 25'b1111101100010111000111001;
    rom[23305] = 25'b1111101100010111000010110;
    rom[23306] = 25'b1111101100010110111110101;
    rom[23307] = 25'b1111101100010110111010100;
    rom[23308] = 25'b1111101100010110110110100;
    rom[23309] = 25'b1111101100010110110010101;
    rom[23310] = 25'b1111101100010110101110110;
    rom[23311] = 25'b1111101100010110101011001;
    rom[23312] = 25'b1111101100010110100111101;
    rom[23313] = 25'b1111101100010110100100001;
    rom[23314] = 25'b1111101100010110100000110;
    rom[23315] = 25'b1111101100010110011101101;
    rom[23316] = 25'b1111101100010110011010011;
    rom[23317] = 25'b1111101100010110010111100;
    rom[23318] = 25'b1111101100010110010100100;
    rom[23319] = 25'b1111101100010110010001110;
    rom[23320] = 25'b1111101100010110001111000;
    rom[23321] = 25'b1111101100010110001100011;
    rom[23322] = 25'b1111101100010110001010000;
    rom[23323] = 25'b1111101100010110000111101;
    rom[23324] = 25'b1111101100010110000101011;
    rom[23325] = 25'b1111101100010110000011001;
    rom[23326] = 25'b1111101100010110000001001;
    rom[23327] = 25'b1111101100010101111111010;
    rom[23328] = 25'b1111101100010101111101011;
    rom[23329] = 25'b1111101100010101111011110;
    rom[23330] = 25'b1111101100010101111010001;
    rom[23331] = 25'b1111101100010101111000101;
    rom[23332] = 25'b1111101100010101110111010;
    rom[23333] = 25'b1111101100010101110101111;
    rom[23334] = 25'b1111101100010101110100110;
    rom[23335] = 25'b1111101100010101110011101;
    rom[23336] = 25'b1111101100010101110010110;
    rom[23337] = 25'b1111101100010101110001111;
    rom[23338] = 25'b1111101100010101110001001;
    rom[23339] = 25'b1111101100010101110000101;
    rom[23340] = 25'b1111101100010101110000000;
    rom[23341] = 25'b1111101100010101101111101;
    rom[23342] = 25'b1111101100010101101111011;
    rom[23343] = 25'b1111101100010101101111010;
    rom[23344] = 25'b1111101100010101101111001;
    rom[23345] = 25'b1111101100010101101111010;
    rom[23346] = 25'b1111101100010101101111011;
    rom[23347] = 25'b1111101100010101101111101;
    rom[23348] = 25'b1111101100010101110000000;
    rom[23349] = 25'b1111101100010101110000100;
    rom[23350] = 25'b1111101100010101110001000;
    rom[23351] = 25'b1111101100010101110001110;
    rom[23352] = 25'b1111101100010101110010100;
    rom[23353] = 25'b1111101100010101110011100;
    rom[23354] = 25'b1111101100010101110100100;
    rom[23355] = 25'b1111101100010101110101101;
    rom[23356] = 25'b1111101100010101110111000;
    rom[23357] = 25'b1111101100010101111000011;
    rom[23358] = 25'b1111101100010101111001110;
    rom[23359] = 25'b1111101100010101111011011;
    rom[23360] = 25'b1111101100010101111101001;
    rom[23361] = 25'b1111101100010101111110111;
    rom[23362] = 25'b1111101100010110000000111;
    rom[23363] = 25'b1111101100010110000010110;
    rom[23364] = 25'b1111101100010110000101000;
    rom[23365] = 25'b1111101100010110000111010;
    rom[23366] = 25'b1111101100010110001001101;
    rom[23367] = 25'b1111101100010110001100000;
    rom[23368] = 25'b1111101100010110001110101;
    rom[23369] = 25'b1111101100010110010001011;
    rom[23370] = 25'b1111101100010110010100001;
    rom[23371] = 25'b1111101100010110010111001;
    rom[23372] = 25'b1111101100010110011010001;
    rom[23373] = 25'b1111101100010110011101010;
    rom[23374] = 25'b1111101100010110100000100;
    rom[23375] = 25'b1111101100010110100011111;
    rom[23376] = 25'b1111101100010110100111011;
    rom[23377] = 25'b1111101100010110101011000;
    rom[23378] = 25'b1111101100010110101110110;
    rom[23379] = 25'b1111101100010110110010011;
    rom[23380] = 25'b1111101100010110110110011;
    rom[23381] = 25'b1111101100010110111010100;
    rom[23382] = 25'b1111101100010110111110101;
    rom[23383] = 25'b1111101100010111000010111;
    rom[23384] = 25'b1111101100010111000111001;
    rom[23385] = 25'b1111101100010111001011101;
    rom[23386] = 25'b1111101100010111010000011;
    rom[23387] = 25'b1111101100010111010101000;
    rom[23388] = 25'b1111101100010111011001111;
    rom[23389] = 25'b1111101100010111011110110;
    rom[23390] = 25'b1111101100010111100011110;
    rom[23391] = 25'b1111101100010111101001000;
    rom[23392] = 25'b1111101100010111101110010;
    rom[23393] = 25'b1111101100010111110011101;
    rom[23394] = 25'b1111101100010111111001001;
    rom[23395] = 25'b1111101100010111111110110;
    rom[23396] = 25'b1111101100011000000100011;
    rom[23397] = 25'b1111101100011000001010010;
    rom[23398] = 25'b1111101100011000010000010;
    rom[23399] = 25'b1111101100011000010110010;
    rom[23400] = 25'b1111101100011000011100011;
    rom[23401] = 25'b1111101100011000100010101;
    rom[23402] = 25'b1111101100011000101001000;
    rom[23403] = 25'b1111101100011000101111101;
    rom[23404] = 25'b1111101100011000110110010;
    rom[23405] = 25'b1111101100011000111100111;
    rom[23406] = 25'b1111101100011001000011110;
    rom[23407] = 25'b1111101100011001001010110;
    rom[23408] = 25'b1111101100011001010001111;
    rom[23409] = 25'b1111101100011001011001000;
    rom[23410] = 25'b1111101100011001100000011;
    rom[23411] = 25'b1111101100011001100111110;
    rom[23412] = 25'b1111101100011001101111001;
    rom[23413] = 25'b1111101100011001110110111;
    rom[23414] = 25'b1111101100011001111110101;
    rom[23415] = 25'b1111101100011010000110011;
    rom[23416] = 25'b1111101100011010001110100;
    rom[23417] = 25'b1111101100011010010110100;
    rom[23418] = 25'b1111101100011010011110110;
    rom[23419] = 25'b1111101100011010100111000;
    rom[23420] = 25'b1111101100011010101111011;
    rom[23421] = 25'b1111101100011010111000000;
    rom[23422] = 25'b1111101100011011000000110;
    rom[23423] = 25'b1111101100011011001001011;
    rom[23424] = 25'b1111101100011011010010011;
    rom[23425] = 25'b1111101100011011011011010;
    rom[23426] = 25'b1111101100011011100100011;
    rom[23427] = 25'b1111101100011011101101101;
    rom[23428] = 25'b1111101100011011110111000;
    rom[23429] = 25'b1111101100011100000000011;
    rom[23430] = 25'b1111101100011100001010000;
    rom[23431] = 25'b1111101100011100010011101;
    rom[23432] = 25'b1111101100011100011101011;
    rom[23433] = 25'b1111101100011100100111011;
    rom[23434] = 25'b1111101100011100110001011;
    rom[23435] = 25'b1111101100011100111011100;
    rom[23436] = 25'b1111101100011101000101110;
    rom[23437] = 25'b1111101100011101010000001;
    rom[23438] = 25'b1111101100011101011010101;
    rom[23439] = 25'b1111101100011101100101001;
    rom[23440] = 25'b1111101100011101101111111;
    rom[23441] = 25'b1111101100011101111010110;
    rom[23442] = 25'b1111101100011110000101101;
    rom[23443] = 25'b1111101100011110010000101;
    rom[23444] = 25'b1111101100011110011011111;
    rom[23445] = 25'b1111101100011110100111001;
    rom[23446] = 25'b1111101100011110110010100;
    rom[23447] = 25'b1111101100011110111110000;
    rom[23448] = 25'b1111101100011111001001101;
    rom[23449] = 25'b1111101100011111010101011;
    rom[23450] = 25'b1111101100011111100001001;
    rom[23451] = 25'b1111101100011111101101010;
    rom[23452] = 25'b1111101100011111111001010;
    rom[23453] = 25'b1111101100100000000101011;
    rom[23454] = 25'b1111101100100000010001110;
    rom[23455] = 25'b1111101100100000011110001;
    rom[23456] = 25'b1111101100100000101010101;
    rom[23457] = 25'b1111101100100000110111011;
    rom[23458] = 25'b1111101100100001000100001;
    rom[23459] = 25'b1111101100100001010001000;
    rom[23460] = 25'b1111101100100001011110000;
    rom[23461] = 25'b1111101100100001101011001;
    rom[23462] = 25'b1111101100100001111000011;
    rom[23463] = 25'b1111101100100010000101101;
    rom[23464] = 25'b1111101100100010010011001;
    rom[23465] = 25'b1111101100100010100000110;
    rom[23466] = 25'b1111101100100010101110011;
    rom[23467] = 25'b1111101100100010111100001;
    rom[23468] = 25'b1111101100100011001010001;
    rom[23469] = 25'b1111101100100011011000001;
    rom[23470] = 25'b1111101100100011100110010;
    rom[23471] = 25'b1111101100100011110100100;
    rom[23472] = 25'b1111101100100100000010111;
    rom[23473] = 25'b1111101100100100010001011;
    rom[23474] = 25'b1111101100100100100000000;
    rom[23475] = 25'b1111101100100100101110110;
    rom[23476] = 25'b1111101100100100111101101;
    rom[23477] = 25'b1111101100100101001100100;
    rom[23478] = 25'b1111101100100101011011101;
    rom[23479] = 25'b1111101100100101101010110;
    rom[23480] = 25'b1111101100100101111010000;
    rom[23481] = 25'b1111101100100110001001011;
    rom[23482] = 25'b1111101100100110011001000;
    rom[23483] = 25'b1111101100100110101000101;
    rom[23484] = 25'b1111101100100110111000011;
    rom[23485] = 25'b1111101100100111001000010;
    rom[23486] = 25'b1111101100100111011000010;
    rom[23487] = 25'b1111101100100111101000011;
    rom[23488] = 25'b1111101100100111111000101;
    rom[23489] = 25'b1111101100101000001000111;
    rom[23490] = 25'b1111101100101000011001011;
    rom[23491] = 25'b1111101100101000101010000;
    rom[23492] = 25'b1111101100101000111010101;
    rom[23493] = 25'b1111101100101001001011100;
    rom[23494] = 25'b1111101100101001011100011;
    rom[23495] = 25'b1111101100101001101101011;
    rom[23496] = 25'b1111101100101001111110100;
    rom[23497] = 25'b1111101100101010001111111;
    rom[23498] = 25'b1111101100101010100001010;
    rom[23499] = 25'b1111101100101010110010101;
    rom[23500] = 25'b1111101100101011000100011;
    rom[23501] = 25'b1111101100101011010110001;
    rom[23502] = 25'b1111101100101011100111111;
    rom[23503] = 25'b1111101100101011111001111;
    rom[23504] = 25'b1111101100101100001100000;
    rom[23505] = 25'b1111101100101100011110001;
    rom[23506] = 25'b1111101100101100110000100;
    rom[23507] = 25'b1111101100101101000010111;
    rom[23508] = 25'b1111101100101101010101100;
    rom[23509] = 25'b1111101100101101101000001;
    rom[23510] = 25'b1111101100101101111010111;
    rom[23511] = 25'b1111101100101110001101110;
    rom[23512] = 25'b1111101100101110100000110;
    rom[23513] = 25'b1111101100101110110100000;
    rom[23514] = 25'b1111101100101111000111010;
    rom[23515] = 25'b1111101100101111011010100;
    rom[23516] = 25'b1111101100101111101110000;
    rom[23517] = 25'b1111101100110000000001100;
    rom[23518] = 25'b1111101100110000010101010;
    rom[23519] = 25'b1111101100110000101001001;
    rom[23520] = 25'b1111101100110000111101000;
    rom[23521] = 25'b1111101100110001010001001;
    rom[23522] = 25'b1111101100110001100101010;
    rom[23523] = 25'b1111101100110001111001100;
    rom[23524] = 25'b1111101100110010001110000;
    rom[23525] = 25'b1111101100110010100010100;
    rom[23526] = 25'b1111101100110010110111010;
    rom[23527] = 25'b1111101100110011001011111;
    rom[23528] = 25'b1111101100110011100000111;
    rom[23529] = 25'b1111101100110011110101111;
    rom[23530] = 25'b1111101100110100001011000;
    rom[23531] = 25'b1111101100110100100000001;
    rom[23532] = 25'b1111101100110100110101100;
    rom[23533] = 25'b1111101100110101001010111;
    rom[23534] = 25'b1111101100110101100000100;
    rom[23535] = 25'b1111101100110101110110010;
    rom[23536] = 25'b1111101100110110001100000;
    rom[23537] = 25'b1111101100110110100010000;
    rom[23538] = 25'b1111101100110110111000000;
    rom[23539] = 25'b1111101100110111001110010;
    rom[23540] = 25'b1111101100110111100100100;
    rom[23541] = 25'b1111101100110111111010111;
    rom[23542] = 25'b1111101100111000010001011;
    rom[23543] = 25'b1111101100111000101000001;
    rom[23544] = 25'b1111101100111000111110110;
    rom[23545] = 25'b1111101100111001010101101;
    rom[23546] = 25'b1111101100111001101100101;
    rom[23547] = 25'b1111101100111010000011110;
    rom[23548] = 25'b1111101100111010011011000;
    rom[23549] = 25'b1111101100111010110010010;
    rom[23550] = 25'b1111101100111011001001110;
    rom[23551] = 25'b1111101100111011100001011;
    rom[23552] = 25'b1111101100111011111001000;
    rom[23553] = 25'b1111101100111100010000110;
    rom[23554] = 25'b1111101100111100101000110;
    rom[23555] = 25'b1111101100111101000000110;
    rom[23556] = 25'b1111101100111101011001000;
    rom[23557] = 25'b1111101100111101110001010;
    rom[23558] = 25'b1111101100111110001001101;
    rom[23559] = 25'b1111101100111110100010001;
    rom[23560] = 25'b1111101100111110111010110;
    rom[23561] = 25'b1111101100111111010011100;
    rom[23562] = 25'b1111101100111111101100011;
    rom[23563] = 25'b1111101101000000000101011;
    rom[23564] = 25'b1111101101000000011110100;
    rom[23565] = 25'b1111101101000000110111110;
    rom[23566] = 25'b1111101101000001010001000;
    rom[23567] = 25'b1111101101000001101010011;
    rom[23568] = 25'b1111101101000010000100000;
    rom[23569] = 25'b1111101101000010011101110;
    rom[23570] = 25'b1111101101000010110111100;
    rom[23571] = 25'b1111101101000011010001011;
    rom[23572] = 25'b1111101101000011101011100;
    rom[23573] = 25'b1111101101000100000101101;
    rom[23574] = 25'b1111101101000100100000000;
    rom[23575] = 25'b1111101101000100111010010;
    rom[23576] = 25'b1111101101000101010100111;
    rom[23577] = 25'b1111101101000101101111011;
    rom[23578] = 25'b1111101101000110001010010;
    rom[23579] = 25'b1111101101000110100101000;
    rom[23580] = 25'b1111101101000111000000000;
    rom[23581] = 25'b1111101101000111011011010;
    rom[23582] = 25'b1111101101000111110110011;
    rom[23583] = 25'b1111101101001000010001110;
    rom[23584] = 25'b1111101101001000101101010;
    rom[23585] = 25'b1111101101001001001000110;
    rom[23586] = 25'b1111101101001001100100100;
    rom[23587] = 25'b1111101101001010000000010;
    rom[23588] = 25'b1111101101001010011100010;
    rom[23589] = 25'b1111101101001010111000010;
    rom[23590] = 25'b1111101101001011010100011;
    rom[23591] = 25'b1111101101001011110000101;
    rom[23592] = 25'b1111101101001100001101000;
    rom[23593] = 25'b1111101101001100101001101;
    rom[23594] = 25'b1111101101001101000110010;
    rom[23595] = 25'b1111101101001101100011000;
    rom[23596] = 25'b1111101101001101111111111;
    rom[23597] = 25'b1111101101001110011100111;
    rom[23598] = 25'b1111101101001110111010000;
    rom[23599] = 25'b1111101101001111010111010;
    rom[23600] = 25'b1111101101001111110100100;
    rom[23601] = 25'b1111101101010000010010000;
    rom[23602] = 25'b1111101101010000101111101;
    rom[23603] = 25'b1111101101010001001101010;
    rom[23604] = 25'b1111101101010001101011001;
    rom[23605] = 25'b1111101101010010001001000;
    rom[23606] = 25'b1111101101010010100111001;
    rom[23607] = 25'b1111101101010011000101010;
    rom[23608] = 25'b1111101101010011100011100;
    rom[23609] = 25'b1111101101010100000010000;
    rom[23610] = 25'b1111101101010100100000100;
    rom[23611] = 25'b1111101101010100111111001;
    rom[23612] = 25'b1111101101010101011110000;
    rom[23613] = 25'b1111101101010101111100110;
    rom[23614] = 25'b1111101101010110011011110;
    rom[23615] = 25'b1111101101010110111011000;
    rom[23616] = 25'b1111101101010111011010001;
    rom[23617] = 25'b1111101101010111111001100;
    rom[23618] = 25'b1111101101011000011001000;
    rom[23619] = 25'b1111101101011000111000101;
    rom[23620] = 25'b1111101101011001011000011;
    rom[23621] = 25'b1111101101011001111000001;
    rom[23622] = 25'b1111101101011010011000001;
    rom[23623] = 25'b1111101101011010111000001;
    rom[23624] = 25'b1111101101011011011000011;
    rom[23625] = 25'b1111101101011011111000101;
    rom[23626] = 25'b1111101101011100011001001;
    rom[23627] = 25'b1111101101011100111001101;
    rom[23628] = 25'b1111101101011101011010010;
    rom[23629] = 25'b1111101101011101111011000;
    rom[23630] = 25'b1111101101011110011011111;
    rom[23631] = 25'b1111101101011110111101000;
    rom[23632] = 25'b1111101101011111011110001;
    rom[23633] = 25'b1111101101011111111111011;
    rom[23634] = 25'b1111101101100000100000110;
    rom[23635] = 25'b1111101101100001000010010;
    rom[23636] = 25'b1111101101100001100011111;
    rom[23637] = 25'b1111101101100010000101101;
    rom[23638] = 25'b1111101101100010100111011;
    rom[23639] = 25'b1111101101100011001001011;
    rom[23640] = 25'b1111101101100011101011100;
    rom[23641] = 25'b1111101101100100001101101;
    rom[23642] = 25'b1111101101100100110000000;
    rom[23643] = 25'b1111101101100101010010100;
    rom[23644] = 25'b1111101101100101110101000;
    rom[23645] = 25'b1111101101100110010111101;
    rom[23646] = 25'b1111101101100110111010100;
    rom[23647] = 25'b1111101101100111011101011;
    rom[23648] = 25'b1111101101101000000000100;
    rom[23649] = 25'b1111101101101000100011100;
    rom[23650] = 25'b1111101101101001000110111;
    rom[23651] = 25'b1111101101101001101010010;
    rom[23652] = 25'b1111101101101010001101110;
    rom[23653] = 25'b1111101101101010110001011;
    rom[23654] = 25'b1111101101101011010101001;
    rom[23655] = 25'b1111101101101011111001000;
    rom[23656] = 25'b1111101101101100011100111;
    rom[23657] = 25'b1111101101101101000001000;
    rom[23658] = 25'b1111101101101101100101010;
    rom[23659] = 25'b1111101101101110001001101;
    rom[23660] = 25'b1111101101101110101110000;
    rom[23661] = 25'b1111101101101111010010101;
    rom[23662] = 25'b1111101101101111110111011;
    rom[23663] = 25'b1111101101110000011100001;
    rom[23664] = 25'b1111101101110001000001001;
    rom[23665] = 25'b1111101101110001100110001;
    rom[23666] = 25'b1111101101110010001011010;
    rom[23667] = 25'b1111101101110010110000101;
    rom[23668] = 25'b1111101101110011010110000;
    rom[23669] = 25'b1111101101110011111011100;
    rom[23670] = 25'b1111101101110100100001001;
    rom[23671] = 25'b1111101101110101000111000;
    rom[23672] = 25'b1111101101110101101100110;
    rom[23673] = 25'b1111101101110110010010110;
    rom[23674] = 25'b1111101101110110111000111;
    rom[23675] = 25'b1111101101110111011111001;
    rom[23676] = 25'b1111101101111000000101101;
    rom[23677] = 25'b1111101101111000101100000;
    rom[23678] = 25'b1111101101111001010010101;
    rom[23679] = 25'b1111101101111001111001010;
    rom[23680] = 25'b1111101101111010100000001;
    rom[23681] = 25'b1111101101111011000111001;
    rom[23682] = 25'b1111101101111011101110010;
    rom[23683] = 25'b1111101101111100010101011;
    rom[23684] = 25'b1111101101111100111100101;
    rom[23685] = 25'b1111101101111101100100000;
    rom[23686] = 25'b1111101101111110001011101;
    rom[23687] = 25'b1111101101111110110011011;
    rom[23688] = 25'b1111101101111111011011001;
    rom[23689] = 25'b1111101110000000000011000;
    rom[23690] = 25'b1111101110000000101011000;
    rom[23691] = 25'b1111101110000001010011001;
    rom[23692] = 25'b1111101110000001111011011;
    rom[23693] = 25'b1111101110000010100011110;
    rom[23694] = 25'b1111101110000011001100010;
    rom[23695] = 25'b1111101110000011110100111;
    rom[23696] = 25'b1111101110000100011101101;
    rom[23697] = 25'b1111101110000101000110100;
    rom[23698] = 25'b1111101110000101101111100;
    rom[23699] = 25'b1111101110000110011000101;
    rom[23700] = 25'b1111101110000111000001110;
    rom[23701] = 25'b1111101110000111101011000;
    rom[23702] = 25'b1111101110001000010100100;
    rom[23703] = 25'b1111101110001000111110000;
    rom[23704] = 25'b1111101110001001100111110;
    rom[23705] = 25'b1111101110001010010001100;
    rom[23706] = 25'b1111101110001010111011100;
    rom[23707] = 25'b1111101110001011100101100;
    rom[23708] = 25'b1111101110001100001111110;
    rom[23709] = 25'b1111101110001100111001111;
    rom[23710] = 25'b1111101110001101100100011;
    rom[23711] = 25'b1111101110001110001110111;
    rom[23712] = 25'b1111101110001110111001100;
    rom[23713] = 25'b1111101110001111100100010;
    rom[23714] = 25'b1111101110010000001111001;
    rom[23715] = 25'b1111101110010000111010001;
    rom[23716] = 25'b1111101110010001100101010;
    rom[23717] = 25'b1111101110010010010000100;
    rom[23718] = 25'b1111101110010010111011110;
    rom[23719] = 25'b1111101110010011100111010;
    rom[23720] = 25'b1111101110010100010010111;
    rom[23721] = 25'b1111101110010100111110100;
    rom[23722] = 25'b1111101110010101101010011;
    rom[23723] = 25'b1111101110010110010110011;
    rom[23724] = 25'b1111101110010111000010011;
    rom[23725] = 25'b1111101110010111101110101;
    rom[23726] = 25'b1111101110011000011010111;
    rom[23727] = 25'b1111101110011001000111010;
    rom[23728] = 25'b1111101110011001110011110;
    rom[23729] = 25'b1111101110011010100000011;
    rom[23730] = 25'b1111101110011011001101010;
    rom[23731] = 25'b1111101110011011111010000;
    rom[23732] = 25'b1111101110011100100111000;
    rom[23733] = 25'b1111101110011101010100010;
    rom[23734] = 25'b1111101110011110000001100;
    rom[23735] = 25'b1111101110011110101110111;
    rom[23736] = 25'b1111101110011111011100010;
    rom[23737] = 25'b1111101110100000001001111;
    rom[23738] = 25'b1111101110100000110111101;
    rom[23739] = 25'b1111101110100001100101011;
    rom[23740] = 25'b1111101110100010010011011;
    rom[23741] = 25'b1111101110100011000001100;
    rom[23742] = 25'b1111101110100011101111101;
    rom[23743] = 25'b1111101110100100011101111;
    rom[23744] = 25'b1111101110100101001100100;
    rom[23745] = 25'b1111101110100101111011000;
    rom[23746] = 25'b1111101110100110101001101;
    rom[23747] = 25'b1111101110100111011000011;
    rom[23748] = 25'b1111101110101000000111010;
    rom[23749] = 25'b1111101110101000110110010;
    rom[23750] = 25'b1111101110101001100101100;
    rom[23751] = 25'b1111101110101010010100110;
    rom[23752] = 25'b1111101110101011000100000;
    rom[23753] = 25'b1111101110101011110011101;
    rom[23754] = 25'b1111101110101100100011010;
    rom[23755] = 25'b1111101110101101010010111;
    rom[23756] = 25'b1111101110101110000010110;
    rom[23757] = 25'b1111101110101110110010110;
    rom[23758] = 25'b1111101110101111100010111;
    rom[23759] = 25'b1111101110110000010011000;
    rom[23760] = 25'b1111101110110001000011011;
    rom[23761] = 25'b1111101110110001110011110;
    rom[23762] = 25'b1111101110110010100100011;
    rom[23763] = 25'b1111101110110011010101000;
    rom[23764] = 25'b1111101110110100000101111;
    rom[23765] = 25'b1111101110110100110110110;
    rom[23766] = 25'b1111101110110101100111110;
    rom[23767] = 25'b1111101110110110011000111;
    rom[23768] = 25'b1111101110110111001010010;
    rom[23769] = 25'b1111101110110111111011100;
    rom[23770] = 25'b1111101110111000101101001;
    rom[23771] = 25'b1111101110111001011110110;
    rom[23772] = 25'b1111101110111010010000100;
    rom[23773] = 25'b1111101110111011000010010;
    rom[23774] = 25'b1111101110111011110100011;
    rom[23775] = 25'b1111101110111100100110011;
    rom[23776] = 25'b1111101110111101011000101;
    rom[23777] = 25'b1111101110111110001011000;
    rom[23778] = 25'b1111101110111110111101011;
    rom[23779] = 25'b1111101110111111101111111;
    rom[23780] = 25'b1111101111000000100010101;
    rom[23781] = 25'b1111101111000001010101011;
    rom[23782] = 25'b1111101111000010001000010;
    rom[23783] = 25'b1111101111000010111011011;
    rom[23784] = 25'b1111101111000011101110101;
    rom[23785] = 25'b1111101111000100100001111;
    rom[23786] = 25'b1111101111000101010101010;
    rom[23787] = 25'b1111101111000110001000110;
    rom[23788] = 25'b1111101111000110111100011;
    rom[23789] = 25'b1111101111000111110000001;
    rom[23790] = 25'b1111101111001000100100000;
    rom[23791] = 25'b1111101111001001011000000;
    rom[23792] = 25'b1111101111001010001100001;
    rom[23793] = 25'b1111101111001011000000010;
    rom[23794] = 25'b1111101111001011110100101;
    rom[23795] = 25'b1111101111001100101001001;
    rom[23796] = 25'b1111101111001101011101101;
    rom[23797] = 25'b1111101111001110010010011;
    rom[23798] = 25'b1111101111001111000111001;
    rom[23799] = 25'b1111101111001111111100000;
    rom[23800] = 25'b1111101111010000110001001;
    rom[23801] = 25'b1111101111010001100110010;
    rom[23802] = 25'b1111101111010010011011100;
    rom[23803] = 25'b1111101111010011010001000;
    rom[23804] = 25'b1111101111010100000110100;
    rom[23805] = 25'b1111101111010100111100001;
    rom[23806] = 25'b1111101111010101110001111;
    rom[23807] = 25'b1111101111010110100111101;
    rom[23808] = 25'b1111101111010111011101101;
    rom[23809] = 25'b1111101111011000010011110;
    rom[23810] = 25'b1111101111011001001010000;
    rom[23811] = 25'b1111101111011010000000010;
    rom[23812] = 25'b1111101111011010110110110;
    rom[23813] = 25'b1111101111011011101101010;
    rom[23814] = 25'b1111101111011100100100000;
    rom[23815] = 25'b1111101111011101011010111;
    rom[23816] = 25'b1111101111011110010001110;
    rom[23817] = 25'b1111101111011111001000110;
    rom[23818] = 25'b1111101111100000000000000;
    rom[23819] = 25'b1111101111100000110111010;
    rom[23820] = 25'b1111101111100001101110101;
    rom[23821] = 25'b1111101111100010100110001;
    rom[23822] = 25'b1111101111100011011101110;
    rom[23823] = 25'b1111101111100100010101100;
    rom[23824] = 25'b1111101111100101001101011;
    rom[23825] = 25'b1111101111100110000101011;
    rom[23826] = 25'b1111101111100110111101011;
    rom[23827] = 25'b1111101111100111110101101;
    rom[23828] = 25'b1111101111101000101101111;
    rom[23829] = 25'b1111101111101001100110011;
    rom[23830] = 25'b1111101111101010011110111;
    rom[23831] = 25'b1111101111101011010111101;
    rom[23832] = 25'b1111101111101100010000100;
    rom[23833] = 25'b1111101111101101001001011;
    rom[23834] = 25'b1111101111101110000010011;
    rom[23835] = 25'b1111101111101110111011101;
    rom[23836] = 25'b1111101111101111110100111;
    rom[23837] = 25'b1111101111110000101110001;
    rom[23838] = 25'b1111101111110001100111101;
    rom[23839] = 25'b1111101111110010100001010;
    rom[23840] = 25'b1111101111110011011011000;
    rom[23841] = 25'b1111101111110100010100111;
    rom[23842] = 25'b1111101111110101001110111;
    rom[23843] = 25'b1111101111110110001000111;
    rom[23844] = 25'b1111101111110111000011001;
    rom[23845] = 25'b1111101111110111111101100;
    rom[23846] = 25'b1111101111111000110111111;
    rom[23847] = 25'b1111101111111001110010011;
    rom[23848] = 25'b1111101111111010101101001;
    rom[23849] = 25'b1111101111111011100111111;
    rom[23850] = 25'b1111101111111100100010110;
    rom[23851] = 25'b1111101111111101011101110;
    rom[23852] = 25'b1111101111111110011000111;
    rom[23853] = 25'b1111101111111111010100001;
    rom[23854] = 25'b1111110000000000001111100;
    rom[23855] = 25'b1111110000000001001011000;
    rom[23856] = 25'b1111110000000010000110101;
    rom[23857] = 25'b1111110000000011000010010;
    rom[23858] = 25'b1111110000000011111110001;
    rom[23859] = 25'b1111110000000100111010001;
    rom[23860] = 25'b1111110000000101110110001;
    rom[23861] = 25'b1111110000000110110010010;
    rom[23862] = 25'b1111110000000111101110101;
    rom[23863] = 25'b1111110000001000101011000;
    rom[23864] = 25'b1111110000001001100111100;
    rom[23865] = 25'b1111110000001010100100001;
    rom[23866] = 25'b1111110000001011100000111;
    rom[23867] = 25'b1111110000001100011101111;
    rom[23868] = 25'b1111110000001101011010110;
    rom[23869] = 25'b1111110000001110010111111;
    rom[23870] = 25'b1111110000001111010101001;
    rom[23871] = 25'b1111110000010000010010011;
    rom[23872] = 25'b1111110000010001001111111;
    rom[23873] = 25'b1111110000010010001101100;
    rom[23874] = 25'b1111110000010011001011001;
    rom[23875] = 25'b1111110000010100001000111;
    rom[23876] = 25'b1111110000010101000110111;
    rom[23877] = 25'b1111110000010110000100111;
    rom[23878] = 25'b1111110000010111000011000;
    rom[23879] = 25'b1111110000011000000001010;
    rom[23880] = 25'b1111110000011000111111101;
    rom[23881] = 25'b1111110000011001111110010;
    rom[23882] = 25'b1111110000011010111100110;
    rom[23883] = 25'b1111110000011011111011100;
    rom[23884] = 25'b1111110000011100111010011;
    rom[23885] = 25'b1111110000011101111001011;
    rom[23886] = 25'b1111110000011110111000011;
    rom[23887] = 25'b1111110000011111110111101;
    rom[23888] = 25'b1111110000100000110110111;
    rom[23889] = 25'b1111110000100001110110010;
    rom[23890] = 25'b1111110000100010110101110;
    rom[23891] = 25'b1111110000100011110101011;
    rom[23892] = 25'b1111110000100100110101010;
    rom[23893] = 25'b1111110000100101110101001;
    rom[23894] = 25'b1111110000100110110101000;
    rom[23895] = 25'b1111110000100111110101010;
    rom[23896] = 25'b1111110000101000110101100;
    rom[23897] = 25'b1111110000101001110101110;
    rom[23898] = 25'b1111110000101010110110010;
    rom[23899] = 25'b1111110000101011110110110;
    rom[23900] = 25'b1111110000101100110111100;
    rom[23901] = 25'b1111110000101101111000010;
    rom[23902] = 25'b1111110000101110111001010;
    rom[23903] = 25'b1111110000101111111010001;
    rom[23904] = 25'b1111110000110000111011011;
    rom[23905] = 25'b1111110000110001111100100;
    rom[23906] = 25'b1111110000110010111101111;
    rom[23907] = 25'b1111110000110011111111100;
    rom[23908] = 25'b1111110000110101000001000;
    rom[23909] = 25'b1111110000110110000010110;
    rom[23910] = 25'b1111110000110111000100101;
    rom[23911] = 25'b1111110000111000000110100;
    rom[23912] = 25'b1111110000111001001000101;
    rom[23913] = 25'b1111110000111010001010110;
    rom[23914] = 25'b1111110000111011001101000;
    rom[23915] = 25'b1111110000111100001111011;
    rom[23916] = 25'b1111110000111101010010000;
    rom[23917] = 25'b1111110000111110010100101;
    rom[23918] = 25'b1111110000111111010111011;
    rom[23919] = 25'b1111110001000000011010010;
    rom[23920] = 25'b1111110001000001011101001;
    rom[23921] = 25'b1111110001000010100000010;
    rom[23922] = 25'b1111110001000011100011100;
    rom[23923] = 25'b1111110001000100100110110;
    rom[23924] = 25'b1111110001000101101010010;
    rom[23925] = 25'b1111110001000110101101110;
    rom[23926] = 25'b1111110001000111110001011;
    rom[23927] = 25'b1111110001001000110101001;
    rom[23928] = 25'b1111110001001001111001000;
    rom[23929] = 25'b1111110001001010111101000;
    rom[23930] = 25'b1111110001001100000001010;
    rom[23931] = 25'b1111110001001101000101011;
    rom[23932] = 25'b1111110001001110001001110;
    rom[23933] = 25'b1111110001001111001110001;
    rom[23934] = 25'b1111110001010000010010110;
    rom[23935] = 25'b1111110001010001010111100;
    rom[23936] = 25'b1111110001010010011100010;
    rom[23937] = 25'b1111110001010011100001001;
    rom[23938] = 25'b1111110001010100100110001;
    rom[23939] = 25'b1111110001010101101011010;
    rom[23940] = 25'b1111110001010110110000100;
    rom[23941] = 25'b1111110001010111110101111;
    rom[23942] = 25'b1111110001011000111011010;
    rom[23943] = 25'b1111110001011010000001000;
    rom[23944] = 25'b1111110001011011000110101;
    rom[23945] = 25'b1111110001011100001100011;
    rom[23946] = 25'b1111110001011101010010011;
    rom[23947] = 25'b1111110001011110011000011;
    rom[23948] = 25'b1111110001011111011110100;
    rom[23949] = 25'b1111110001100000100100111;
    rom[23950] = 25'b1111110001100001101011001;
    rom[23951] = 25'b1111110001100010110001101;
    rom[23952] = 25'b1111110001100011111000010;
    rom[23953] = 25'b1111110001100100111111000;
    rom[23954] = 25'b1111110001100110000101111;
    rom[23955] = 25'b1111110001100111001100110;
    rom[23956] = 25'b1111110001101000010011110;
    rom[23957] = 25'b1111110001101001011011000;
    rom[23958] = 25'b1111110001101010100010010;
    rom[23959] = 25'b1111110001101011101001101;
    rom[23960] = 25'b1111110001101100110001001;
    rom[23961] = 25'b1111110001101101111000110;
    rom[23962] = 25'b1111110001101111000000100;
    rom[23963] = 25'b1111110001110000001000011;
    rom[23964] = 25'b1111110001110001010000010;
    rom[23965] = 25'b1111110001110010011000011;
    rom[23966] = 25'b1111110001110011100000100;
    rom[23967] = 25'b1111110001110100101000110;
    rom[23968] = 25'b1111110001110101110001001;
    rom[23969] = 25'b1111110001110110111001110;
    rom[23970] = 25'b1111110001111000000010010;
    rom[23971] = 25'b1111110001111001001011000;
    rom[23972] = 25'b1111110001111010010011111;
    rom[23973] = 25'b1111110001111011011100111;
    rom[23974] = 25'b1111110001111100100110000;
    rom[23975] = 25'b1111110001111101101111001;
    rom[23976] = 25'b1111110001111110111000100;
    rom[23977] = 25'b1111110010000000000001111;
    rom[23978] = 25'b1111110010000001001011011;
    rom[23979] = 25'b1111110010000010010101000;
    rom[23980] = 25'b1111110010000011011110110;
    rom[23981] = 25'b1111110010000100101000101;
    rom[23982] = 25'b1111110010000101110010101;
    rom[23983] = 25'b1111110010000110111100101;
    rom[23984] = 25'b1111110010001000000110110;
    rom[23985] = 25'b1111110010001001010001001;
    rom[23986] = 25'b1111110010001010011011100;
    rom[23987] = 25'b1111110010001011100110001;
    rom[23988] = 25'b1111110010001100110000101;
    rom[23989] = 25'b1111110010001101111011011;
    rom[23990] = 25'b1111110010001111000110010;
    rom[23991] = 25'b1111110010010000010001001;
    rom[23992] = 25'b1111110010010001011100010;
    rom[23993] = 25'b1111110010010010100111100;
    rom[23994] = 25'b1111110010010011110010110;
    rom[23995] = 25'b1111110010010100111110001;
    rom[23996] = 25'b1111110010010110001001110;
    rom[23997] = 25'b1111110010010111010101010;
    rom[23998] = 25'b1111110010011000100001000;
    rom[23999] = 25'b1111110010011001101100111;
    rom[24000] = 25'b1111110010011010111000111;
    rom[24001] = 25'b1111110010011100000100111;
    rom[24002] = 25'b1111110010011101010001001;
    rom[24003] = 25'b1111110010011110011101011;
    rom[24004] = 25'b1111110010011111101001110;
    rom[24005] = 25'b1111110010100000110110010;
    rom[24006] = 25'b1111110010100010000010111;
    rom[24007] = 25'b1111110010100011001111101;
    rom[24008] = 25'b1111110010100100011100100;
    rom[24009] = 25'b1111110010100101101001011;
    rom[24010] = 25'b1111110010100110110110100;
    rom[24011] = 25'b1111110010101000000011101;
    rom[24012] = 25'b1111110010101001010000111;
    rom[24013] = 25'b1111110010101010011110011;
    rom[24014] = 25'b1111110010101011101011111;
    rom[24015] = 25'b1111110010101100111001011;
    rom[24016] = 25'b1111110010101110000111001;
    rom[24017] = 25'b1111110010101111010100111;
    rom[24018] = 25'b1111110010110000100010111;
    rom[24019] = 25'b1111110010110001110001000;
    rom[24020] = 25'b1111110010110010111111001;
    rom[24021] = 25'b1111110010110100001101011;
    rom[24022] = 25'b1111110010110101011011110;
    rom[24023] = 25'b1111110010110110101010010;
    rom[24024] = 25'b1111110010110111111000111;
    rom[24025] = 25'b1111110010111001000111100;
    rom[24026] = 25'b1111110010111010010110010;
    rom[24027] = 25'b1111110010111011100101010;
    rom[24028] = 25'b1111110010111100110100010;
    rom[24029] = 25'b1111110010111110000011011;
    rom[24030] = 25'b1111110010111111010010101;
    rom[24031] = 25'b1111110011000000100010000;
    rom[24032] = 25'b1111110011000001110001011;
    rom[24033] = 25'b1111110011000011000001000;
    rom[24034] = 25'b1111110011000100010000101;
    rom[24035] = 25'b1111110011000101100000100;
    rom[24036] = 25'b1111110011000110110000011;
    rom[24037] = 25'b1111110011001000000000011;
    rom[24038] = 25'b1111110011001001010000100;
    rom[24039] = 25'b1111110011001010100000110;
    rom[24040] = 25'b1111110011001011110001000;
    rom[24041] = 25'b1111110011001101000001100;
    rom[24042] = 25'b1111110011001110010010000;
    rom[24043] = 25'b1111110011001111100010101;
    rom[24044] = 25'b1111110011010000110011011;
    rom[24045] = 25'b1111110011010010000100010;
    rom[24046] = 25'b1111110011010011010101010;
    rom[24047] = 25'b1111110011010100100110010;
    rom[24048] = 25'b1111110011010101110111100;
    rom[24049] = 25'b1111110011010111001000110;
    rom[24050] = 25'b1111110011011000011010010;
    rom[24051] = 25'b1111110011011001101011110;
    rom[24052] = 25'b1111110011011010111101011;
    rom[24053] = 25'b1111110011011100001111001;
    rom[24054] = 25'b1111110011011101100000111;
    rom[24055] = 25'b1111110011011110110010111;
    rom[24056] = 25'b1111110011100000000100111;
    rom[24057] = 25'b1111110011100001010111001;
    rom[24058] = 25'b1111110011100010101001011;
    rom[24059] = 25'b1111110011100011111011110;
    rom[24060] = 25'b1111110011100101001110001;
    rom[24061] = 25'b1111110011100110100000110;
    rom[24062] = 25'b1111110011100111110011100;
    rom[24063] = 25'b1111110011101001000110010;
    rom[24064] = 25'b1111110011101010011001001;
    rom[24065] = 25'b1111110011101011101100001;
    rom[24066] = 25'b1111110011101100111111010;
    rom[24067] = 25'b1111110011101110010010100;
    rom[24068] = 25'b1111110011101111100101110;
    rom[24069] = 25'b1111110011110000111001010;
    rom[24070] = 25'b1111110011110010001100110;
    rom[24071] = 25'b1111110011110011100000011;
    rom[24072] = 25'b1111110011110100110100010;
    rom[24073] = 25'b1111110011110110001000001;
    rom[24074] = 25'b1111110011110111011100000;
    rom[24075] = 25'b1111110011111000110000001;
    rom[24076] = 25'b1111110011111010000100010;
    rom[24077] = 25'b1111110011111011011000100;
    rom[24078] = 25'b1111110011111100101101000;
    rom[24079] = 25'b1111110011111110000001100;
    rom[24080] = 25'b1111110011111111010110000;
    rom[24081] = 25'b1111110100000000101010110;
    rom[24082] = 25'b1111110100000001111111101;
    rom[24083] = 25'b1111110100000011010100100;
    rom[24084] = 25'b1111110100000100101001100;
    rom[24085] = 25'b1111110100000101111110101;
    rom[24086] = 25'b1111110100000111010011111;
    rom[24087] = 25'b1111110100001000101001001;
    rom[24088] = 25'b1111110100001001111110101;
    rom[24089] = 25'b1111110100001011010100001;
    rom[24090] = 25'b1111110100001100101001110;
    rom[24091] = 25'b1111110100001101111111101;
    rom[24092] = 25'b1111110100001111010101011;
    rom[24093] = 25'b1111110100010000101011011;
    rom[24094] = 25'b1111110100010010000001100;
    rom[24095] = 25'b1111110100010011010111101;
    rom[24096] = 25'b1111110100010100101101111;
    rom[24097] = 25'b1111110100010110000100010;
    rom[24098] = 25'b1111110100010111011010110;
    rom[24099] = 25'b1111110100011000110001011;
    rom[24100] = 25'b1111110100011010001000001;
    rom[24101] = 25'b1111110100011011011110111;
    rom[24102] = 25'b1111110100011100110101110;
    rom[24103] = 25'b1111110100011110001100110;
    rom[24104] = 25'b1111110100011111100011111;
    rom[24105] = 25'b1111110100100000111011001;
    rom[24106] = 25'b1111110100100010010010011;
    rom[24107] = 25'b1111110100100011101001111;
    rom[24108] = 25'b1111110100100101000001011;
    rom[24109] = 25'b1111110100100110011001000;
    rom[24110] = 25'b1111110100100111110000110;
    rom[24111] = 25'b1111110100101001001000101;
    rom[24112] = 25'b1111110100101010100000100;
    rom[24113] = 25'b1111110100101011111000100;
    rom[24114] = 25'b1111110100101101010000110;
    rom[24115] = 25'b1111110100101110101001000;
    rom[24116] = 25'b1111110100110000000001010;
    rom[24117] = 25'b1111110100110001011001110;
    rom[24118] = 25'b1111110100110010110010011;
    rom[24119] = 25'b1111110100110100001011000;
    rom[24120] = 25'b1111110100110101100011110;
    rom[24121] = 25'b1111110100110110111100101;
    rom[24122] = 25'b1111110100111000010101101;
    rom[24123] = 25'b1111110100111001101110101;
    rom[24124] = 25'b1111110100111011000111110;
    rom[24125] = 25'b1111110100111100100001000;
    rom[24126] = 25'b1111110100111101111010011;
    rom[24127] = 25'b1111110100111111010100000;
    rom[24128] = 25'b1111110101000000101101100;
    rom[24129] = 25'b1111110101000010000111010;
    rom[24130] = 25'b1111110101000011100001000;
    rom[24131] = 25'b1111110101000100111010111;
    rom[24132] = 25'b1111110101000110010100111;
    rom[24133] = 25'b1111110101000111101110111;
    rom[24134] = 25'b1111110101001001001001001;
    rom[24135] = 25'b1111110101001010100011100;
    rom[24136] = 25'b1111110101001011111101111;
    rom[24137] = 25'b1111110101001101011000011;
    rom[24138] = 25'b1111110101001110110010111;
    rom[24139] = 25'b1111110101010000001101101;
    rom[24140] = 25'b1111110101010001101000100;
    rom[24141] = 25'b1111110101010011000011011;
    rom[24142] = 25'b1111110101010100011110011;
    rom[24143] = 25'b1111110101010101111001011;
    rom[24144] = 25'b1111110101010111010100101;
    rom[24145] = 25'b1111110101011000110000000;
    rom[24146] = 25'b1111110101011010001011011;
    rom[24147] = 25'b1111110101011011100110111;
    rom[24148] = 25'b1111110101011101000010100;
    rom[24149] = 25'b1111110101011110011110001;
    rom[24150] = 25'b1111110101011111111010000;
    rom[24151] = 25'b1111110101100001010101111;
    rom[24152] = 25'b1111110101100010110010000;
    rom[24153] = 25'b1111110101100100001110000;
    rom[24154] = 25'b1111110101100101101010010;
    rom[24155] = 25'b1111110101100111000110100;
    rom[24156] = 25'b1111110101101000100010111;
    rom[24157] = 25'b1111110101101001111111100;
    rom[24158] = 25'b1111110101101011011100001;
    rom[24159] = 25'b1111110101101100111000110;
    rom[24160] = 25'b1111110101101110010101101;
    rom[24161] = 25'b1111110101101111110010100;
    rom[24162] = 25'b1111110101110001001111100;
    rom[24163] = 25'b1111110101110010101100101;
    rom[24164] = 25'b1111110101110100001001110;
    rom[24165] = 25'b1111110101110101100111001;
    rom[24166] = 25'b1111110101110111000100100;
    rom[24167] = 25'b1111110101111000100010000;
    rom[24168] = 25'b1111110101111001111111101;
    rom[24169] = 25'b1111110101111011011101010;
    rom[24170] = 25'b1111110101111100111011001;
    rom[24171] = 25'b1111110101111110011001000;
    rom[24172] = 25'b1111110101111111110111000;
    rom[24173] = 25'b1111110110000001010101001;
    rom[24174] = 25'b1111110110000010110011011;
    rom[24175] = 25'b1111110110000100010001100;
    rom[24176] = 25'b1111110110000101110000000;
    rom[24177] = 25'b1111110110000111001110100;
    rom[24178] = 25'b1111110110001000101101001;
    rom[24179] = 25'b1111110110001010001011110;
    rom[24180] = 25'b1111110110001011101010100;
    rom[24181] = 25'b1111110110001101001001011;
    rom[24182] = 25'b1111110110001110101000011;
    rom[24183] = 25'b1111110110010000000111100;
    rom[24184] = 25'b1111110110010001100110101;
    rom[24185] = 25'b1111110110010011000101111;
    rom[24186] = 25'b1111110110010100100101010;
    rom[24187] = 25'b1111110110010110000100101;
    rom[24188] = 25'b1111110110010111100100010;
    rom[24189] = 25'b1111110110011001000100000;
    rom[24190] = 25'b1111110110011010100011101;
    rom[24191] = 25'b1111110110011100000011101;
    rom[24192] = 25'b1111110110011101100011100;
    rom[24193] = 25'b1111110110011111000011101;
    rom[24194] = 25'b1111110110100000100011101;
    rom[24195] = 25'b1111110110100010000100000;
    rom[24196] = 25'b1111110110100011100100010;
    rom[24197] = 25'b1111110110100101000100110;
    rom[24198] = 25'b1111110110100110100101010;
    rom[24199] = 25'b1111110110101000000101111;
    rom[24200] = 25'b1111110110101001100110101;
    rom[24201] = 25'b1111110110101011000111011;
    rom[24202] = 25'b1111110110101100101000010;
    rom[24203] = 25'b1111110110101110001001010;
    rom[24204] = 25'b1111110110101111101010011;
    rom[24205] = 25'b1111110110110001001011101;
    rom[24206] = 25'b1111110110110010101100111;
    rom[24207] = 25'b1111110110110100001110011;
    rom[24208] = 25'b1111110110110101101111110;
    rom[24209] = 25'b1111110110110111010001011;
    rom[24210] = 25'b1111110110111000110011000;
    rom[24211] = 25'b1111110110111010010100110;
    rom[24212] = 25'b1111110110111011110110101;
    rom[24213] = 25'b1111110110111101011000101;
    rom[24214] = 25'b1111110110111110111010101;
    rom[24215] = 25'b1111110111000000011100111;
    rom[24216] = 25'b1111110111000001111111001;
    rom[24217] = 25'b1111110111000011100001100;
    rom[24218] = 25'b1111110111000101000011111;
    rom[24219] = 25'b1111110111000110100110100;
    rom[24220] = 25'b1111110111001000001001001;
    rom[24221] = 25'b1111110111001001101011110;
    rom[24222] = 25'b1111110111001011001110101;
    rom[24223] = 25'b1111110111001100110001100;
    rom[24224] = 25'b1111110111001110010100100;
    rom[24225] = 25'b1111110111001111110111100;
    rom[24226] = 25'b1111110111010001011010111;
    rom[24227] = 25'b1111110111010010111110001;
    rom[24228] = 25'b1111110111010100100001100;
    rom[24229] = 25'b1111110111010110000100111;
    rom[24230] = 25'b1111110111010111101000100;
    rom[24231] = 25'b1111110111011001001100001;
    rom[24232] = 25'b1111110111011010101111111;
    rom[24233] = 25'b1111110111011100010011110;
    rom[24234] = 25'b1111110111011101110111110;
    rom[24235] = 25'b1111110111011111011011110;
    rom[24236] = 25'b1111110111100000111111111;
    rom[24237] = 25'b1111110111100010100100000;
    rom[24238] = 25'b1111110111100100001000011;
    rom[24239] = 25'b1111110111100101101100110;
    rom[24240] = 25'b1111110111100111010001010;
    rom[24241] = 25'b1111110111101000110101111;
    rom[24242] = 25'b1111110111101010011010100;
    rom[24243] = 25'b1111110111101011111111010;
    rom[24244] = 25'b1111110111101101100100001;
    rom[24245] = 25'b1111110111101111001001001;
    rom[24246] = 25'b1111110111110000101110001;
    rom[24247] = 25'b1111110111110010010011010;
    rom[24248] = 25'b1111110111110011111000100;
    rom[24249] = 25'b1111110111110101011101111;
    rom[24250] = 25'b1111110111110111000011010;
    rom[24251] = 25'b1111110111111000101000110;
    rom[24252] = 25'b1111110111111010001110011;
    rom[24253] = 25'b1111110111111011110100001;
    rom[24254] = 25'b1111110111111101011001110;
    rom[24255] = 25'b1111110111111110111111101;
    rom[24256] = 25'b1111111000000000100101101;
    rom[24257] = 25'b1111111000000010001011110;
    rom[24258] = 25'b1111111000000011110001111;
    rom[24259] = 25'b1111111000000101011000000;
    rom[24260] = 25'b1111111000000110111110011;
    rom[24261] = 25'b1111111000001000100100111;
    rom[24262] = 25'b1111111000001010001011010;
    rom[24263] = 25'b1111111000001011110001111;
    rom[24264] = 25'b1111111000001101011000101;
    rom[24265] = 25'b1111111000001110111111011;
    rom[24266] = 25'b1111111000010000100110010;
    rom[24267] = 25'b1111111000010010001101010;
    rom[24268] = 25'b1111111000010011110100010;
    rom[24269] = 25'b1111111000010101011011011;
    rom[24270] = 25'b1111111000010111000010101;
    rom[24271] = 25'b1111111000011000101001111;
    rom[24272] = 25'b1111111000011010010001011;
    rom[24273] = 25'b1111111000011011111000111;
    rom[24274] = 25'b1111111000011101100000011;
    rom[24275] = 25'b1111111000011111001000000;
    rom[24276] = 25'b1111111000100000101111110;
    rom[24277] = 25'b1111111000100010010111101;
    rom[24278] = 25'b1111111000100011111111101;
    rom[24279] = 25'b1111111000100101100111101;
    rom[24280] = 25'b1111111000100111001111110;
    rom[24281] = 25'b1111111000101000111000000;
    rom[24282] = 25'b1111111000101010100000010;
    rom[24283] = 25'b1111111000101100001000101;
    rom[24284] = 25'b1111111000101101110001001;
    rom[24285] = 25'b1111111000101111011001110;
    rom[24286] = 25'b1111111000110001000010010;
    rom[24287] = 25'b1111111000110010101011001;
    rom[24288] = 25'b1111111000110100010011111;
    rom[24289] = 25'b1111111000110101111100110;
    rom[24290] = 25'b1111111000110111100101110;
    rom[24291] = 25'b1111111000111001001110111;
    rom[24292] = 25'b1111111000111010111000000;
    rom[24293] = 25'b1111111000111100100001010;
    rom[24294] = 25'b1111111000111110001010101;
    rom[24295] = 25'b1111111000111111110100000;
    rom[24296] = 25'b1111111001000001011101100;
    rom[24297] = 25'b1111111001000011000111001;
    rom[24298] = 25'b1111111001000100110000111;
    rom[24299] = 25'b1111111001000110011010101;
    rom[24300] = 25'b1111111001001000000100100;
    rom[24301] = 25'b1111111001001001101110100;
    rom[24302] = 25'b1111111001001011011000100;
    rom[24303] = 25'b1111111001001101000010101;
    rom[24304] = 25'b1111111001001110101100111;
    rom[24305] = 25'b1111111001010000010111001;
    rom[24306] = 25'b1111111001010010000001100;
    rom[24307] = 25'b1111111001010011101100000;
    rom[24308] = 25'b1111111001010101010110100;
    rom[24309] = 25'b1111111001010111000001001;
    rom[24310] = 25'b1111111001011000101011111;
    rom[24311] = 25'b1111111001011010010110110;
    rom[24312] = 25'b1111111001011100000001101;
    rom[24313] = 25'b1111111001011101101100101;
    rom[24314] = 25'b1111111001011111010111101;
    rom[24315] = 25'b1111111001100001000010111;
    rom[24316] = 25'b1111111001100010101110000;
    rom[24317] = 25'b1111111001100100011001011;
    rom[24318] = 25'b1111111001100110000100110;
    rom[24319] = 25'b1111111001100111110000010;
    rom[24320] = 25'b1111111001101001011011110;
    rom[24321] = 25'b1111111001101011000111100;
    rom[24322] = 25'b1111111001101100110011010;
    rom[24323] = 25'b1111111001101110011111000;
    rom[24324] = 25'b1111111001110000001011000;
    rom[24325] = 25'b1111111001110001110110111;
    rom[24326] = 25'b1111111001110011100011000;
    rom[24327] = 25'b1111111001110101001111010;
    rom[24328] = 25'b1111111001110110111011011;
    rom[24329] = 25'b1111111001111000100111110;
    rom[24330] = 25'b1111111001111010010100001;
    rom[24331] = 25'b1111111001111100000000101;
    rom[24332] = 25'b1111111001111101101101010;
    rom[24333] = 25'b1111111001111111011001111;
    rom[24334] = 25'b1111111010000001000110101;
    rom[24335] = 25'b1111111010000010110011011;
    rom[24336] = 25'b1111111010000100100000010;
    rom[24337] = 25'b1111111010000110001101011;
    rom[24338] = 25'b1111111010000111111010100;
    rom[24339] = 25'b1111111010001001100111100;
    rom[24340] = 25'b1111111010001011010100110;
    rom[24341] = 25'b1111111010001101000010001;
    rom[24342] = 25'b1111111010001110101111100;
    rom[24343] = 25'b1111111010010000011101000;
    rom[24344] = 25'b1111111010010010001010101;
    rom[24345] = 25'b1111111010010011111000010;
    rom[24346] = 25'b1111111010010101100110000;
    rom[24347] = 25'b1111111010010111010011110;
    rom[24348] = 25'b1111111010011001000001101;
    rom[24349] = 25'b1111111010011010101111101;
    rom[24350] = 25'b1111111010011100011101110;
    rom[24351] = 25'b1111111010011110001011111;
    rom[24352] = 25'b1111111010011111111010000;
    rom[24353] = 25'b1111111010100001101000011;
    rom[24354] = 25'b1111111010100011010110110;
    rom[24355] = 25'b1111111010100101000101001;
    rom[24356] = 25'b1111111010100110110011101;
    rom[24357] = 25'b1111111010101000100010011;
    rom[24358] = 25'b1111111010101010010001000;
    rom[24359] = 25'b1111111010101011111111111;
    rom[24360] = 25'b1111111010101101101110101;
    rom[24361] = 25'b1111111010101111011101101;
    rom[24362] = 25'b1111111010110001001100101;
    rom[24363] = 25'b1111111010110010111011110;
    rom[24364] = 25'b1111111010110100101010111;
    rom[24365] = 25'b1111111010110110011010001;
    rom[24366] = 25'b1111111010111000001001100;
    rom[24367] = 25'b1111111010111001111000111;
    rom[24368] = 25'b1111111010111011101000011;
    rom[24369] = 25'b1111111010111101011000000;
    rom[24370] = 25'b1111111010111111000111101;
    rom[24371] = 25'b1111111011000000110111011;
    rom[24372] = 25'b1111111011000010100111001;
    rom[24373] = 25'b1111111011000100010111000;
    rom[24374] = 25'b1111111011000110000111000;
    rom[24375] = 25'b1111111011000111110111000;
    rom[24376] = 25'b1111111011001001100111001;
    rom[24377] = 25'b1111111011001011010111011;
    rom[24378] = 25'b1111111011001101000111101;
    rom[24379] = 25'b1111111011001110111000000;
    rom[24380] = 25'b1111111011010000101000011;
    rom[24381] = 25'b1111111011010010011000111;
    rom[24382] = 25'b1111111011010100001001100;
    rom[24383] = 25'b1111111011010101111010001;
    rom[24384] = 25'b1111111011010111101010111;
    rom[24385] = 25'b1111111011011001011011110;
    rom[24386] = 25'b1111111011011011001100101;
    rom[24387] = 25'b1111111011011100111101101;
    rom[24388] = 25'b1111111011011110101110101;
    rom[24389] = 25'b1111111011100000011111110;
    rom[24390] = 25'b1111111011100010010001000;
    rom[24391] = 25'b1111111011100100000010010;
    rom[24392] = 25'b1111111011100101110011100;
    rom[24393] = 25'b1111111011100111100101000;
    rom[24394] = 25'b1111111011101001010110101;
    rom[24395] = 25'b1111111011101011001000001;
    rom[24396] = 25'b1111111011101100111001110;
    rom[24397] = 25'b1111111011101110101011100;
    rom[24398] = 25'b1111111011110000011101010;
    rom[24399] = 25'b1111111011110010001111010;
    rom[24400] = 25'b1111111011110100000001001;
    rom[24401] = 25'b1111111011110101110011001;
    rom[24402] = 25'b1111111011110111100101010;
    rom[24403] = 25'b1111111011111001010111100;
    rom[24404] = 25'b1111111011111011001001110;
    rom[24405] = 25'b1111111011111100111100001;
    rom[24406] = 25'b1111111011111110101110100;
    rom[24407] = 25'b1111111100000000100001000;
    rom[24408] = 25'b1111111100000010010011100;
    rom[24409] = 25'b1111111100000100000110001;
    rom[24410] = 25'b1111111100000101111000111;
    rom[24411] = 25'b1111111100000111101011101;
    rom[24412] = 25'b1111111100001001011110100;
    rom[24413] = 25'b1111111100001011010001011;
    rom[24414] = 25'b1111111100001101000100011;
    rom[24415] = 25'b1111111100001110110111100;
    rom[24416] = 25'b1111111100010000101010101;
    rom[24417] = 25'b1111111100010010011101111;
    rom[24418] = 25'b1111111100010100010001001;
    rom[24419] = 25'b1111111100010110000100100;
    rom[24420] = 25'b1111111100010111110111111;
    rom[24421] = 25'b1111111100011001101011100;
    rom[24422] = 25'b1111111100011011011111000;
    rom[24423] = 25'b1111111100011101010010101;
    rom[24424] = 25'b1111111100011111000110011;
    rom[24425] = 25'b1111111100100000111010001;
    rom[24426] = 25'b1111111100100010101110001;
    rom[24427] = 25'b1111111100100100100010000;
    rom[24428] = 25'b1111111100100110010110000;
    rom[24429] = 25'b1111111100101000001010001;
    rom[24430] = 25'b1111111100101001111110010;
    rom[24431] = 25'b1111111100101011110010100;
    rom[24432] = 25'b1111111100101101100110111;
    rom[24433] = 25'b1111111100101111011011010;
    rom[24434] = 25'b1111111100110001001111101;
    rom[24435] = 25'b1111111100110011000100001;
    rom[24436] = 25'b1111111100110100111000110;
    rom[24437] = 25'b1111111100110110101101011;
    rom[24438] = 25'b1111111100111000100010001;
    rom[24439] = 25'b1111111100111010010110111;
    rom[24440] = 25'b1111111100111100001011110;
    rom[24441] = 25'b1111111100111110000000110;
    rom[24442] = 25'b1111111100111111110101110;
    rom[24443] = 25'b1111111101000001101010111;
    rom[24444] = 25'b1111111101000011011111111;
    rom[24445] = 25'b1111111101000101010101001;
    rom[24446] = 25'b1111111101000111001010011;
    rom[24447] = 25'b1111111101001000111111110;
    rom[24448] = 25'b1111111101001010110101010;
    rom[24449] = 25'b1111111101001100101010101;
    rom[24450] = 25'b1111111101001110100000010;
    rom[24451] = 25'b1111111101010000010101111;
    rom[24452] = 25'b1111111101010010001011101;
    rom[24453] = 25'b1111111101010100000001011;
    rom[24454] = 25'b1111111101010101110111010;
    rom[24455] = 25'b1111111101010111101101000;
    rom[24456] = 25'b1111111101011001100011001;
    rom[24457] = 25'b1111111101011011011001001;
    rom[24458] = 25'b1111111101011101001111001;
    rom[24459] = 25'b1111111101011111000101011;
    rom[24460] = 25'b1111111101100000111011101;
    rom[24461] = 25'b1111111101100010110010000;
    rom[24462] = 25'b1111111101100100101000011;
    rom[24463] = 25'b1111111101100110011110110;
    rom[24464] = 25'b1111111101101000010101010;
    rom[24465] = 25'b1111111101101010001011111;
    rom[24466] = 25'b1111111101101100000010100;
    rom[24467] = 25'b1111111101101101111001010;
    rom[24468] = 25'b1111111101101111110000000;
    rom[24469] = 25'b1111111101110001100110111;
    rom[24470] = 25'b1111111101110011011101110;
    rom[24471] = 25'b1111111101110101010100110;
    rom[24472] = 25'b1111111101110111001011110;
    rom[24473] = 25'b1111111101111001000011000;
    rom[24474] = 25'b1111111101111010111010001;
    rom[24475] = 25'b1111111101111100110001011;
    rom[24476] = 25'b1111111101111110101000101;
    rom[24477] = 25'b1111111110000000100000000;
    rom[24478] = 25'b1111111110000010010111100;
    rom[24479] = 25'b1111111110000100001111000;
    rom[24480] = 25'b1111111110000110000110101;
    rom[24481] = 25'b1111111110000111111110010;
    rom[24482] = 25'b1111111110001001110101111;
    rom[24483] = 25'b1111111110001011101101101;
    rom[24484] = 25'b1111111110001101100101100;
    rom[24485] = 25'b1111111110001111011101011;
    rom[24486] = 25'b1111111110010001010101010;
    rom[24487] = 25'b1111111110010011001101011;
    rom[24488] = 25'b1111111110010101000101100;
    rom[24489] = 25'b1111111110010110111101101;
    rom[24490] = 25'b1111111110011000110101110;
    rom[24491] = 25'b1111111110011010101110000;
    rom[24492] = 25'b1111111110011100100110011;
    rom[24493] = 25'b1111111110011110011110110;
    rom[24494] = 25'b1111111110100000010111010;
    rom[24495] = 25'b1111111110100010001111111;
    rom[24496] = 25'b1111111110100100001000011;
    rom[24497] = 25'b1111111110100110000001000;
    rom[24498] = 25'b1111111110100111111001110;
    rom[24499] = 25'b1111111110101001110010100;
    rom[24500] = 25'b1111111110101011101011011;
    rom[24501] = 25'b1111111110101101100100011;
    rom[24502] = 25'b1111111110101111011101010;
    rom[24503] = 25'b1111111110110001010110010;
    rom[24504] = 25'b1111111110110011001111011;
    rom[24505] = 25'b1111111110110101001000100;
    rom[24506] = 25'b1111111110110111000001110;
    rom[24507] = 25'b1111111110111000111011000;
    rom[24508] = 25'b1111111110111010110100011;
    rom[24509] = 25'b1111111110111100101101110;
    rom[24510] = 25'b1111111110111110100111010;
    rom[24511] = 25'b1111111111000000100000110;
    rom[24512] = 25'b1111111111000010011010011;
    rom[24513] = 25'b1111111111000100010100000;
    rom[24514] = 25'b1111111111000110001101110;
    rom[24515] = 25'b1111111111001000000111011;
    rom[24516] = 25'b1111111111001010000001010;
    rom[24517] = 25'b1111111111001011111011001;
    rom[24518] = 25'b1111111111001101110101001;
    rom[24519] = 25'b1111111111001111101111001;
    rom[24520] = 25'b1111111111010001101001001;
    rom[24521] = 25'b1111111111010011100011010;
    rom[24522] = 25'b1111111111010101011101011;
    rom[24523] = 25'b1111111111010111010111101;
    rom[24524] = 25'b1111111111011001010010000;
    rom[24525] = 25'b1111111111011011001100011;
    rom[24526] = 25'b1111111111011101000110110;
    rom[24527] = 25'b1111111111011111000001010;
    rom[24528] = 25'b1111111111100000111011111;
    rom[24529] = 25'b1111111111100010110110011;
    rom[24530] = 25'b1111111111100100110001000;
    rom[24531] = 25'b1111111111100110101011110;
    rom[24532] = 25'b1111111111101000100110100;
    rom[24533] = 25'b1111111111101010100001010;
    rom[24534] = 25'b1111111111101100011100001;
    rom[24535] = 25'b1111111111101110010111001;
    rom[24536] = 25'b1111111111110000010010001;
    rom[24537] = 25'b1111111111110010001101001;
    rom[24538] = 25'b1111111111110100001000011;
    rom[24539] = 25'b1111111111110110000011100;
    rom[24540] = 25'b1111111111110111111110101;
    rom[24541] = 25'b1111111111111001111010000;
    rom[24542] = 25'b1111111111111011110101011;
    rom[24543] = 25'b1111111111111101110000101;
    rom[24544] = 25'b1111111111111111101100001;
    rom[24545] = 25'b0000000000000001100111101;
    rom[24546] = 25'b0000000000000011100011001;
    rom[24547] = 25'b0000000000000101011110110;
    rom[24548] = 25'b0000000000000111011010011;
    rom[24549] = 25'b0000000000001001010110001;
    rom[24550] = 25'b0000000000001011010001111;
    rom[24551] = 25'b0000000000001101001101110;
    rom[24552] = 25'b0000000000001111001001101;
    rom[24553] = 25'b0000000000010001000101101;
    rom[24554] = 25'b0000000000010011000001101;
    rom[24555] = 25'b0000000000010100111101110;
    rom[24556] = 25'b0000000000010110111001111;
    rom[24557] = 25'b0000000000011000110110000;
    rom[24558] = 25'b0000000000011010110010010;
    rom[24559] = 25'b0000000000011100101110100;
    rom[24560] = 25'b0000000000011110101010111;
    rom[24561] = 25'b0000000000100000100111010;
    rom[24562] = 25'b0000000000100010100011101;
    rom[24563] = 25'b0000000000100100100000001;
    rom[24564] = 25'b0000000000100110011100101;
    rom[24565] = 25'b0000000000101000011001010;
    rom[24566] = 25'b0000000000101010010101111;
    rom[24567] = 25'b0000000000101100010010101;
    rom[24568] = 25'b0000000000101110001111011;
    rom[24569] = 25'b0000000000110000001100010;
    rom[24570] = 25'b0000000000110010001001001;
    rom[24571] = 25'b0000000000110100000110000;
    rom[24572] = 25'b0000000000110110000010111;
    rom[24573] = 25'b0000000000111000000000000;
    rom[24574] = 25'b0000000000111001111101000;
    rom[24575] = 25'b0000000000111011111010001;
    rom[24576] = 25'b0000000000111101110111011;
    rom[24577] = 25'b0000000000111111110100100;
    rom[24578] = 25'b0000000001000001110001111;
    rom[24579] = 25'b0000000001000011101111001;
    rom[24580] = 25'b0000000001000101101100101;
    rom[24581] = 25'b0000000001000111101010000;
    rom[24582] = 25'b0000000001001001100111011;
    rom[24583] = 25'b0000000001001011100101000;
    rom[24584] = 25'b0000000001001101100010100;
    rom[24585] = 25'b0000000001001111100000010;
    rom[24586] = 25'b0000000001010001011101111;
    rom[24587] = 25'b0000000001010011011011101;
    rom[24588] = 25'b0000000001010101011001011;
    rom[24589] = 25'b0000000001010111010111010;
    rom[24590] = 25'b0000000001011001010101001;
    rom[24591] = 25'b0000000001011011010011001;
    rom[24592] = 25'b0000000001011101010001000;
    rom[24593] = 25'b0000000001011111001111000;
    rom[24594] = 25'b0000000001100001001101001;
    rom[24595] = 25'b0000000001100011001011010;
    rom[24596] = 25'b0000000001100101001001011;
    rom[24597] = 25'b0000000001100111000111101;
    rom[24598] = 25'b0000000001101001000110000;
    rom[24599] = 25'b0000000001101011000100010;
    rom[24600] = 25'b0000000001101101000010101;
    rom[24601] = 25'b0000000001101111000001000;
    rom[24602] = 25'b0000000001110000111111100;
    rom[24603] = 25'b0000000001110010111110000;
    rom[24604] = 25'b0000000001110100111100100;
    rom[24605] = 25'b0000000001110110111011001;
    rom[24606] = 25'b0000000001111000111001110;
    rom[24607] = 25'b0000000001111010111000100;
    rom[24608] = 25'b0000000001111100110111010;
    rom[24609] = 25'b0000000001111110110110001;
    rom[24610] = 25'b0000000010000000110100111;
    rom[24611] = 25'b0000000010000010110011110;
    rom[24612] = 25'b0000000010000100110010110;
    rom[24613] = 25'b0000000010000110110001110;
    rom[24614] = 25'b0000000010001000110000110;
    rom[24615] = 25'b0000000010001010101111111;
    rom[24616] = 25'b0000000010001100101110111;
    rom[24617] = 25'b0000000010001110101110001;
    rom[24618] = 25'b0000000010010000101101011;
    rom[24619] = 25'b0000000010010010101100100;
    rom[24620] = 25'b0000000010010100101011111;
    rom[24621] = 25'b0000000010010110101011001;
    rom[24622] = 25'b0000000010011000101010100;
    rom[24623] = 25'b0000000010011010101010000;
    rom[24624] = 25'b0000000010011100101001100;
    rom[24625] = 25'b0000000010011110101001000;
    rom[24626] = 25'b0000000010100000101000100;
    rom[24627] = 25'b0000000010100010101000010;
    rom[24628] = 25'b0000000010100100100111111;
    rom[24629] = 25'b0000000010100110100111100;
    rom[24630] = 25'b0000000010101000100111010;
    rom[24631] = 25'b0000000010101010100111000;
    rom[24632] = 25'b0000000010101100100110111;
    rom[24633] = 25'b0000000010101110100110110;
    rom[24634] = 25'b0000000010110000100110101;
    rom[24635] = 25'b0000000010110010100110101;
    rom[24636] = 25'b0000000010110100100110101;
    rom[24637] = 25'b0000000010110110100110101;
    rom[24638] = 25'b0000000010111000100110110;
    rom[24639] = 25'b0000000010111010100110111;
    rom[24640] = 25'b0000000010111100100111000;
    rom[24641] = 25'b0000000010111110100111010;
    rom[24642] = 25'b0000000011000000100111100;
    rom[24643] = 25'b0000000011000010100111110;
    rom[24644] = 25'b0000000011000100101000001;
    rom[24645] = 25'b0000000011000110101000100;
    rom[24646] = 25'b0000000011001000101000111;
    rom[24647] = 25'b0000000011001010101001011;
    rom[24648] = 25'b0000000011001100101001111;
    rom[24649] = 25'b0000000011001110101010011;
    rom[24650] = 25'b0000000011010000101010111;
    rom[24651] = 25'b0000000011010010101011101;
    rom[24652] = 25'b0000000011010100101100010;
    rom[24653] = 25'b0000000011010110101101000;
    rom[24654] = 25'b0000000011011000101101101;
    rom[24655] = 25'b0000000011011010101110100;
    rom[24656] = 25'b0000000011011100101111010;
    rom[24657] = 25'b0000000011011110110000001;
    rom[24658] = 25'b0000000011100000110001001;
    rom[24659] = 25'b0000000011100010110010000;
    rom[24660] = 25'b0000000011100100110010111;
    rom[24661] = 25'b0000000011100110110100000;
    rom[24662] = 25'b0000000011101000110101000;
    rom[24663] = 25'b0000000011101010110110001;
    rom[24664] = 25'b0000000011101100110111010;
    rom[24665] = 25'b0000000011101110111000011;
    rom[24666] = 25'b0000000011110000111001101;
    rom[24667] = 25'b0000000011110010111010111;
    rom[24668] = 25'b0000000011110100111100001;
    rom[24669] = 25'b0000000011110110111101011;
    rom[24670] = 25'b0000000011111000111110110;
    rom[24671] = 25'b0000000011111011000000001;
    rom[24672] = 25'b0000000011111101000001101;
    rom[24673] = 25'b0000000011111111000011000;
    rom[24674] = 25'b0000000100000001000100101;
    rom[24675] = 25'b0000000100000011000110001;
    rom[24676] = 25'b0000000100000101000111110;
    rom[24677] = 25'b0000000100000111001001010;
    rom[24678] = 25'b0000000100001001001011000;
    rom[24679] = 25'b0000000100001011001100101;
    rom[24680] = 25'b0000000100001101001110010;
    rom[24681] = 25'b0000000100001111010000001;
    rom[24682] = 25'b0000000100010001010001111;
    rom[24683] = 25'b0000000100010011010011110;
    rom[24684] = 25'b0000000100010101010101100;
    rom[24685] = 25'b0000000100010111010111100;
    rom[24686] = 25'b0000000100011001011001011;
    rom[24687] = 25'b0000000100011011011011011;
    rom[24688] = 25'b0000000100011101011101011;
    rom[24689] = 25'b0000000100011111011111011;
    rom[24690] = 25'b0000000100100001100001011;
    rom[24691] = 25'b0000000100100011100011100;
    rom[24692] = 25'b0000000100100101100101101;
    rom[24693] = 25'b0000000100100111100111111;
    rom[24694] = 25'b0000000100101001101010000;
    rom[24695] = 25'b0000000100101011101100010;
    rom[24696] = 25'b0000000100101101101110100;
    rom[24697] = 25'b0000000100101111110000111;
    rom[24698] = 25'b0000000100110001110011001;
    rom[24699] = 25'b0000000100110011110101100;
    rom[24700] = 25'b0000000100110101111000000;
    rom[24701] = 25'b0000000100110111111010011;
    rom[24702] = 25'b0000000100111001111100110;
    rom[24703] = 25'b0000000100111011111111010;
    rom[24704] = 25'b0000000100111110000001111;
    rom[24705] = 25'b0000000101000000000100011;
    rom[24706] = 25'b0000000101000010000111000;
    rom[24707] = 25'b0000000101000100001001101;
    rom[24708] = 25'b0000000101000110001100010;
    rom[24709] = 25'b0000000101001000001111000;
    rom[24710] = 25'b0000000101001010010001101;
    rom[24711] = 25'b0000000101001100010100011;
    rom[24712] = 25'b0000000101001110010111010;
    rom[24713] = 25'b0000000101010000011010000;
    rom[24714] = 25'b0000000101010010011100110;
    rom[24715] = 25'b0000000101010100011111110;
    rom[24716] = 25'b0000000101010110100010100;
    rom[24717] = 25'b0000000101011000100101100;
    rom[24718] = 25'b0000000101011010101000011;
    rom[24719] = 25'b0000000101011100101011011;
    rom[24720] = 25'b0000000101011110101110100;
    rom[24721] = 25'b0000000101100000110001100;
    rom[24722] = 25'b0000000101100010110100101;
    rom[24723] = 25'b0000000101100100110111101;
    rom[24724] = 25'b0000000101100110111010110;
    rom[24725] = 25'b0000000101101000111101111;
    rom[24726] = 25'b0000000101101011000001001;
    rom[24727] = 25'b0000000101101101000100011;
    rom[24728] = 25'b0000000101101111000111100;
    rom[24729] = 25'b0000000101110001001010111;
    rom[24730] = 25'b0000000101110011001110001;
    rom[24731] = 25'b0000000101110101010001100;
    rom[24732] = 25'b0000000101110111010100110;
    rom[24733] = 25'b0000000101111001011000001;
    rom[24734] = 25'b0000000101111011011011100;
    rom[24735] = 25'b0000000101111101011111000;
    rom[24736] = 25'b0000000101111111100010011;
    rom[24737] = 25'b0000000110000001100101111;
    rom[24738] = 25'b0000000110000011101001011;
    rom[24739] = 25'b0000000110000101101101000;
    rom[24740] = 25'b0000000110000111110000101;
    rom[24741] = 25'b0000000110001001110100001;
    rom[24742] = 25'b0000000110001011110111110;
    rom[24743] = 25'b0000000110001101111011011;
    rom[24744] = 25'b0000000110001111111111001;
    rom[24745] = 25'b0000000110010010000010110;
    rom[24746] = 25'b0000000110010100000110100;
    rom[24747] = 25'b0000000110010110001010010;
    rom[24748] = 25'b0000000110011000001110000;
    rom[24749] = 25'b0000000110011010010001110;
    rom[24750] = 25'b0000000110011100010101100;
    rom[24751] = 25'b0000000110011110011001011;
    rom[24752] = 25'b0000000110100000011101010;
    rom[24753] = 25'b0000000110100010100001001;
    rom[24754] = 25'b0000000110100100100101001;
    rom[24755] = 25'b0000000110100110101000111;
    rom[24756] = 25'b0000000110101000101100111;
    rom[24757] = 25'b0000000110101010110000111;
    rom[24758] = 25'b0000000110101100110100111;
    rom[24759] = 25'b0000000110101110111000111;
    rom[24760] = 25'b0000000110110000111101000;
    rom[24761] = 25'b0000000110110011000001000;
    rom[24762] = 25'b0000000110110101000101001;
    rom[24763] = 25'b0000000110110111001001010;
    rom[24764] = 25'b0000000110111001001101011;
    rom[24765] = 25'b0000000110111011010001100;
    rom[24766] = 25'b0000000110111101010101101;
    rom[24767] = 25'b0000000110111111011001111;
    rom[24768] = 25'b0000000111000001011110000;
    rom[24769] = 25'b0000000111000011100010010;
    rom[24770] = 25'b0000000111000101100110101;
    rom[24771] = 25'b0000000111000111101010111;
    rom[24772] = 25'b0000000111001001101111001;
    rom[24773] = 25'b0000000111001011110011100;
    rom[24774] = 25'b0000000111001101110111111;
    rom[24775] = 25'b0000000111001111111100001;
    rom[24776] = 25'b0000000111010010000000101;
    rom[24777] = 25'b0000000111010100000101000;
    rom[24778] = 25'b0000000111010110001001011;
    rom[24779] = 25'b0000000111011000001101111;
    rom[24780] = 25'b0000000111011010010010010;
    rom[24781] = 25'b0000000111011100010110110;
    rom[24782] = 25'b0000000111011110011011010;
    rom[24783] = 25'b0000000111100000011111110;
    rom[24784] = 25'b0000000111100010100100011;
    rom[24785] = 25'b0000000111100100101000111;
    rom[24786] = 25'b0000000111100110101101100;
    rom[24787] = 25'b0000000111101000110010000;
    rom[24788] = 25'b0000000111101010110110101;
    rom[24789] = 25'b0000000111101100111011010;
    rom[24790] = 25'b0000000111101110111111111;
    rom[24791] = 25'b0000000111110001000100100;
    rom[24792] = 25'b0000000111110011001001010;
    rom[24793] = 25'b0000000111110101001101111;
    rom[24794] = 25'b0000000111110111010010101;
    rom[24795] = 25'b0000000111111001010111011;
    rom[24796] = 25'b0000000111111011011100000;
    rom[24797] = 25'b0000000111111101100000111;
    rom[24798] = 25'b0000000111111111100101101;
    rom[24799] = 25'b0000001000000001101010011;
    rom[24800] = 25'b0000001000000011101111010;
    rom[24801] = 25'b0000001000000101110100000;
    rom[24802] = 25'b0000001000000111111000110;
    rom[24803] = 25'b0000001000001001111101110;
    rom[24804] = 25'b0000001000001100000010101;
    rom[24805] = 25'b0000001000001110000111100;
    rom[24806] = 25'b0000001000010000001100011;
    rom[24807] = 25'b0000001000010010010001010;
    rom[24808] = 25'b0000001000010100010110001;
    rom[24809] = 25'b0000001000010110011011001;
    rom[24810] = 25'b0000001000011000100000000;
    rom[24811] = 25'b0000001000011010100101000;
    rom[24812] = 25'b0000001000011100101010000;
    rom[24813] = 25'b0000001000011110101111000;
    rom[24814] = 25'b0000001000100000110100000;
    rom[24815] = 25'b0000001000100010111001000;
    rom[24816] = 25'b0000001000100100111110000;
    rom[24817] = 25'b0000001000100111000011001;
    rom[24818] = 25'b0000001000101001001000001;
    rom[24819] = 25'b0000001000101011001101010;
    rom[24820] = 25'b0000001000101101010010010;
    rom[24821] = 25'b0000001000101111010111011;
    rom[24822] = 25'b0000001000110001011100100;
    rom[24823] = 25'b0000001000110011100001101;
    rom[24824] = 25'b0000001000110101100110110;
    rom[24825] = 25'b0000001000110111101011111;
    rom[24826] = 25'b0000001000111001110001000;
    rom[24827] = 25'b0000001000111011110110010;
    rom[24828] = 25'b0000001000111101111011011;
    rom[24829] = 25'b0000001001000000000000100;
    rom[24830] = 25'b0000001001000010000101110;
    rom[24831] = 25'b0000001001000100001011000;
    rom[24832] = 25'b0000001001000110010000001;
    rom[24833] = 25'b0000001001001000010101011;
    rom[24834] = 25'b0000001001001010011010101;
    rom[24835] = 25'b0000001001001100011111111;
    rom[24836] = 25'b0000001001001110100101001;
    rom[24837] = 25'b0000001001010000101010011;
    rom[24838] = 25'b0000001001010010101111101;
    rom[24839] = 25'b0000001001010100110100111;
    rom[24840] = 25'b0000001001010110111010001;
    rom[24841] = 25'b0000001001011000111111100;
    rom[24842] = 25'b0000001001011011000100110;
    rom[24843] = 25'b0000001001011101001010001;
    rom[24844] = 25'b0000001001011111001111011;
    rom[24845] = 25'b0000001001100001010100110;
    rom[24846] = 25'b0000001001100011011010001;
    rom[24847] = 25'b0000001001100101011111100;
    rom[24848] = 25'b0000001001100111100100111;
    rom[24849] = 25'b0000001001101001101010010;
    rom[24850] = 25'b0000001001101011101111100;
    rom[24851] = 25'b0000001001101101110100111;
    rom[24852] = 25'b0000001001101111111010010;
    rom[24853] = 25'b0000001001110001111111110;
    rom[24854] = 25'b0000001001110100000101001;
    rom[24855] = 25'b0000001001110110001010011;
    rom[24856] = 25'b0000001001111000001111111;
    rom[24857] = 25'b0000001001111010010101011;
    rom[24858] = 25'b0000001001111100011010101;
    rom[24859] = 25'b0000001001111110100000001;
    rom[24860] = 25'b0000001010000000100101101;
    rom[24861] = 25'b0000001010000010101011000;
    rom[24862] = 25'b0000001010000100110000011;
    rom[24863] = 25'b0000001010000110110101111;
    rom[24864] = 25'b0000001010001000111011010;
    rom[24865] = 25'b0000001010001011000000110;
    rom[24866] = 25'b0000001010001101000110010;
    rom[24867] = 25'b0000001010001111001011101;
    rom[24868] = 25'b0000001010010001010001001;
    rom[24869] = 25'b0000001010010011010110100;
    rom[24870] = 25'b0000001010010101011100000;
    rom[24871] = 25'b0000001010010111100001100;
    rom[24872] = 25'b0000001010011001100111000;
    rom[24873] = 25'b0000001010011011101100011;
    rom[24874] = 25'b0000001010011101110010000;
    rom[24875] = 25'b0000001010011111110111011;
    rom[24876] = 25'b0000001010100001111100111;
    rom[24877] = 25'b0000001010100100000010011;
    rom[24878] = 25'b0000001010100110000111111;
    rom[24879] = 25'b0000001010101000001101011;
    rom[24880] = 25'b0000001010101010010010111;
    rom[24881] = 25'b0000001010101100011000011;
    rom[24882] = 25'b0000001010101110011101111;
    rom[24883] = 25'b0000001010110000100011010;
    rom[24884] = 25'b0000001010110010101000111;
    rom[24885] = 25'b0000001010110100101110010;
    rom[24886] = 25'b0000001010110110110011111;
    rom[24887] = 25'b0000001010111000111001010;
    rom[24888] = 25'b0000001010111010111110111;
    rom[24889] = 25'b0000001010111101000100010;
    rom[24890] = 25'b0000001010111111001001111;
    rom[24891] = 25'b0000001011000001001111010;
    rom[24892] = 25'b0000001011000011010100111;
    rom[24893] = 25'b0000001011000101011010010;
    rom[24894] = 25'b0000001011000111011111111;
    rom[24895] = 25'b0000001011001001100101010;
    rom[24896] = 25'b0000001011001011101010110;
    rom[24897] = 25'b0000001011001101110000010;
    rom[24898] = 25'b0000001011001111110101110;
    rom[24899] = 25'b0000001011010001111011010;
    rom[24900] = 25'b0000001011010100000000110;
    rom[24901] = 25'b0000001011010110000110001;
    rom[24902] = 25'b0000001011011000001011110;
    rom[24903] = 25'b0000001011011010010001001;
    rom[24904] = 25'b0000001011011100010110101;
    rom[24905] = 25'b0000001011011110011100000;
    rom[24906] = 25'b0000001011100000100001101;
    rom[24907] = 25'b0000001011100010100111000;
    rom[24908] = 25'b0000001011100100101100100;
    rom[24909] = 25'b0000001011100110110010000;
    rom[24910] = 25'b0000001011101000110111011;
    rom[24911] = 25'b0000001011101010111100111;
    rom[24912] = 25'b0000001011101101000010010;
    rom[24913] = 25'b0000001011101111000111110;
    rom[24914] = 25'b0000001011110001001101010;
    rom[24915] = 25'b0000001011110011010010100;
    rom[24916] = 25'b0000001011110101011000000;
    rom[24917] = 25'b0000001011110111011101100;
    rom[24918] = 25'b0000001011111001100010110;
    rom[24919] = 25'b0000001011111011101000010;
    rom[24920] = 25'b0000001011111101101101110;
    rom[24921] = 25'b0000001011111111110011001;
    rom[24922] = 25'b0000001100000001111000011;
    rom[24923] = 25'b0000001100000011111101111;
    rom[24924] = 25'b0000001100000110000011010;
    rom[24925] = 25'b0000001100001000001000101;
    rom[24926] = 25'b0000001100001010001110000;
    rom[24927] = 25'b0000001100001100010011010;
    rom[24928] = 25'b0000001100001110011000101;
    rom[24929] = 25'b0000001100010000011110000;
    rom[24930] = 25'b0000001100010010100011011;
    rom[24931] = 25'b0000001100010100101000101;
    rom[24932] = 25'b0000001100010110101110000;
    rom[24933] = 25'b0000001100011000110011011;
    rom[24934] = 25'b0000001100011010111000101;
    rom[24935] = 25'b0000001100011100111101111;
    rom[24936] = 25'b0000001100011111000011010;
    rom[24937] = 25'b0000001100100001001000100;
    rom[24938] = 25'b0000001100100011001101110;
    rom[24939] = 25'b0000001100100101010011000;
    rom[24940] = 25'b0000001100100111011000010;
    rom[24941] = 25'b0000001100101001011101100;
    rom[24942] = 25'b0000001100101011100010110;
    rom[24943] = 25'b0000001100101101101000000;
    rom[24944] = 25'b0000001100101111101101001;
    rom[24945] = 25'b0000001100110001110010011;
    rom[24946] = 25'b0000001100110011110111101;
    rom[24947] = 25'b0000001100110101111100110;
    rom[24948] = 25'b0000001100111000000001111;
    rom[24949] = 25'b0000001100111010000111001;
    rom[24950] = 25'b0000001100111100001100001;
    rom[24951] = 25'b0000001100111110010001011;
    rom[24952] = 25'b0000001101000000010110100;
    rom[24953] = 25'b0000001101000010011011101;
    rom[24954] = 25'b0000001101000100100000101;
    rom[24955] = 25'b0000001101000110100101110;
    rom[24956] = 25'b0000001101001000101010111;
    rom[24957] = 25'b0000001101001010101111111;
    rom[24958] = 25'b0000001101001100110101000;
    rom[24959] = 25'b0000001101001110111010000;
    rom[24960] = 25'b0000001101010000111111000;
    rom[24961] = 25'b0000001101010011000100000;
    rom[24962] = 25'b0000001101010101001001000;
    rom[24963] = 25'b0000001101010111001110000;
    rom[24964] = 25'b0000001101011001010011000;
    rom[24965] = 25'b0000001101011011011000000;
    rom[24966] = 25'b0000001101011101011100111;
    rom[24967] = 25'b0000001101011111100001111;
    rom[24968] = 25'b0000001101100001100110110;
    rom[24969] = 25'b0000001101100011101011101;
    rom[24970] = 25'b0000001101100101110000100;
    rom[24971] = 25'b0000001101100111110101011;
    rom[24972] = 25'b0000001101101001111010010;
    rom[24973] = 25'b0000001101101011111111000;
    rom[24974] = 25'b0000001101101110000011111;
    rom[24975] = 25'b0000001101110000001000101;
    rom[24976] = 25'b0000001101110010001101100;
    rom[24977] = 25'b0000001101110100010010010;
    rom[24978] = 25'b0000001101110110010111000;
    rom[24979] = 25'b0000001101111000011011110;
    rom[24980] = 25'b0000001101111010100000100;
    rom[24981] = 25'b0000001101111100100101001;
    rom[24982] = 25'b0000001101111110101001111;
    rom[24983] = 25'b0000001110000000101110100;
    rom[24984] = 25'b0000001110000010110011001;
    rom[24985] = 25'b0000001110000100110111110;
    rom[24986] = 25'b0000001110000110111100100;
    rom[24987] = 25'b0000001110001001000001000;
    rom[24988] = 25'b0000001110001011000101101;
    rom[24989] = 25'b0000001110001101001010010;
    rom[24990] = 25'b0000001110001111001110110;
    rom[24991] = 25'b0000001110010001010011010;
    rom[24992] = 25'b0000001110010011010111110;
    rom[24993] = 25'b0000001110010101011100010;
    rom[24994] = 25'b0000001110010111100000110;
    rom[24995] = 25'b0000001110011001100101001;
    rom[24996] = 25'b0000001110011011101001100;
    rom[24997] = 25'b0000001110011101101110000;
    rom[24998] = 25'b0000001110011111110010011;
    rom[24999] = 25'b0000001110100001110110110;
    rom[25000] = 25'b0000001110100011111011000;
    rom[25001] = 25'b0000001110100101111111011;
    rom[25002] = 25'b0000001110101000000011110;
    rom[25003] = 25'b0000001110101010001000000;
    rom[25004] = 25'b0000001110101100001100010;
    rom[25005] = 25'b0000001110101110010000100;
    rom[25006] = 25'b0000001110110000010100110;
    rom[25007] = 25'b0000001110110010011000111;
    rom[25008] = 25'b0000001110110100011101001;
    rom[25009] = 25'b0000001110110110100001010;
    rom[25010] = 25'b0000001110111000100101011;
    rom[25011] = 25'b0000001110111010101001100;
    rom[25012] = 25'b0000001110111100101101101;
    rom[25013] = 25'b0000001110111110110001101;
    rom[25014] = 25'b0000001111000000110101110;
    rom[25015] = 25'b0000001111000010111001101;
    rom[25016] = 25'b0000001111000100111101110;
    rom[25017] = 25'b0000001111000111000001101;
    rom[25018] = 25'b0000001111001001000101101;
    rom[25019] = 25'b0000001111001011001001100;
    rom[25020] = 25'b0000001111001101001101011;
    rom[25021] = 25'b0000001111001111010001010;
    rom[25022] = 25'b0000001111010001010101001;
    rom[25023] = 25'b0000001111010011011000111;
    rom[25024] = 25'b0000001111010101011100110;
    rom[25025] = 25'b0000001111010111100000100;
    rom[25026] = 25'b0000001111011001100100010;
    rom[25027] = 25'b0000001111011011101000000;
    rom[25028] = 25'b0000001111011101101011101;
    rom[25029] = 25'b0000001111011111101111011;
    rom[25030] = 25'b0000001111100001110011000;
    rom[25031] = 25'b0000001111100011110110101;
    rom[25032] = 25'b0000001111100101111010010;
    rom[25033] = 25'b0000001111100111111101110;
    rom[25034] = 25'b0000001111101010000001010;
    rom[25035] = 25'b0000001111101100000100110;
    rom[25036] = 25'b0000001111101110001000010;
    rom[25037] = 25'b0000001111110000001011110;
    rom[25038] = 25'b0000001111110010001111001;
    rom[25039] = 25'b0000001111110100010010100;
    rom[25040] = 25'b0000001111110110010101111;
    rom[25041] = 25'b0000001111111000011001010;
    rom[25042] = 25'b0000001111111010011100100;
    rom[25043] = 25'b0000001111111100011111111;
    rom[25044] = 25'b0000001111111110100011000;
    rom[25045] = 25'b0000010000000000100110011;
    rom[25046] = 25'b0000010000000010101001100;
    rom[25047] = 25'b0000010000000100101100101;
    rom[25048] = 25'b0000010000000110101111110;
    rom[25049] = 25'b0000010000001000110010111;
    rom[25050] = 25'b0000010000001010110110000;
    rom[25051] = 25'b0000010000001100111001000;
    rom[25052] = 25'b0000010000001110111100000;
    rom[25053] = 25'b0000010000010000111111000;
    rom[25054] = 25'b0000010000010011000010000;
    rom[25055] = 25'b0000010000010101000100111;
    rom[25056] = 25'b0000010000010111000111110;
    rom[25057] = 25'b0000010000011001001010110;
    rom[25058] = 25'b0000010000011011001101100;
    rom[25059] = 25'b0000010000011101010000010;
    rom[25060] = 25'b0000010000011111010011000;
    rom[25061] = 25'b0000010000100001010101110;
    rom[25062] = 25'b0000010000100011011000100;
    rom[25063] = 25'b0000010000100101011011001;
    rom[25064] = 25'b0000010000100111011101110;
    rom[25065] = 25'b0000010000101001100000011;
    rom[25066] = 25'b0000010000101011100010111;
    rom[25067] = 25'b0000010000101101100101100;
    rom[25068] = 25'b0000010000101111101000000;
    rom[25069] = 25'b0000010000110001101010100;
    rom[25070] = 25'b0000010000110011101100111;
    rom[25071] = 25'b0000010000110101101111010;
    rom[25072] = 25'b0000010000110111110001101;
    rom[25073] = 25'b0000010000111001110100000;
    rom[25074] = 25'b0000010000111011110110010;
    rom[25075] = 25'b0000010000111101111000100;
    rom[25076] = 25'b0000010000111111111010110;
    rom[25077] = 25'b0000010001000001111101000;
    rom[25078] = 25'b0000010001000011111111001;
    rom[25079] = 25'b0000010001000110000001010;
    rom[25080] = 25'b0000010001001000000011011;
    rom[25081] = 25'b0000010001001010000101010;
    rom[25082] = 25'b0000010001001100000111011;
    rom[25083] = 25'b0000010001001110001001010;
    rom[25084] = 25'b0000010001010000001011010;
    rom[25085] = 25'b0000010001010010001101010;
    rom[25086] = 25'b0000010001010100001111000;
    rom[25087] = 25'b0000010001010110010000111;
    rom[25088] = 25'b0000010001011000010010101;
    rom[25089] = 25'b0000010001011010010100011;
    rom[25090] = 25'b0000010001011100010110001;
    rom[25091] = 25'b0000010001011110010111110;
    rom[25092] = 25'b0000010001100000011001100;
    rom[25093] = 25'b0000010001100010011011000;
    rom[25094] = 25'b0000010001100100011100101;
    rom[25095] = 25'b0000010001100110011110001;
    rom[25096] = 25'b0000010001101000011111101;
    rom[25097] = 25'b0000010001101010100001000;
    rom[25098] = 25'b0000010001101100100010100;
    rom[25099] = 25'b0000010001101110100011110;
    rom[25100] = 25'b0000010001110000100101001;
    rom[25101] = 25'b0000010001110010100110100;
    rom[25102] = 25'b0000010001110100100111110;
    rom[25103] = 25'b0000010001110110101000111;
    rom[25104] = 25'b0000010001111000101010000;
    rom[25105] = 25'b0000010001111010101011010;
    rom[25106] = 25'b0000010001111100101100010;
    rom[25107] = 25'b0000010001111110101101011;
    rom[25108] = 25'b0000010010000000101110010;
    rom[25109] = 25'b0000010010000010101111010;
    rom[25110] = 25'b0000010010000100110000010;
    rom[25111] = 25'b0000010010000110110001001;
    rom[25112] = 25'b0000010010001000110001111;
    rom[25113] = 25'b0000010010001010110010101;
    rom[25114] = 25'b0000010010001100110011011;
    rom[25115] = 25'b0000010010001110110100001;
    rom[25116] = 25'b0000010010010000110100110;
    rom[25117] = 25'b0000010010010010110101011;
    rom[25118] = 25'b0000010010010100110110000;
    rom[25119] = 25'b0000010010010110110110101;
    rom[25120] = 25'b0000010010011000110111001;
    rom[25121] = 25'b0000010010011010110111100;
    rom[25122] = 25'b0000010010011100110111111;
    rom[25123] = 25'b0000010010011110111000010;
    rom[25124] = 25'b0000010010100000111000100;
    rom[25125] = 25'b0000010010100010111000111;
    rom[25126] = 25'b0000010010100100111001001;
    rom[25127] = 25'b0000010010100110111001010;
    rom[25128] = 25'b0000010010101000111001011;
    rom[25129] = 25'b0000010010101010111001100;
    rom[25130] = 25'b0000010010101100111001100;
    rom[25131] = 25'b0000010010101110111001100;
    rom[25132] = 25'b0000010010110000111001100;
    rom[25133] = 25'b0000010010110010111001011;
    rom[25134] = 25'b0000010010110100111001010;
    rom[25135] = 25'b0000010010110110111001001;
    rom[25136] = 25'b0000010010111000111000111;
    rom[25137] = 25'b0000010010111010111000101;
    rom[25138] = 25'b0000010010111100111000010;
    rom[25139] = 25'b0000010010111110110111111;
    rom[25140] = 25'b0000010011000000110111100;
    rom[25141] = 25'b0000010011000010110111000;
    rom[25142] = 25'b0000010011000100110110011;
    rom[25143] = 25'b0000010011000110110101111;
    rom[25144] = 25'b0000010011001000110101010;
    rom[25145] = 25'b0000010011001010110100101;
    rom[25146] = 25'b0000010011001100110100000;
    rom[25147] = 25'b0000010011001110110011001;
    rom[25148] = 25'b0000010011010000110010011;
    rom[25149] = 25'b0000010011010010110001100;
    rom[25150] = 25'b0000010011010100110000101;
    rom[25151] = 25'b0000010011010110101111101;
    rom[25152] = 25'b0000010011011000101110101;
    rom[25153] = 25'b0000010011011010101101100;
    rom[25154] = 25'b0000010011011100101100100;
    rom[25155] = 25'b0000010011011110101011010;
    rom[25156] = 25'b0000010011100000101010001;
    rom[25157] = 25'b0000010011100010101000111;
    rom[25158] = 25'b0000010011100100100111100;
    rom[25159] = 25'b0000010011100110100110010;
    rom[25160] = 25'b0000010011101000100100111;
    rom[25161] = 25'b0000010011101010100011011;
    rom[25162] = 25'b0000010011101100100001110;
    rom[25163] = 25'b0000010011101110100000010;
    rom[25164] = 25'b0000010011110000011110101;
    rom[25165] = 25'b0000010011110010011101000;
    rom[25166] = 25'b0000010011110100011011010;
    rom[25167] = 25'b0000010011110110011001100;
    rom[25168] = 25'b0000010011111000010111101;
    rom[25169] = 25'b0000010011111010010101110;
    rom[25170] = 25'b0000010011111100010011110;
    rom[25171] = 25'b0000010011111110010001111;
    rom[25172] = 25'b0000010100000000001111110;
    rom[25173] = 25'b0000010100000010001101110;
    rom[25174] = 25'b0000010100000100001011100;
    rom[25175] = 25'b0000010100000110001001010;
    rom[25176] = 25'b0000010100001000000111001;
    rom[25177] = 25'b0000010100001010000100110;
    rom[25178] = 25'b0000010100001100000010011;
    rom[25179] = 25'b0000010100001110000000000;
    rom[25180] = 25'b0000010100001111111101100;
    rom[25181] = 25'b0000010100010001111011000;
    rom[25182] = 25'b0000010100010011111000011;
    rom[25183] = 25'b0000010100010101110101110;
    rom[25184] = 25'b0000010100010111110011000;
    rom[25185] = 25'b0000010100011001110000011;
    rom[25186] = 25'b0000010100011011101101100;
    rom[25187] = 25'b0000010100011101101010101;
    rom[25188] = 25'b0000010100011111100111101;
    rom[25189] = 25'b0000010100100001100100110;
    rom[25190] = 25'b0000010100100011100001101;
    rom[25191] = 25'b0000010100100101011110101;
    rom[25192] = 25'b0000010100100111011011011;
    rom[25193] = 25'b0000010100101001011000010;
    rom[25194] = 25'b0000010100101011010100111;
    rom[25195] = 25'b0000010100101101010001101;
    rom[25196] = 25'b0000010100101111001110010;
    rom[25197] = 25'b0000010100110001001010110;
    rom[25198] = 25'b0000010100110011000111010;
    rom[25199] = 25'b0000010100110101000011110;
    rom[25200] = 25'b0000010100110111000000001;
    rom[25201] = 25'b0000010100111000111100011;
    rom[25202] = 25'b0000010100111010111000110;
    rom[25203] = 25'b0000010100111100110100111;
    rom[25204] = 25'b0000010100111110110001000;
    rom[25205] = 25'b0000010101000000101101001;
    rom[25206] = 25'b0000010101000010101001001;
    rom[25207] = 25'b0000010101000100100101000;
    rom[25208] = 25'b0000010101000110100001000;
    rom[25209] = 25'b0000010101001000011100111;
    rom[25210] = 25'b0000010101001010011000100;
    rom[25211] = 25'b0000010101001100010100010;
    rom[25212] = 25'b0000010101001110001111111;
    rom[25213] = 25'b0000010101010000001011100;
    rom[25214] = 25'b0000010101010010000111000;
    rom[25215] = 25'b0000010101010100000010100;
    rom[25216] = 25'b0000010101010101111110000;
    rom[25217] = 25'b0000010101010111111001010;
    rom[25218] = 25'b0000010101011001110100101;
    rom[25219] = 25'b0000010101011011101111110;
    rom[25220] = 25'b0000010101011101101011000;
    rom[25221] = 25'b0000010101011111100110000;
    rom[25222] = 25'b0000010101100001100001000;
    rom[25223] = 25'b0000010101100011011100000;
    rom[25224] = 25'b0000010101100101010110111;
    rom[25225] = 25'b0000010101100111010001110;
    rom[25226] = 25'b0000010101101001001100100;
    rom[25227] = 25'b0000010101101011000111010;
    rom[25228] = 25'b0000010101101101000001111;
    rom[25229] = 25'b0000010101101110111100100;
    rom[25230] = 25'b0000010101110000110111000;
    rom[25231] = 25'b0000010101110010110001011;
    rom[25232] = 25'b0000010101110100101011110;
    rom[25233] = 25'b0000010101110110100110001;
    rom[25234] = 25'b0000010101111000100000011;
    rom[25235] = 25'b0000010101111010011010101;
    rom[25236] = 25'b0000010101111100010100101;
    rom[25237] = 25'b0000010101111110001110110;
    rom[25238] = 25'b0000010110000000001000110;
    rom[25239] = 25'b0000010110000010000010101;
    rom[25240] = 25'b0000010110000011111100100;
    rom[25241] = 25'b0000010110000101110110010;
    rom[25242] = 25'b0000010110000111110000000;
    rom[25243] = 25'b0000010110001001101001101;
    rom[25244] = 25'b0000010110001011100011010;
    rom[25245] = 25'b0000010110001101011100110;
    rom[25246] = 25'b0000010110001111010110010;
    rom[25247] = 25'b0000010110010001001111100;
    rom[25248] = 25'b0000010110010011001000111;
    rom[25249] = 25'b0000010110010101000010001;
    rom[25250] = 25'b0000010110010110111011010;
    rom[25251] = 25'b0000010110011000110100011;
    rom[25252] = 25'b0000010110011010101101011;
    rom[25253] = 25'b0000010110011100100110011;
    rom[25254] = 25'b0000010110011110011111010;
    rom[25255] = 25'b0000010110100000011000001;
    rom[25256] = 25'b0000010110100010010000111;
    rom[25257] = 25'b0000010110100100001001100;
    rom[25258] = 25'b0000010110100110000010010;
    rom[25259] = 25'b0000010110100111111010110;
    rom[25260] = 25'b0000010110101001110011010;
    rom[25261] = 25'b0000010110101011101011101;
    rom[25262] = 25'b0000010110101101100011111;
    rom[25263] = 25'b0000010110101111011100001;
    rom[25264] = 25'b0000010110110001010100011;
    rom[25265] = 25'b0000010110110011001100100;
    rom[25266] = 25'b0000010110110101000100100;
    rom[25267] = 25'b0000010110110110111100100;
    rom[25268] = 25'b0000010110111000110100011;
    rom[25269] = 25'b0000010110111010101100010;
    rom[25270] = 25'b0000010110111100100100000;
    rom[25271] = 25'b0000010110111110011011101;
    rom[25272] = 25'b0000010111000000010011010;
    rom[25273] = 25'b0000010111000010001010110;
    rom[25274] = 25'b0000010111000100000010010;
    rom[25275] = 25'b0000010111000101111001101;
    rom[25276] = 25'b0000010111000111110001000;
    rom[25277] = 25'b0000010111001001101000001;
    rom[25278] = 25'b0000010111001011011111011;
    rom[25279] = 25'b0000010111001101010110100;
    rom[25280] = 25'b0000010111001111001101100;
    rom[25281] = 25'b0000010111010001000100100;
    rom[25282] = 25'b0000010111010010111011011;
    rom[25283] = 25'b0000010111010100110010001;
    rom[25284] = 25'b0000010111010110101000111;
    rom[25285] = 25'b0000010111011000011111011;
    rom[25286] = 25'b0000010111011010010110000;
    rom[25287] = 25'b0000010111011100001100100;
    rom[25288] = 25'b0000010111011110000011000;
    rom[25289] = 25'b0000010111011111111001010;
    rom[25290] = 25'b0000010111100001101111100;
    rom[25291] = 25'b0000010111100011100101101;
    rom[25292] = 25'b0000010111100101011011110;
    rom[25293] = 25'b0000010111100111010001110;
    rom[25294] = 25'b0000010111101001000111110;
    rom[25295] = 25'b0000010111101010111101101;
    rom[25296] = 25'b0000010111101100110011100;
    rom[25297] = 25'b0000010111101110101001001;
    rom[25298] = 25'b0000010111110000011110110;
    rom[25299] = 25'b0000010111110010010100011;
    rom[25300] = 25'b0000010111110100001001111;
    rom[25301] = 25'b0000010111110101111111010;
    rom[25302] = 25'b0000010111110111110100100;
    rom[25303] = 25'b0000010111111001101001111;
    rom[25304] = 25'b0000010111111011011110111;
    rom[25305] = 25'b0000010111111101010100000;
    rom[25306] = 25'b0000010111111111001001000;
    rom[25307] = 25'b0000011000000000111110000;
    rom[25308] = 25'b0000011000000010110010110;
    rom[25309] = 25'b0000011000000100100111100;
    rom[25310] = 25'b0000011000000110011100010;
    rom[25311] = 25'b0000011000001000010000111;
    rom[25312] = 25'b0000011000001010000101011;
    rom[25313] = 25'b0000011000001011111001111;
    rom[25314] = 25'b0000011000001101101110001;
    rom[25315] = 25'b0000011000001111100010100;
    rom[25316] = 25'b0000011000010001010110101;
    rom[25317] = 25'b0000011000010011001010110;
    rom[25318] = 25'b0000011000010100111110110;
    rom[25319] = 25'b0000011000010110110010110;
    rom[25320] = 25'b0000011000011000100110101;
    rom[25321] = 25'b0000011000011010011010011;
    rom[25322] = 25'b0000011000011100001110001;
    rom[25323] = 25'b0000011000011110000001110;
    rom[25324] = 25'b0000011000011111110101010;
    rom[25325] = 25'b0000011000100001101000110;
    rom[25326] = 25'b0000011000100011011100000;
    rom[25327] = 25'b0000011000100101001111011;
    rom[25328] = 25'b0000011000100111000010100;
    rom[25329] = 25'b0000011000101000110101101;
    rom[25330] = 25'b0000011000101010101000110;
    rom[25331] = 25'b0000011000101100011011110;
    rom[25332] = 25'b0000011000101110001110101;
    rom[25333] = 25'b0000011000110000000001011;
    rom[25334] = 25'b0000011000110001110100000;
    rom[25335] = 25'b0000011000110011100110101;
    rom[25336] = 25'b0000011000110101011001001;
    rom[25337] = 25'b0000011000110111001011101;
    rom[25338] = 25'b0000011000111000111101111;
    rom[25339] = 25'b0000011000111010110000010;
    rom[25340] = 25'b0000011000111100100010011;
    rom[25341] = 25'b0000011000111110010100011;
    rom[25342] = 25'b0000011001000000000110100;
    rom[25343] = 25'b0000011001000001111000011;
    rom[25344] = 25'b0000011001000011101010001;
    rom[25345] = 25'b0000011001000101011011111;
    rom[25346] = 25'b0000011001000111001101100;
    rom[25347] = 25'b0000011001001000111111001;
    rom[25348] = 25'b0000011001001010110000101;
    rom[25349] = 25'b0000011001001100100010000;
    rom[25350] = 25'b0000011001001110010011010;
    rom[25351] = 25'b0000011001010000000100100;
    rom[25352] = 25'b0000011001010001110101101;
    rom[25353] = 25'b0000011001010011100110101;
    rom[25354] = 25'b0000011001010101010111101;
    rom[25355] = 25'b0000011001010111001000100;
    rom[25356] = 25'b0000011001011000111001010;
    rom[25357] = 25'b0000011001011010101001111;
    rom[25358] = 25'b0000011001011100011010100;
    rom[25359] = 25'b0000011001011110001011000;
    rom[25360] = 25'b0000011001011111111011011;
    rom[25361] = 25'b0000011001100001101011110;
    rom[25362] = 25'b0000011001100011011100000;
    rom[25363] = 25'b0000011001100101001100001;
    rom[25364] = 25'b0000011001100110111100001;
    rom[25365] = 25'b0000011001101000101100001;
    rom[25366] = 25'b0000011001101010011100000;
    rom[25367] = 25'b0000011001101100001011110;
    rom[25368] = 25'b0000011001101101111011011;
    rom[25369] = 25'b0000011001101111101011000;
    rom[25370] = 25'b0000011001110001011010100;
    rom[25371] = 25'b0000011001110011001001111;
    rom[25372] = 25'b0000011001110100111001010;
    rom[25373] = 25'b0000011001110110101000011;
    rom[25374] = 25'b0000011001111000010111100;
    rom[25375] = 25'b0000011001111010000110101;
    rom[25376] = 25'b0000011001111011110101100;
    rom[25377] = 25'b0000011001111101100100011;
    rom[25378] = 25'b0000011001111111010011001;
    rom[25379] = 25'b0000011010000001000001110;
    rom[25380] = 25'b0000011010000010110000010;
    rom[25381] = 25'b0000011010000100011110110;
    rom[25382] = 25'b0000011010000110001101001;
    rom[25383] = 25'b0000011010000111111011011;
    rom[25384] = 25'b0000011010001001101001101;
    rom[25385] = 25'b0000011010001011010111110;
    rom[25386] = 25'b0000011010001101000101110;
    rom[25387] = 25'b0000011010001110110011101;
    rom[25388] = 25'b0000011010010000100001011;
    rom[25389] = 25'b0000011010010010001111001;
    rom[25390] = 25'b0000011010010011111100110;
    rom[25391] = 25'b0000011010010101101010010;
    rom[25392] = 25'b0000011010010111010111101;
    rom[25393] = 25'b0000011010011001000101000;
    rom[25394] = 25'b0000011010011010110010001;
    rom[25395] = 25'b0000011010011100011111011;
    rom[25396] = 25'b0000011010011110001100011;
    rom[25397] = 25'b0000011010011111111001011;
    rom[25398] = 25'b0000011010100001100110001;
    rom[25399] = 25'b0000011010100011010010111;
    rom[25400] = 25'b0000011010100100111111100;
    rom[25401] = 25'b0000011010100110101100000;
    rom[25402] = 25'b0000011010101000011000100;
    rom[25403] = 25'b0000011010101010000100111;
    rom[25404] = 25'b0000011010101011110001001;
    rom[25405] = 25'b0000011010101101011101010;
    rom[25406] = 25'b0000011010101111001001010;
    rom[25407] = 25'b0000011010110000110101010;
    rom[25408] = 25'b0000011010110010100001001;
    rom[25409] = 25'b0000011010110100001100110;
    rom[25410] = 25'b0000011010110101111000100;
    rom[25411] = 25'b0000011010110111100100000;
    rom[25412] = 25'b0000011010111001001111100;
    rom[25413] = 25'b0000011010111010111010111;
    rom[25414] = 25'b0000011010111100100110000;
    rom[25415] = 25'b0000011010111110010001010;
    rom[25416] = 25'b0000011010111111111100010;
    rom[25417] = 25'b0000011011000001100111010;
    rom[25418] = 25'b0000011011000011010010000;
    rom[25419] = 25'b0000011011000100111100110;
    rom[25420] = 25'b0000011011000110100111011;
    rom[25421] = 25'b0000011011001000010010000;
    rom[25422] = 25'b0000011011001001111100100;
    rom[25423] = 25'b0000011011001011100110110;
    rom[25424] = 25'b0000011011001101010001000;
    rom[25425] = 25'b0000011011001110111011001;
    rom[25426] = 25'b0000011011010000100101001;
    rom[25427] = 25'b0000011011010010001111001;
    rom[25428] = 25'b0000011011010011111000111;
    rom[25429] = 25'b0000011011010101100010101;
    rom[25430] = 25'b0000011011010111001100010;
    rom[25431] = 25'b0000011011011000110101110;
    rom[25432] = 25'b0000011011011010011111001;
    rom[25433] = 25'b0000011011011100001000011;
    rom[25434] = 25'b0000011011011101110001101;
    rom[25435] = 25'b0000011011011111011010110;
    rom[25436] = 25'b0000011011100001000011110;
    rom[25437] = 25'b0000011011100010101100101;
    rom[25438] = 25'b0000011011100100010101011;
    rom[25439] = 25'b0000011011100101111110000;
    rom[25440] = 25'b0000011011100111100110100;
    rom[25441] = 25'b0000011011101001001111000;
    rom[25442] = 25'b0000011011101010110111011;
    rom[25443] = 25'b0000011011101100011111101;
    rom[25444] = 25'b0000011011101110000111110;
    rom[25445] = 25'b0000011011101111101111111;
    rom[25446] = 25'b0000011011110001010111110;
    rom[25447] = 25'b0000011011110010111111100;
    rom[25448] = 25'b0000011011110100100111010;
    rom[25449] = 25'b0000011011110110001110111;
    rom[25450] = 25'b0000011011110111110110011;
    rom[25451] = 25'b0000011011111001011101110;
    rom[25452] = 25'b0000011011111011000101001;
    rom[25453] = 25'b0000011011111100101100010;
    rom[25454] = 25'b0000011011111110010011010;
    rom[25455] = 25'b0000011011111111111010010;
    rom[25456] = 25'b0000011100000001100001001;
    rom[25457] = 25'b0000011100000011000111111;
    rom[25458] = 25'b0000011100000100101110100;
    rom[25459] = 25'b0000011100000110010101000;
    rom[25460] = 25'b0000011100000111111011100;
    rom[25461] = 25'b0000011100001001100001110;
    rom[25462] = 25'b0000011100001011001000000;
    rom[25463] = 25'b0000011100001100101110000;
    rom[25464] = 25'b0000011100001110010100000;
    rom[25465] = 25'b0000011100001111111001110;
    rom[25466] = 25'b0000011100010001011111101;
    rom[25467] = 25'b0000011100010011000101010;
    rom[25468] = 25'b0000011100010100101010110;
    rom[25469] = 25'b0000011100010110010000010;
    rom[25470] = 25'b0000011100010111110101100;
    rom[25471] = 25'b0000011100011001011010101;
    rom[25472] = 25'b0000011100011010111111111;
    rom[25473] = 25'b0000011100011100100100110;
    rom[25474] = 25'b0000011100011110001001101;
    rom[25475] = 25'b0000011100011111101110011;
    rom[25476] = 25'b0000011100100001010011000;
    rom[25477] = 25'b0000011100100010110111100;
    rom[25478] = 25'b0000011100100100011100000;
    rom[25479] = 25'b0000011100100110000000010;
    rom[25480] = 25'b0000011100100111100100100;
    rom[25481] = 25'b0000011100101001001000100;
    rom[25482] = 25'b0000011100101010101100100;
    rom[25483] = 25'b0000011100101100010000010;
    rom[25484] = 25'b0000011100101101110100000;
    rom[25485] = 25'b0000011100101111010111110;
    rom[25486] = 25'b0000011100110000111011001;
    rom[25487] = 25'b0000011100110010011110101;
    rom[25488] = 25'b0000011100110100000001111;
    rom[25489] = 25'b0000011100110101100101000;
    rom[25490] = 25'b0000011100110111001000000;
    rom[25491] = 25'b0000011100111000101011000;
    rom[25492] = 25'b0000011100111010001101111;
    rom[25493] = 25'b0000011100111011110000100;
    rom[25494] = 25'b0000011100111101010011001;
    rom[25495] = 25'b0000011100111110110101100;
    rom[25496] = 25'b0000011101000000010111111;
    rom[25497] = 25'b0000011101000001111010001;
    rom[25498] = 25'b0000011101000011011100010;
    rom[25499] = 25'b0000011101000100111110010;
    rom[25500] = 25'b0000011101000110100000001;
    rom[25501] = 25'b0000011101001000000001111;
    rom[25502] = 25'b0000011101001001100011100;
    rom[25503] = 25'b0000011101001011000101001;
    rom[25504] = 25'b0000011101001100100110100;
    rom[25505] = 25'b0000011101001110000111111;
    rom[25506] = 25'b0000011101001111101001000;
    rom[25507] = 25'b0000011101010001001010001;
    rom[25508] = 25'b0000011101010010101011000;
    rom[25509] = 25'b0000011101010100001011111;
    rom[25510] = 25'b0000011101010101101100100;
    rom[25511] = 25'b0000011101010111001101001;
    rom[25512] = 25'b0000011101011000101101101;
    rom[25513] = 25'b0000011101011010001101111;
    rom[25514] = 25'b0000011101011011101110010;
    rom[25515] = 25'b0000011101011101001110010;
    rom[25516] = 25'b0000011101011110101110010;
    rom[25517] = 25'b0000011101100000001110001;
    rom[25518] = 25'b0000011101100001101101111;
    rom[25519] = 25'b0000011101100011001101100;
    rom[25520] = 25'b0000011101100100101101000;
    rom[25521] = 25'b0000011101100110001100011;
    rom[25522] = 25'b0000011101100111101011101;
    rom[25523] = 25'b0000011101101001001010111;
    rom[25524] = 25'b0000011101101010101001111;
    rom[25525] = 25'b0000011101101100001000110;
    rom[25526] = 25'b0000011101101101100111101;
    rom[25527] = 25'b0000011101101111000110001;
    rom[25528] = 25'b0000011101110000100100110;
    rom[25529] = 25'b0000011101110010000011010;
    rom[25530] = 25'b0000011101110011100001011;
    rom[25531] = 25'b0000011101110100111111101;
    rom[25532] = 25'b0000011101110110011101110;
    rom[25533] = 25'b0000011101110111111011101;
    rom[25534] = 25'b0000011101111001011001011;
    rom[25535] = 25'b0000011101111010110111001;
    rom[25536] = 25'b0000011101111100010100101;
    rom[25537] = 25'b0000011101111101110010001;
    rom[25538] = 25'b0000011101111111001111011;
    rom[25539] = 25'b0000011110000000101100101;
    rom[25540] = 25'b0000011110000010001001101;
    rom[25541] = 25'b0000011110000011100110100;
    rom[25542] = 25'b0000011110000101000011011;
    rom[25543] = 25'b0000011110000110100000001;
    rom[25544] = 25'b0000011110000111111100101;
    rom[25545] = 25'b0000011110001001011001001;
    rom[25546] = 25'b0000011110001010110101011;
    rom[25547] = 25'b0000011110001100010001100;
    rom[25548] = 25'b0000011110001101101101101;
    rom[25549] = 25'b0000011110001111001001100;
    rom[25550] = 25'b0000011110010000100101011;
    rom[25551] = 25'b0000011110010010000001000;
    rom[25552] = 25'b0000011110010011011100101;
    rom[25553] = 25'b0000011110010100111000001;
    rom[25554] = 25'b0000011110010110010011010;
    rom[25555] = 25'b0000011110010111101110100;
    rom[25556] = 25'b0000011110011001001001101;
    rom[25557] = 25'b0000011110011010100100100;
    rom[25558] = 25'b0000011110011011111111011;
    rom[25559] = 25'b0000011110011101011001111;
    rom[25560] = 25'b0000011110011110110100100;
    rom[25561] = 25'b0000011110100000001110111;
    rom[25562] = 25'b0000011110100001101001010;
    rom[25563] = 25'b0000011110100011000011011;
    rom[25564] = 25'b0000011110100100011101011;
    rom[25565] = 25'b0000011110100101110111010;
    rom[25566] = 25'b0000011110100111010001000;
    rom[25567] = 25'b0000011110101000101010101;
    rom[25568] = 25'b0000011110101010000100001;
    rom[25569] = 25'b0000011110101011011101100;
    rom[25570] = 25'b0000011110101100110110110;
    rom[25571] = 25'b0000011110101110001111111;
    rom[25572] = 25'b0000011110101111101000111;
    rom[25573] = 25'b0000011110110001000001110;
    rom[25574] = 25'b0000011110110010011010100;
    rom[25575] = 25'b0000011110110011110011001;
    rom[25576] = 25'b0000011110110101001011100;
    rom[25577] = 25'b0000011110110110100011111;
    rom[25578] = 25'b0000011110110111111100001;
    rom[25579] = 25'b0000011110111001010100010;
    rom[25580] = 25'b0000011110111010101100001;
    rom[25581] = 25'b0000011110111100000100000;
    rom[25582] = 25'b0000011110111101011011101;
    rom[25583] = 25'b0000011110111110110011001;
    rom[25584] = 25'b0000011111000000001010101;
    rom[25585] = 25'b0000011111000001100001111;
    rom[25586] = 25'b0000011111000010111001000;
    rom[25587] = 25'b0000011111000100010000000;
    rom[25588] = 25'b0000011111000101100110111;
    rom[25589] = 25'b0000011111000110111101101;
    rom[25590] = 25'b0000011111001000010100011;
    rom[25591] = 25'b0000011111001001101010110;
    rom[25592] = 25'b0000011111001011000001001;
    rom[25593] = 25'b0000011111001100010111011;
    rom[25594] = 25'b0000011111001101101101100;
    rom[25595] = 25'b0000011111001111000011011;
    rom[25596] = 25'b0000011111010000011001010;
    rom[25597] = 25'b0000011111010001101110111;
    rom[25598] = 25'b0000011111010011000100011;
    rom[25599] = 25'b0000011111010100011001111;
    rom[25600] = 25'b0000011111010101101111001;
    rom[25601] = 25'b0000011111010111000100010;
    rom[25602] = 25'b0000011111011000011001010;
    rom[25603] = 25'b0000011111011001101110001;
    rom[25604] = 25'b0000011111011011000010111;
    rom[25605] = 25'b0000011111011100010111100;
    rom[25606] = 25'b0000011111011101101100000;
    rom[25607] = 25'b0000011111011111000000011;
    rom[25608] = 25'b0000011111100000010100100;
    rom[25609] = 25'b0000011111100001101000100;
    rom[25610] = 25'b0000011111100010111100100;
    rom[25611] = 25'b0000011111100100010000010;
    rom[25612] = 25'b0000011111100101100011111;
    rom[25613] = 25'b0000011111100110110111011;
    rom[25614] = 25'b0000011111101000001010110;
    rom[25615] = 25'b0000011111101001011110000;
    rom[25616] = 25'b0000011111101010110001001;
    rom[25617] = 25'b0000011111101100000100000;
    rom[25618] = 25'b0000011111101101010110111;
    rom[25619] = 25'b0000011111101110101001100;
    rom[25620] = 25'b0000011111101111111100001;
    rom[25621] = 25'b0000011111110001001110011;
    rom[25622] = 25'b0000011111110010100000110;
    rom[25623] = 25'b0000011111110011110010111;
    rom[25624] = 25'b0000011111110101000100110;
    rom[25625] = 25'b0000011111110110010110110;
    rom[25626] = 25'b0000011111110111101000011;
    rom[25627] = 25'b0000011111111000111001111;
    rom[25628] = 25'b0000011111111010001011011;
    rom[25629] = 25'b0000011111111011011100101;
    rom[25630] = 25'b0000011111111100101101110;
    rom[25631] = 25'b0000011111111101111110111;
    rom[25632] = 25'b0000011111111111001111110;
    rom[25633] = 25'b0000100000000000100000011;
    rom[25634] = 25'b0000100000000001110001000;
    rom[25635] = 25'b0000100000000011000001011;
    rom[25636] = 25'b0000100000000100010001110;
    rom[25637] = 25'b0000100000000101100001111;
    rom[25638] = 25'b0000100000000110110001111;
    rom[25639] = 25'b0000100000001000000001110;
    rom[25640] = 25'b0000100000001001010001100;
    rom[25641] = 25'b0000100000001010100001001;
    rom[25642] = 25'b0000100000001011110000101;
    rom[25643] = 25'b0000100000001100111111111;
    rom[25644] = 25'b0000100000001110001111000;
    rom[25645] = 25'b0000100000001111011110001;
    rom[25646] = 25'b0000100000010000101100111;
    rom[25647] = 25'b0000100000010001111011101;
    rom[25648] = 25'b0000100000010011001010010;
    rom[25649] = 25'b0000100000010100011000110;
    rom[25650] = 25'b0000100000010101100111000;
    rom[25651] = 25'b0000100000010110110101001;
    rom[25652] = 25'b0000100000011000000011001;
    rom[25653] = 25'b0000100000011001010001001;
    rom[25654] = 25'b0000100000011010011110110;
    rom[25655] = 25'b0000100000011011101100011;
    rom[25656] = 25'b0000100000011100111001110;
    rom[25657] = 25'b0000100000011110000111001;
    rom[25658] = 25'b0000100000011111010100010;
    rom[25659] = 25'b0000100000100000100001010;
    rom[25660] = 25'b0000100000100001101110000;
    rom[25661] = 25'b0000100000100010111010111;
    rom[25662] = 25'b0000100000100100000111011;
    rom[25663] = 25'b0000100000100101010011110;
    rom[25664] = 25'b0000100000100110100000001;
    rom[25665] = 25'b0000100000100111101100010;
    rom[25666] = 25'b0000100000101000111000001;
    rom[25667] = 25'b0000100000101010000100000;
    rom[25668] = 25'b0000100000101011001111110;
    rom[25669] = 25'b0000100000101100011011010;
    rom[25670] = 25'b0000100000101101100110101;
    rom[25671] = 25'b0000100000101110110001111;
    rom[25672] = 25'b0000100000101111111101000;
    rom[25673] = 25'b0000100000110001001000000;
    rom[25674] = 25'b0000100000110010010010110;
    rom[25675] = 25'b0000100000110011011101011;
    rom[25676] = 25'b0000100000110100100111111;
    rom[25677] = 25'b0000100000110101110010010;
    rom[25678] = 25'b0000100000110110111100100;
    rom[25679] = 25'b0000100000111000000110100;
    rom[25680] = 25'b0000100000111001010000011;
    rom[25681] = 25'b0000100000111010011010001;
    rom[25682] = 25'b0000100000111011100011110;
    rom[25683] = 25'b0000100000111100101101010;
    rom[25684] = 25'b0000100000111101110110101;
    rom[25685] = 25'b0000100000111110111111110;
    rom[25686] = 25'b0000100001000000001000110;
    rom[25687] = 25'b0000100001000001010001101;
    rom[25688] = 25'b0000100001000010011010010;
    rom[25689] = 25'b0000100001000011100010111;
    rom[25690] = 25'b0000100001000100101011011;
    rom[25691] = 25'b0000100001000101110011101;
    rom[25692] = 25'b0000100001000110111011110;
    rom[25693] = 25'b0000100001001000000011101;
    rom[25694] = 25'b0000100001001001001011011;
    rom[25695] = 25'b0000100001001010010011001;
    rom[25696] = 25'b0000100001001011011010101;
    rom[25697] = 25'b0000100001001100100010000;
    rom[25698] = 25'b0000100001001101101001010;
    rom[25699] = 25'b0000100001001110110000010;
    rom[25700] = 25'b0000100001001111110111001;
    rom[25701] = 25'b0000100001010000111101111;
    rom[25702] = 25'b0000100001010010000100100;
    rom[25703] = 25'b0000100001010011001011000;
    rom[25704] = 25'b0000100001010100010001010;
    rom[25705] = 25'b0000100001010101010111011;
    rom[25706] = 25'b0000100001010110011101011;
    rom[25707] = 25'b0000100001010111100011010;
    rom[25708] = 25'b0000100001011000101000111;
    rom[25709] = 25'b0000100001011001101110011;
    rom[25710] = 25'b0000100001011010110011110;
    rom[25711] = 25'b0000100001011011111000111;
    rom[25712] = 25'b0000100001011100111110000;
    rom[25713] = 25'b0000100001011110000011000;
    rom[25714] = 25'b0000100001011111000111110;
    rom[25715] = 25'b0000100001100000001100011;
    rom[25716] = 25'b0000100001100001010000110;
    rom[25717] = 25'b0000100001100010010101000;
    rom[25718] = 25'b0000100001100011011001001;
    rom[25719] = 25'b0000100001100100011101001;
    rom[25720] = 25'b0000100001100101100000111;
    rom[25721] = 25'b0000100001100110100100101;
    rom[25722] = 25'b0000100001100111101000001;
    rom[25723] = 25'b0000100001101000101011100;
    rom[25724] = 25'b0000100001101001101110110;
    rom[25725] = 25'b0000100001101010110001110;
    rom[25726] = 25'b0000100001101011110100101;
    rom[25727] = 25'b0000100001101100110111010;
    rom[25728] = 25'b0000100001101101111001111;
    rom[25729] = 25'b0000100001101110111100010;
    rom[25730] = 25'b0000100001101111111110101;
    rom[25731] = 25'b0000100001110001000000110;
    rom[25732] = 25'b0000100001110010000010101;
    rom[25733] = 25'b0000100001110011000100011;
    rom[25734] = 25'b0000100001110100000110000;
    rom[25735] = 25'b0000100001110101000111100;
    rom[25736] = 25'b0000100001110110001000111;
    rom[25737] = 25'b0000100001110111001010000;
    rom[25738] = 25'b0000100001111000001011000;
    rom[25739] = 25'b0000100001111001001011111;
    rom[25740] = 25'b0000100001111010001100100;
    rom[25741] = 25'b0000100001111011001101000;
    rom[25742] = 25'b0000100001111100001101011;
    rom[25743] = 25'b0000100001111101001101101;
    rom[25744] = 25'b0000100001111110001101101;
    rom[25745] = 25'b0000100001111111001101100;
    rom[25746] = 25'b0000100010000000001101010;
    rom[25747] = 25'b0000100010000001001100111;
    rom[25748] = 25'b0000100010000010001100010;
    rom[25749] = 25'b0000100010000011001011100;
    rom[25750] = 25'b0000100010000100001010100;
    rom[25751] = 25'b0000100010000101001001100;
    rom[25752] = 25'b0000100010000110001000010;
    rom[25753] = 25'b0000100010000111000110110;
    rom[25754] = 25'b0000100010001000000101010;
    rom[25755] = 25'b0000100010001001000011100;
    rom[25756] = 25'b0000100010001010000001101;
    rom[25757] = 25'b0000100010001010111111101;
    rom[25758] = 25'b0000100010001011111101011;
    rom[25759] = 25'b0000100010001100111011000;
    rom[25760] = 25'b0000100010001101111000100;
    rom[25761] = 25'b0000100010001110110101111;
    rom[25762] = 25'b0000100010001111110011000;
    rom[25763] = 25'b0000100010010000110000000;
    rom[25764] = 25'b0000100010010001101100110;
    rom[25765] = 25'b0000100010010010101001100;
    rom[25766] = 25'b0000100010010011100101111;
    rom[25767] = 25'b0000100010010100100010010;
    rom[25768] = 25'b0000100010010101011110100;
    rom[25769] = 25'b0000100010010110011010011;
    rom[25770] = 25'b0000100010010111010110010;
    rom[25771] = 25'b0000100010011000010010000;
    rom[25772] = 25'b0000100010011001001101100;
    rom[25773] = 25'b0000100010011010001000111;
    rom[25774] = 25'b0000100010011011000100000;
    rom[25775] = 25'b0000100010011011111111000;
    rom[25776] = 25'b0000100010011100111001111;
    rom[25777] = 25'b0000100010011101110100101;
    rom[25778] = 25'b0000100010011110101111001;
    rom[25779] = 25'b0000100010011111101001100;
    rom[25780] = 25'b0000100010100000100011110;
    rom[25781] = 25'b0000100010100001011101110;
    rom[25782] = 25'b0000100010100010010111101;
    rom[25783] = 25'b0000100010100011010001011;
    rom[25784] = 25'b0000100010100100001010111;
    rom[25785] = 25'b0000100010100101000100010;
    rom[25786] = 25'b0000100010100101111101100;
    rom[25787] = 25'b0000100010100110110110100;
    rom[25788] = 25'b0000100010100111101111011;
    rom[25789] = 25'b0000100010101000101000001;
    rom[25790] = 25'b0000100010101001100000101;
    rom[25791] = 25'b0000100010101010011001000;
    rom[25792] = 25'b0000100010101011010001010;
    rom[25793] = 25'b0000100010101100001001010;
    rom[25794] = 25'b0000100010101101000001001;
    rom[25795] = 25'b0000100010101101111000111;
    rom[25796] = 25'b0000100010101110110000011;
    rom[25797] = 25'b0000100010101111100111110;
    rom[25798] = 25'b0000100010110000011111000;
    rom[25799] = 25'b0000100010110001010110000;
    rom[25800] = 25'b0000100010110010001100111;
    rom[25801] = 25'b0000100010110011000011100;
    rom[25802] = 25'b0000100010110011111010000;
    rom[25803] = 25'b0000100010110100110000011;
    rom[25804] = 25'b0000100010110101100110101;
    rom[25805] = 25'b0000100010110110011100101;
    rom[25806] = 25'b0000100010110111010010100;
    rom[25807] = 25'b0000100010111000001000010;
    rom[25808] = 25'b0000100010111000111101110;
    rom[25809] = 25'b0000100010111001110011000;
    rom[25810] = 25'b0000100010111010101000010;
    rom[25811] = 25'b0000100010111011011101010;
    rom[25812] = 25'b0000100010111100010010001;
    rom[25813] = 25'b0000100010111101000110110;
    rom[25814] = 25'b0000100010111101111011010;
    rom[25815] = 25'b0000100010111110101111101;
    rom[25816] = 25'b0000100010111111100011110;
    rom[25817] = 25'b0000100011000000010111110;
    rom[25818] = 25'b0000100011000001001011101;
    rom[25819] = 25'b0000100011000001111111010;
    rom[25820] = 25'b0000100011000010110010101;
    rom[25821] = 25'b0000100011000011100110000;
    rom[25822] = 25'b0000100011000100011001001;
    rom[25823] = 25'b0000100011000101001100000;
    rom[25824] = 25'b0000100011000101111110111;
    rom[25825] = 25'b0000100011000110110001100;
    rom[25826] = 25'b0000100011000111100100000;
    rom[25827] = 25'b0000100011001000010110010;
    rom[25828] = 25'b0000100011001001001000010;
    rom[25829] = 25'b0000100011001001111010010;
    rom[25830] = 25'b0000100011001010101100000;
    rom[25831] = 25'b0000100011001011011101101;
    rom[25832] = 25'b0000100011001100001111000;
    rom[25833] = 25'b0000100011001101000000010;
    rom[25834] = 25'b0000100011001101110001010;
    rom[25835] = 25'b0000100011001110100010001;
    rom[25836] = 25'b0000100011001111010010111;
    rom[25837] = 25'b0000100011010000000011011;
    rom[25838] = 25'b0000100011010000110011110;
    rom[25839] = 25'b0000100011010001100100000;
    rom[25840] = 25'b0000100011010010010100000;
    rom[25841] = 25'b0000100011010011000011111;
    rom[25842] = 25'b0000100011010011110011101;
    rom[25843] = 25'b0000100011010100100011000;
    rom[25844] = 25'b0000100011010101010010011;
    rom[25845] = 25'b0000100011010110000001100;
    rom[25846] = 25'b0000100011010110110000100;
    rom[25847] = 25'b0000100011010111011111010;
    rom[25848] = 25'b0000100011011000001101111;
    rom[25849] = 25'b0000100011011000111100011;
    rom[25850] = 25'b0000100011011001101010101;
    rom[25851] = 25'b0000100011011010011000110;
    rom[25852] = 25'b0000100011011011000110110;
    rom[25853] = 25'b0000100011011011110100011;
    rom[25854] = 25'b0000100011011100100001111;
    rom[25855] = 25'b0000100011011101001111011;
    rom[25856] = 25'b0000100011011101111100101;
    rom[25857] = 25'b0000100011011110101001101;
    rom[25858] = 25'b0000100011011111010110100;
    rom[25859] = 25'b0000100011100000000011001;
    rom[25860] = 25'b0000100011100000101111110;
    rom[25861] = 25'b0000100011100001011100000;
    rom[25862] = 25'b0000100011100010001000001;
    rom[25863] = 25'b0000100011100010110100001;
    rom[25864] = 25'b0000100011100011100000000;
    rom[25865] = 25'b0000100011100100001011100;
    rom[25866] = 25'b0000100011100100110111001;
    rom[25867] = 25'b0000100011100101100010011;
    rom[25868] = 25'b0000100011100110001101011;
    rom[25869] = 25'b0000100011100110111000011;
    rom[25870] = 25'b0000100011100111100011000;
    rom[25871] = 25'b0000100011101000001101101;
    rom[25872] = 25'b0000100011101000111000000;
    rom[25873] = 25'b0000100011101001100010010;
    rom[25874] = 25'b0000100011101010001100010;
    rom[25875] = 25'b0000100011101010110110000;
    rom[25876] = 25'b0000100011101011011111110;
    rom[25877] = 25'b0000100011101100001001001;
    rom[25878] = 25'b0000100011101100110010100;
    rom[25879] = 25'b0000100011101101011011101;
    rom[25880] = 25'b0000100011101110000100100;
    rom[25881] = 25'b0000100011101110101101011;
    rom[25882] = 25'b0000100011101111010101111;
    rom[25883] = 25'b0000100011101111111110011;
    rom[25884] = 25'b0000100011110000100110101;
    rom[25885] = 25'b0000100011110001001110100;
    rom[25886] = 25'b0000100011110001110110011;
    rom[25887] = 25'b0000100011110010011110001;
    rom[25888] = 25'b0000100011110011000101101;
    rom[25889] = 25'b0000100011110011101100111;
    rom[25890] = 25'b0000100011110100010100000;
    rom[25891] = 25'b0000100011110100111011000;
    rom[25892] = 25'b0000100011110101100001111;
    rom[25893] = 25'b0000100011110110001000011;
    rom[25894] = 25'b0000100011110110101110110;
    rom[25895] = 25'b0000100011110111010101001;
    rom[25896] = 25'b0000100011110111111011001;
    rom[25897] = 25'b0000100011111000100001000;
    rom[25898] = 25'b0000100011111001000110101;
    rom[25899] = 25'b0000100011111001101100001;
    rom[25900] = 25'b0000100011111010010001100;
    rom[25901] = 25'b0000100011111010110110101;
    rom[25902] = 25'b0000100011111011011011101;
    rom[25903] = 25'b0000100011111100000000011;
    rom[25904] = 25'b0000100011111100100100111;
    rom[25905] = 25'b0000100011111101001001011;
    rom[25906] = 25'b0000100011111101101101100;
    rom[25907] = 25'b0000100011111110010001101;
    rom[25908] = 25'b0000100011111110110101100;
    rom[25909] = 25'b0000100011111111011001001;
    rom[25910] = 25'b0000100011111111111100101;
    rom[25911] = 25'b0000100100000000011111111;
    rom[25912] = 25'b0000100100000001000011000;
    rom[25913] = 25'b0000100100000001100110000;
    rom[25914] = 25'b0000100100000010001000110;
    rom[25915] = 25'b0000100100000010101011010;
    rom[25916] = 25'b0000100100000011001101110;
    rom[25917] = 25'b0000100100000011101111111;
    rom[25918] = 25'b0000100100000100010001111;
    rom[25919] = 25'b0000100100000100110011110;
    rom[25920] = 25'b0000100100000101010101011;
    rom[25921] = 25'b0000100100000101110110111;
    rom[25922] = 25'b0000100100000110011000001;
    rom[25923] = 25'b0000100100000110111001001;
    rom[25924] = 25'b0000100100000111011010001;
    rom[25925] = 25'b0000100100000111111010110;
    rom[25926] = 25'b0000100100001000011011010;
    rom[25927] = 25'b0000100100001000111011110;
    rom[25928] = 25'b0000100100001001011011111;
    rom[25929] = 25'b0000100100001001111011110;
    rom[25930] = 25'b0000100100001010011011101;
    rom[25931] = 25'b0000100100001010111011001;
    rom[25932] = 25'b0000100100001011011010101;
    rom[25933] = 25'b0000100100001011111001111;
    rom[25934] = 25'b0000100100001100011000111;
    rom[25935] = 25'b0000100100001100110111110;
    rom[25936] = 25'b0000100100001101010110011;
    rom[25937] = 25'b0000100100001101110100111;
    rom[25938] = 25'b0000100100001110010011001;
    rom[25939] = 25'b0000100100001110110001010;
    rom[25940] = 25'b0000100100001111001111001;
    rom[25941] = 25'b0000100100001111101100111;
    rom[25942] = 25'b0000100100010000001010011;
    rom[25943] = 25'b0000100100010000100111110;
    rom[25944] = 25'b0000100100010001000100111;
    rom[25945] = 25'b0000100100010001100001111;
    rom[25946] = 25'b0000100100010001111110110;
    rom[25947] = 25'b0000100100010010011011010;
    rom[25948] = 25'b0000100100010010110111101;
    rom[25949] = 25'b0000100100010011010100000;
    rom[25950] = 25'b0000100100010011110000000;
    rom[25951] = 25'b0000100100010100001011110;
    rom[25952] = 25'b0000100100010100100111100;
    rom[25953] = 25'b0000100100010101000010111;
    rom[25954] = 25'b0000100100010101011110001;
    rom[25955] = 25'b0000100100010101111001010;
    rom[25956] = 25'b0000100100010110010100001;
    rom[25957] = 25'b0000100100010110101110111;
    rom[25958] = 25'b0000100100010111001001011;
    rom[25959] = 25'b0000100100010111100011110;
    rom[25960] = 25'b0000100100010111111101111;
    rom[25961] = 25'b0000100100011000010111110;
    rom[25962] = 25'b0000100100011000110001100;
    rom[25963] = 25'b0000100100011001001011001;
    rom[25964] = 25'b0000100100011001100100011;
    rom[25965] = 25'b0000100100011001111101101;
    rom[25966] = 25'b0000100100011010010110101;
    rom[25967] = 25'b0000100100011010101111011;
    rom[25968] = 25'b0000100100011011001000000;
    rom[25969] = 25'b0000100100011011100000011;
    rom[25970] = 25'b0000100100011011111000110;
    rom[25971] = 25'b0000100100011100010000110;
    rom[25972] = 25'b0000100100011100101000100;
    rom[25973] = 25'b0000100100011101000000001;
    rom[25974] = 25'b0000100100011101010111101;
    rom[25975] = 25'b0000100100011101101110111;
    rom[25976] = 25'b0000100100011110000110000;
    rom[25977] = 25'b0000100100011110011100111;
    rom[25978] = 25'b0000100100011110110011101;
    rom[25979] = 25'b0000100100011111001010001;
    rom[25980] = 25'b0000100100011111100000010;
    rom[25981] = 25'b0000100100011111110110011;
    rom[25982] = 25'b0000100100100000001100011;
    rom[25983] = 25'b0000100100100000100010001;
    rom[25984] = 25'b0000100100100000110111101;
    rom[25985] = 25'b0000100100100001001101000;
    rom[25986] = 25'b0000100100100001100010001;
    rom[25987] = 25'b0000100100100001110111000;
    rom[25988] = 25'b0000100100100010001011111;
    rom[25989] = 25'b0000100100100010100000011;
    rom[25990] = 25'b0000100100100010110100110;
    rom[25991] = 25'b0000100100100011001000111;
    rom[25992] = 25'b0000100100100011011100111;
    rom[25993] = 25'b0000100100100011110000110;
    rom[25994] = 25'b0000100100100100000100011;
    rom[25995] = 25'b0000100100100100010111101;
    rom[25996] = 25'b0000100100100100101010111;
    rom[25997] = 25'b0000100100100100111101111;
    rom[25998] = 25'b0000100100100101010000110;
    rom[25999] = 25'b0000100100100101100011010;
    rom[26000] = 25'b0000100100100101110101110;
    rom[26001] = 25'b0000100100100110001000000;
    rom[26002] = 25'b0000100100100110011010000;
    rom[26003] = 25'b0000100100100110101011111;
    rom[26004] = 25'b0000100100100110111101100;
    rom[26005] = 25'b0000100100100111001111000;
    rom[26006] = 25'b0000100100100111100000001;
    rom[26007] = 25'b0000100100100111110001010;
    rom[26008] = 25'b0000100100101000000010001;
    rom[26009] = 25'b0000100100101000010010110;
    rom[26010] = 25'b0000100100101000100011010;
    rom[26011] = 25'b0000100100101000110011100;
    rom[26012] = 25'b0000100100101001000011101;
    rom[26013] = 25'b0000100100101001010011100;
    rom[26014] = 25'b0000100100101001100011001;
    rom[26015] = 25'b0000100100101001110010101;
    rom[26016] = 25'b0000100100101010000001111;
    rom[26017] = 25'b0000100100101010010001000;
    rom[26018] = 25'b0000100100101010011111111;
    rom[26019] = 25'b0000100100101010101110101;
    rom[26020] = 25'b0000100100101010111101001;
    rom[26021] = 25'b0000100100101011001011011;
    rom[26022] = 25'b0000100100101011011001100;
    rom[26023] = 25'b0000100100101011100111011;
    rom[26024] = 25'b0000100100101011110101001;
    rom[26025] = 25'b0000100100101100000010101;
    rom[26026] = 25'b0000100100101100010000000;
    rom[26027] = 25'b0000100100101100011101001;
    rom[26028] = 25'b0000100100101100101010000;
    rom[26029] = 25'b0000100100101100110110110;
    rom[26030] = 25'b0000100100101101000011010;
    rom[26031] = 25'b0000100100101101001111100;
    rom[26032] = 25'b0000100100101101011011101;
    rom[26033] = 25'b0000100100101101100111101;
    rom[26034] = 25'b0000100100101101110011010;
    rom[26035] = 25'b0000100100101101111110111;
    rom[26036] = 25'b0000100100101110001010010;
    rom[26037] = 25'b0000100100101110010101010;
    rom[26038] = 25'b0000100100101110100000010;
    rom[26039] = 25'b0000100100101110101011000;
    rom[26040] = 25'b0000100100101110110101100;
    rom[26041] = 25'b0000100100101110111111110;
    rom[26042] = 25'b0000100100101111001010000;
    rom[26043] = 25'b0000100100101111010011111;
    rom[26044] = 25'b0000100100101111011101101;
    rom[26045] = 25'b0000100100101111100111001;
    rom[26046] = 25'b0000100100101111110000100;
    rom[26047] = 25'b0000100100101111111001101;
    rom[26048] = 25'b0000100100110000000010101;
    rom[26049] = 25'b0000100100110000001011010;
    rom[26050] = 25'b0000100100110000010011111;
    rom[26051] = 25'b0000100100110000011100001;
    rom[26052] = 25'b0000100100110000100100010;
    rom[26053] = 25'b0000100100110000101100010;
    rom[26054] = 25'b0000100100110000110011111;
    rom[26055] = 25'b0000100100110000111011100;
    rom[26056] = 25'b0000100100110001000010110;
    rom[26057] = 25'b0000100100110001001001111;
    rom[26058] = 25'b0000100100110001010000111;
    rom[26059] = 25'b0000100100110001010111100;
    rom[26060] = 25'b0000100100110001011110001;
    rom[26061] = 25'b0000100100110001100100011;
    rom[26062] = 25'b0000100100110001101010100;
    rom[26063] = 25'b0000100100110001110000011;
    rom[26064] = 25'b0000100100110001110110001;
    rom[26065] = 25'b0000100100110001111011101;
    rom[26066] = 25'b0000100100110010000000111;
    rom[26067] = 25'b0000100100110010000110000;
    rom[26068] = 25'b0000100100110010001010111;
    rom[26069] = 25'b0000100100110010001111101;
    rom[26070] = 25'b0000100100110010010100001;
    rom[26071] = 25'b0000100100110010011000100;
    rom[26072] = 25'b0000100100110010011100100;
    rom[26073] = 25'b0000100100110010100000011;
    rom[26074] = 25'b0000100100110010100100000;
    rom[26075] = 25'b0000100100110010100111101;
    rom[26076] = 25'b0000100100110010101010111;
    rom[26077] = 25'b0000100100110010101101111;
    rom[26078] = 25'b0000100100110010110000111;
    rom[26079] = 25'b0000100100110010110011100;
    rom[26080] = 25'b0000100100110010110101111;
    rom[26081] = 25'b0000100100110010111000010;
    rom[26082] = 25'b0000100100110010111010010;
    rom[26083] = 25'b0000100100110010111100001;
    rom[26084] = 25'b0000100100110010111101110;
    rom[26085] = 25'b0000100100110010111111010;
    rom[26086] = 25'b0000100100110011000000011;
    rom[26087] = 25'b0000100100110011000001100;
    rom[26088] = 25'b0000100100110011000010010;
    rom[26089] = 25'b0000100100110011000011000;
    rom[26090] = 25'b0000100100110011000011011;
    rom[26091] = 25'b0000100100110011000011101;
    rom[26092] = 25'b0000100100110011000011101;
    rom[26093] = 25'b0000100100110011000011011;
    rom[26094] = 25'b0000100100110011000011000;
    rom[26095] = 25'b0000100100110011000010011;
    rom[26096] = 25'b0000100100110011000001100;
    rom[26097] = 25'b0000100100110011000000100;
    rom[26098] = 25'b0000100100110010111111010;
    rom[26099] = 25'b0000100100110010111101111;
    rom[26100] = 25'b0000100100110010111100011;
    rom[26101] = 25'b0000100100110010111010100;
    rom[26102] = 25'b0000100100110010111000011;
    rom[26103] = 25'b0000100100110010110110001;
    rom[26104] = 25'b0000100100110010110011110;
    rom[26105] = 25'b0000100100110010110001000;
    rom[26106] = 25'b0000100100110010101110010;
    rom[26107] = 25'b0000100100110010101011001;
    rom[26108] = 25'b0000100100110010100111111;
    rom[26109] = 25'b0000100100110010100100011;
    rom[26110] = 25'b0000100100110010100000101;
    rom[26111] = 25'b0000100100110010011100110;
    rom[26112] = 25'b0000100100110010011000101;
    rom[26113] = 25'b0000100100110010010100011;
    rom[26114] = 25'b0000100100110010001111111;
    rom[26115] = 25'b0000100100110010001011001;
    rom[26116] = 25'b0000100100110010000110001;
    rom[26117] = 25'b0000100100110010000001000;
    rom[26118] = 25'b0000100100110001111011110;
    rom[26119] = 25'b0000100100110001110110001;
    rom[26120] = 25'b0000100100110001110000011;
    rom[26121] = 25'b0000100100110001101010011;
    rom[26122] = 25'b0000100100110001100100010;
    rom[26123] = 25'b0000100100110001011101111;
    rom[26124] = 25'b0000100100110001010111010;
    rom[26125] = 25'b0000100100110001010000100;
    rom[26126] = 25'b0000100100110001001001100;
    rom[26127] = 25'b0000100100110001000010010;
    rom[26128] = 25'b0000100100110000111010111;
    rom[26129] = 25'b0000100100110000110011010;
    rom[26130] = 25'b0000100100110000101011011;
    rom[26131] = 25'b0000100100110000100011011;
    rom[26132] = 25'b0000100100110000011011000;
    rom[26133] = 25'b0000100100110000010010101;
    rom[26134] = 25'b0000100100110000001010000;
    rom[26135] = 25'b0000100100110000000001001;
    rom[26136] = 25'b0000100100101111110111111;
    rom[26137] = 25'b0000100100101111101110101;
    rom[26138] = 25'b0000100100101111100101001;
    rom[26139] = 25'b0000100100101111011011011;
    rom[26140] = 25'b0000100100101111010001100;
    rom[26141] = 25'b0000100100101111000111011;
    rom[26142] = 25'b0000100100101110111101000;
    rom[26143] = 25'b0000100100101110110010100;
    rom[26144] = 25'b0000100100101110100111110;
    rom[26145] = 25'b0000100100101110011100110;
    rom[26146] = 25'b0000100100101110010001101;
    rom[26147] = 25'b0000100100101110000110001;
    rom[26148] = 25'b0000100100101101111010101;
    rom[26149] = 25'b0000100100101101101110110;
    rom[26150] = 25'b0000100100101101100010110;
    rom[26151] = 25'b0000100100101101010110100;
    rom[26152] = 25'b0000100100101101001010000;
    rom[26153] = 25'b0000100100101100111101011;
    rom[26154] = 25'b0000100100101100110000100;
    rom[26155] = 25'b0000100100101100100011100;
    rom[26156] = 25'b0000100100101100010110010;
    rom[26157] = 25'b0000100100101100001000101;
    rom[26158] = 25'b0000100100101011111010111;
    rom[26159] = 25'b0000100100101011101101000;
    rom[26160] = 25'b0000100100101011011110111;
    rom[26161] = 25'b0000100100101011010000101;
    rom[26162] = 25'b0000100100101011000010000;
    rom[26163] = 25'b0000100100101010110011010;
    rom[26164] = 25'b0000100100101010100100010;
    rom[26165] = 25'b0000100100101010010101001;
    rom[26166] = 25'b0000100100101010000101110;
    rom[26167] = 25'b0000100100101001110110001;
    rom[26168] = 25'b0000100100101001100110011;
    rom[26169] = 25'b0000100100101001010110010;
    rom[26170] = 25'b0000100100101001000110000;
    rom[26171] = 25'b0000100100101000110101101;
    rom[26172] = 25'b0000100100101000100100111;
    rom[26173] = 25'b0000100100101000010100001;
    rom[26174] = 25'b0000100100101000000011000;
    rom[26175] = 25'b0000100100100111110001101;
    rom[26176] = 25'b0000100100100111100000001;
    rom[26177] = 25'b0000100100100111001110011;
    rom[26178] = 25'b0000100100100110111100100;
    rom[26179] = 25'b0000100100100110101010011;
    rom[26180] = 25'b0000100100100110011000000;
    rom[26181] = 25'b0000100100100110000101011;
    rom[26182] = 25'b0000100100100101110010101;
    rom[26183] = 25'b0000100100100101011111101;
    rom[26184] = 25'b0000100100100101001100011;
    rom[26185] = 25'b0000100100100100111001000;
    rom[26186] = 25'b0000100100100100100101011;
    rom[26187] = 25'b0000100100100100010001100;
    rom[26188] = 25'b0000100100100011111101011;
    rom[26189] = 25'b0000100100100011101001001;
    rom[26190] = 25'b0000100100100011010100110;
    rom[26191] = 25'b0000100100100011000000000;
    rom[26192] = 25'b0000100100100010101011000;
    rom[26193] = 25'b0000100100100010010110000;
    rom[26194] = 25'b0000100100100010000000101;
    rom[26195] = 25'b0000100100100001101011001;
    rom[26196] = 25'b0000100100100001010101011;
    rom[26197] = 25'b0000100100100000111111010;
    rom[26198] = 25'b0000100100100000101001001;
    rom[26199] = 25'b0000100100100000010010110;
    rom[26200] = 25'b0000100100011111111100000;
    rom[26201] = 25'b0000100100011111100101010;
    rom[26202] = 25'b0000100100011111001110010;
    rom[26203] = 25'b0000100100011110110110111;
    rom[26204] = 25'b0000100100011110011111011;
    rom[26205] = 25'b0000100100011110000111110;
    rom[26206] = 25'b0000100100011101101111111;
    rom[26207] = 25'b0000100100011101010111101;
    rom[26208] = 25'b0000100100011100111111011;
    rom[26209] = 25'b0000100100011100100110111;
    rom[26210] = 25'b0000100100011100001110001;
    rom[26211] = 25'b0000100100011011110101001;
    rom[26212] = 25'b0000100100011011011011111;
    rom[26213] = 25'b0000100100011011000010100;
    rom[26214] = 25'b0000100100011010101000111;
    rom[26215] = 25'b0000100100011010001111000;
    rom[26216] = 25'b0000100100011001110100111;
    rom[26217] = 25'b0000100100011001011010110;
    rom[26218] = 25'b0000100100011001000000001;
    rom[26219] = 25'b0000100100011000100101100;
    rom[26220] = 25'b0000100100011000001010101;
    rom[26221] = 25'b0000100100010111101111100;
    rom[26222] = 25'b0000100100010111010100001;
    rom[26223] = 25'b0000100100010110111000101;
    rom[26224] = 25'b0000100100010110011100110;
    rom[26225] = 25'b0000100100010110000000111;
    rom[26226] = 25'b0000100100010101100100101;
    rom[26227] = 25'b0000100100010101001000001;
    rom[26228] = 25'b0000100100010100101011100;
    rom[26229] = 25'b0000100100010100001110110;
    rom[26230] = 25'b0000100100010011110001101;
    rom[26231] = 25'b0000100100010011010100011;
    rom[26232] = 25'b0000100100010010110110111;
    rom[26233] = 25'b0000100100010010011001001;
    rom[26234] = 25'b0000100100010001111011001;
    rom[26235] = 25'b0000100100010001011101000;
    rom[26236] = 25'b0000100100010000111110101;
    rom[26237] = 25'b0000100100010000100000000;
    rom[26238] = 25'b0000100100010000000001010;
    rom[26239] = 25'b0000100100001111100010010;
    rom[26240] = 25'b0000100100001111000011000;
    rom[26241] = 25'b0000100100001110100011100;
    rom[26242] = 25'b0000100100001110000011111;
    rom[26243] = 25'b0000100100001101100100000;
    rom[26244] = 25'b0000100100001101000011111;
    rom[26245] = 25'b0000100100001100100011101;
    rom[26246] = 25'b0000100100001100000011001;
    rom[26247] = 25'b0000100100001011100010010;
    rom[26248] = 25'b0000100100001011000001011;
    rom[26249] = 25'b0000100100001010100000001;
    rom[26250] = 25'b0000100100001001111110110;
    rom[26251] = 25'b0000100100001001011101001;
    rom[26252] = 25'b0000100100001000111011011;
    rom[26253] = 25'b0000100100001000011001010;
    rom[26254] = 25'b0000100100000111110111000;
    rom[26255] = 25'b0000100100000111010100100;
    rom[26256] = 25'b0000100100000110110001110;
    rom[26257] = 25'b0000100100000110001110111;
    rom[26258] = 25'b0000100100000101101011110;
    rom[26259] = 25'b0000100100000101001000011;
    rom[26260] = 25'b0000100100000100100100111;
    rom[26261] = 25'b0000100100000100000001000;
    rom[26262] = 25'b0000100100000011011101000;
    rom[26263] = 25'b0000100100000010111000110;
    rom[26264] = 25'b0000100100000010010100011;
    rom[26265] = 25'b0000100100000001101111101;
    rom[26266] = 25'b0000100100000001001010110;
    rom[26267] = 25'b0000100100000000100101110;
    rom[26268] = 25'b0000100100000000000000011;
    rom[26269] = 25'b0000100011111111011010111;
    rom[26270] = 25'b0000100011111110110101001;
    rom[26271] = 25'b0000100011111110001111001;
    rom[26272] = 25'b0000100011111101101000111;
    rom[26273] = 25'b0000100011111101000010100;
    rom[26274] = 25'b0000100011111100011011111;
    rom[26275] = 25'b0000100011111011110101001;
    rom[26276] = 25'b0000100011111011001110000;
    rom[26277] = 25'b0000100011111010100110110;
    rom[26278] = 25'b0000100011111001111111010;
    rom[26279] = 25'b0000100011111001010111100;
    rom[26280] = 25'b0000100011111000101111101;
    rom[26281] = 25'b0000100011111000000111011;
    rom[26282] = 25'b0000100011110111011111000;
    rom[26283] = 25'b0000100011110110110110100;
    rom[26284] = 25'b0000100011110110001101101;
    rom[26285] = 25'b0000100011110101100100100;
    rom[26286] = 25'b0000100011110100111011011;
    rom[26287] = 25'b0000100011110100010001110;
    rom[26288] = 25'b0000100011110011101000001;
    rom[26289] = 25'b0000100011110010111110010;
    rom[26290] = 25'b0000100011110010010100001;
    rom[26291] = 25'b0000100011110001101001110;
    rom[26292] = 25'b0000100011110000111111010;
    rom[26293] = 25'b0000100011110000010100100;
    rom[26294] = 25'b0000100011101111101001011;
    rom[26295] = 25'b0000100011101110111110001;
    rom[26296] = 25'b0000100011101110010010110;
    rom[26297] = 25'b0000100011101101100111001;
    rom[26298] = 25'b0000100011101100111011010;
    rom[26299] = 25'b0000100011101100001111001;
    rom[26300] = 25'b0000100011101011100010110;
    rom[26301] = 25'b0000100011101010110110010;
    rom[26302] = 25'b0000100011101010001001100;
    rom[26303] = 25'b0000100011101001011100100;
    rom[26304] = 25'b0000100011101000101111010;
    rom[26305] = 25'b0000100011101000000001111;
    rom[26306] = 25'b0000100011100111010100010;
    rom[26307] = 25'b0000100011100110100110011;
    rom[26308] = 25'b0000100011100101111000010;
    rom[26309] = 25'b0000100011100101001010000;
    rom[26310] = 25'b0000100011100100011011100;
    rom[26311] = 25'b0000100011100011101100110;
    rom[26312] = 25'b0000100011100010111101110;
    rom[26313] = 25'b0000100011100010001110101;
    rom[26314] = 25'b0000100011100001011111001;
    rom[26315] = 25'b0000100011100000101111100;
    rom[26316] = 25'b0000100011011111111111110;
    rom[26317] = 25'b0000100011011111001111101;
    rom[26318] = 25'b0000100011011110011111011;
    rom[26319] = 25'b0000100011011101101110111;
    rom[26320] = 25'b0000100011011100111110001;
    rom[26321] = 25'b0000100011011100001101010;
    rom[26322] = 25'b0000100011011011011100001;
    rom[26323] = 25'b0000100011011010101010101;
    rom[26324] = 25'b0000100011011001111001001;
    rom[26325] = 25'b0000100011011001000111010;
    rom[26326] = 25'b0000100011011000010101001;
    rom[26327] = 25'b0000100011010111100010111;
    rom[26328] = 25'b0000100011010110110000011;
    rom[26329] = 25'b0000100011010101111101110;
    rom[26330] = 25'b0000100011010101001010110;
    rom[26331] = 25'b0000100011010100010111101;
    rom[26332] = 25'b0000100011010011100100010;
    rom[26333] = 25'b0000100011010010110000110;
    rom[26334] = 25'b0000100011010001111100111;
    rom[26335] = 25'b0000100011010001001000111;
    rom[26336] = 25'b0000100011010000010100101;
    rom[26337] = 25'b0000100011001111100000001;
    rom[26338] = 25'b0000100011001110101011011;
    rom[26339] = 25'b0000100011001101110110100;
    rom[26340] = 25'b0000100011001101000001011;
    rom[26341] = 25'b0000100011001100001100000;
    rom[26342] = 25'b0000100011001011010110011;
    rom[26343] = 25'b0000100011001010100000101;
    rom[26344] = 25'b0000100011001001101010100;
    rom[26345] = 25'b0000100011001000110100010;
    rom[26346] = 25'b0000100011000111111101111;
    rom[26347] = 25'b0000100011000111000111001;
    rom[26348] = 25'b0000100011000110010000010;
    rom[26349] = 25'b0000100011000101011001001;
    rom[26350] = 25'b0000100011000100100001110;
    rom[26351] = 25'b0000100011000011101010001;
    rom[26352] = 25'b0000100011000010110010011;
    rom[26353] = 25'b0000100011000001111010011;
    rom[26354] = 25'b0000100011000001000010001;
    rom[26355] = 25'b0000100011000000001001101;
    rom[26356] = 25'b0000100010111111010001000;
    rom[26357] = 25'b0000100010111110011000001;
    rom[26358] = 25'b0000100010111101011111000;
    rom[26359] = 25'b0000100010111100100101101;
    rom[26360] = 25'b0000100010111011101100000;
    rom[26361] = 25'b0000100010111010110010001;
    rom[26362] = 25'b0000100010111001111000001;
    rom[26363] = 25'b0000100010111000111110000;
    rom[26364] = 25'b0000100010111000000011100;
    rom[26365] = 25'b0000100010110111001000110;
    rom[26366] = 25'b0000100010110110001101111;
    rom[26367] = 25'b0000100010110101010010110;
    rom[26368] = 25'b0000100010110100010111100;
    rom[26369] = 25'b0000100010110011011011111;
    rom[26370] = 25'b0000100010110010100000001;
    rom[26371] = 25'b0000100010110001100100000;
    rom[26372] = 25'b0000100010110000100111111;
    rom[26373] = 25'b0000100010101111101011011;
    rom[26374] = 25'b0000100010101110101110110;
    rom[26375] = 25'b0000100010101101110001111;
    rom[26376] = 25'b0000100010101100110100101;
    rom[26377] = 25'b0000100010101011110111010;
    rom[26378] = 25'b0000100010101010111001110;
    rom[26379] = 25'b0000100010101001111011111;
    rom[26380] = 25'b0000100010101000111101111;
    rom[26381] = 25'b0000100010100111111111110;
    rom[26382] = 25'b0000100010100111000001010;
    rom[26383] = 25'b0000100010100110000010101;
    rom[26384] = 25'b0000100010100101000011101;
    rom[26385] = 25'b0000100010100100000100100;
    rom[26386] = 25'b0000100010100011000101010;
    rom[26387] = 25'b0000100010100010000101101;
    rom[26388] = 25'b0000100010100001000101111;
    rom[26389] = 25'b0000100010100000000101110;
    rom[26390] = 25'b0000100010011111000101100;
    rom[26391] = 25'b0000100010011110000101001;
    rom[26392] = 25'b0000100010011101000100100;
    rom[26393] = 25'b0000100010011100000011100;
    rom[26394] = 25'b0000100010011011000010011;
    rom[26395] = 25'b0000100010011010000001000;
    rom[26396] = 25'b0000100010011000111111011;
    rom[26397] = 25'b0000100010010111111101101;
    rom[26398] = 25'b0000100010010110111011101;
    rom[26399] = 25'b0000100010010101111001011;
    rom[26400] = 25'b0000100010010100110110111;
    rom[26401] = 25'b0000100010010011110100001;
    rom[26402] = 25'b0000100010010010110001011;
    rom[26403] = 25'b0000100010010001101110001;
    rom[26404] = 25'b0000100010010000101010111;
    rom[26405] = 25'b0000100010001111100111010;
    rom[26406] = 25'b0000100010001110100011011;
    rom[26407] = 25'b0000100010001101011111011;
    rom[26408] = 25'b0000100010001100011011001;
    rom[26409] = 25'b0000100010001011010110101;
    rom[26410] = 25'b0000100010001010010010000;
    rom[26411] = 25'b0000100010001001001101001;
    rom[26412] = 25'b0000100010001000001000000;
    rom[26413] = 25'b0000100010000111000010101;
    rom[26414] = 25'b0000100010000101111101000;
    rom[26415] = 25'b0000100010000100110111001;
    rom[26416] = 25'b0000100010000011110001001;
    rom[26417] = 25'b0000100010000010101010111;
    rom[26418] = 25'b0000100010000001100100011;
    rom[26419] = 25'b0000100010000000011101101;
    rom[26420] = 25'b0000100001111111010110110;
    rom[26421] = 25'b0000100001111110001111101;
    rom[26422] = 25'b0000100001111101001000010;
    rom[26423] = 25'b0000100001111100000000101;
    rom[26424] = 25'b0000100001111010111000111;
    rom[26425] = 25'b0000100001111001110000110;
    rom[26426] = 25'b0000100001111000101000101;
    rom[26427] = 25'b0000100001110111100000000;
    rom[26428] = 25'b0000100001110110010111011;
    rom[26429] = 25'b0000100001110101001110011;
    rom[26430] = 25'b0000100001110100000101010;
    rom[26431] = 25'b0000100001110010111011111;
    rom[26432] = 25'b0000100001110001110010010;
    rom[26433] = 25'b0000100001110000101000011;
    rom[26434] = 25'b0000100001101111011110011;
    rom[26435] = 25'b0000100001101110010100001;
    rom[26436] = 25'b0000100001101101001001101;
    rom[26437] = 25'b0000100001101011111110111;
    rom[26438] = 25'b0000100001101010110011111;
    rom[26439] = 25'b0000100001101001101000110;
    rom[26440] = 25'b0000100001101000011101011;
    rom[26441] = 25'b0000100001100111010001111;
    rom[26442] = 25'b0000100001100110000101111;
    rom[26443] = 25'b0000100001100100111001111;
    rom[26444] = 25'b0000100001100011101101101;
    rom[26445] = 25'b0000100001100010100001001;
    rom[26446] = 25'b0000100001100001010100011;
    rom[26447] = 25'b0000100001100000000111011;
    rom[26448] = 25'b0000100001011110111010010;
    rom[26449] = 25'b0000100001011101101100111;
    rom[26450] = 25'b0000100001011100011111010;
    rom[26451] = 25'b0000100001011011010001011;
    rom[26452] = 25'b0000100001011010000011010;
    rom[26453] = 25'b0000100001011000110101000;
    rom[26454] = 25'b0000100001010111100110100;
    rom[26455] = 25'b0000100001010110010111110;
    rom[26456] = 25'b0000100001010101001000111;
    rom[26457] = 25'b0000100001010011111001101;
    rom[26458] = 25'b0000100001010010101010001;
    rom[26459] = 25'b0000100001010001011010101;
    rom[26460] = 25'b0000100001010000001010110;
    rom[26461] = 25'b0000100001001110111010101;
    rom[26462] = 25'b0000100001001101101010011;
    rom[26463] = 25'b0000100001001100011001111;
    rom[26464] = 25'b0000100001001011001001000;
    rom[26465] = 25'b0000100001001001111000001;
    rom[26466] = 25'b0000100001001000100110111;
    rom[26467] = 25'b0000100001000111010101100;
    rom[26468] = 25'b0000100001000110000011111;
    rom[26469] = 25'b0000100001000100110010000;
    rom[26470] = 25'b0000100001000011011111111;
    rom[26471] = 25'b0000100001000010001101101;
    rom[26472] = 25'b0000100001000000111011000;
    rom[26473] = 25'b0000100000111111101000010;
    rom[26474] = 25'b0000100000111110010101010;
    rom[26475] = 25'b0000100000111101000010001;
    rom[26476] = 25'b0000100000111011101110101;
    rom[26477] = 25'b0000100000111010011011000;
    rom[26478] = 25'b0000100000111001000111001;
    rom[26479] = 25'b0000100000110111110011001;
    rom[26480] = 25'b0000100000110110011110110;
    rom[26481] = 25'b0000100000110101001010001;
    rom[26482] = 25'b0000100000110011110101100;
    rom[26483] = 25'b0000100000110010100000100;
    rom[26484] = 25'b0000100000110001001011010;
    rom[26485] = 25'b0000100000101111110101110;
    rom[26486] = 25'b0000100000101110100000001;
    rom[26487] = 25'b0000100000101101001010010;
    rom[26488] = 25'b0000100000101011110100001;
    rom[26489] = 25'b0000100000101010011101111;
    rom[26490] = 25'b0000100000101001000111010;
    rom[26491] = 25'b0000100000100111110000100;
    rom[26492] = 25'b0000100000100110011001100;
    rom[26493] = 25'b0000100000100101000010010;
    rom[26494] = 25'b0000100000100011101010111;
    rom[26495] = 25'b0000100000100010010011001;
    rom[26496] = 25'b0000100000100000111011010;
    rom[26497] = 25'b0000100000011111100011001;
    rom[26498] = 25'b0000100000011110001010111;
    rom[26499] = 25'b0000100000011100110010010;
    rom[26500] = 25'b0000100000011011011001100;
    rom[26501] = 25'b0000100000011010000000011;
    rom[26502] = 25'b0000100000011000100111010;
    rom[26503] = 25'b0000100000010111001101110;
    rom[26504] = 25'b0000100000010101110100001;
    rom[26505] = 25'b0000100000010100011010001;
    rom[26506] = 25'b0000100000010011000000001;
    rom[26507] = 25'b0000100000010001100101110;
    rom[26508] = 25'b0000100000010000001011001;
    rom[26509] = 25'b0000100000001110110000011;
    rom[26510] = 25'b0000100000001101010101011;
    rom[26511] = 25'b0000100000001011111010001;
    rom[26512] = 25'b0000100000001010011110101;
    rom[26513] = 25'b0000100000001001000011000;
    rom[26514] = 25'b0000100000000111100111001;
    rom[26515] = 25'b0000100000000110001010111;
    rom[26516] = 25'b0000100000000100101110100;
    rom[26517] = 25'b0000100000000011010010000;
    rom[26518] = 25'b0000100000000001110101001;
    rom[26519] = 25'b0000100000000000011000001;
    rom[26520] = 25'b0000011111111110111011000;
    rom[26521] = 25'b0000011111111101011101100;
    rom[26522] = 25'b0000011111111011111111111;
    rom[26523] = 25'b0000011111111010100001111;
    rom[26524] = 25'b0000011111111001000011110;
    rom[26525] = 25'b0000011111110111100101011;
    rom[26526] = 25'b0000011111110110000110111;
    rom[26527] = 25'b0000011111110100101000000;
    rom[26528] = 25'b0000011111110011001001000;
    rom[26529] = 25'b0000011111110001101001110;
    rom[26530] = 25'b0000011111110000001010010;
    rom[26531] = 25'b0000011111101110101010101;
    rom[26532] = 25'b0000011111101101001010101;
    rom[26533] = 25'b0000011111101011101010100;
    rom[26534] = 25'b0000011111101010001010001;
    rom[26535] = 25'b0000011111101000101001101;
    rom[26536] = 25'b0000011111100111001000110;
    rom[26537] = 25'b0000011111100101100111110;
    rom[26538] = 25'b0000011111100100000110100;
    rom[26539] = 25'b0000011111100010100101000;
    rom[26540] = 25'b0000011111100001000011011;
    rom[26541] = 25'b0000011111011111100001100;
    rom[26542] = 25'b0000011111011101111111011;
    rom[26543] = 25'b0000011111011100011101000;
    rom[26544] = 25'b0000011111011010111010011;
    rom[26545] = 25'b0000011111011001010111100;
    rom[26546] = 25'b0000011111010111110100100;
    rom[26547] = 25'b0000011111010110010001010;
    rom[26548] = 25'b0000011111010100101101110;
    rom[26549] = 25'b0000011111010011001010001;
    rom[26550] = 25'b0000011111010001100110001;
    rom[26551] = 25'b0000011111010000000010001;
    rom[26552] = 25'b0000011111001110011101101;
    rom[26553] = 25'b0000011111001100111001001;
    rom[26554] = 25'b0000011111001011010100011;
    rom[26555] = 25'b0000011111001001101111010;
    rom[26556] = 25'b0000011111001000001010000;
    rom[26557] = 25'b0000011111000110100100100;
    rom[26558] = 25'b0000011111000100111110111;
    rom[26559] = 25'b0000011111000011011001000;
    rom[26560] = 25'b0000011111000001110010110;
    rom[26561] = 25'b0000011111000000001100100;
    rom[26562] = 25'b0000011110111110100101111;
    rom[26563] = 25'b0000011110111100111111001;
    rom[26564] = 25'b0000011110111011011000000;
    rom[26565] = 25'b0000011110111001110000110;
    rom[26566] = 25'b0000011110111000001001011;
    rom[26567] = 25'b0000011110110110100001101;
    rom[26568] = 25'b0000011110110100111001110;
    rom[26569] = 25'b0000011110110011010001101;
    rom[26570] = 25'b0000011110110001101001010;
    rom[26571] = 25'b0000011110110000000000110;
    rom[26572] = 25'b0000011110101110010111111;
    rom[26573] = 25'b0000011110101100101110111;
    rom[26574] = 25'b0000011110101011000101101;
    rom[26575] = 25'b0000011110101001011100001;
    rom[26576] = 25'b0000011110100111110010100;
    rom[26577] = 25'b0000011110100110001000100;
    rom[26578] = 25'b0000011110100100011110100;
    rom[26579] = 25'b0000011110100010110100001;
    rom[26580] = 25'b0000011110100001001001100;
    rom[26581] = 25'b0000011110011111011110110;
    rom[26582] = 25'b0000011110011101110011110;
    rom[26583] = 25'b0000011110011100001000100;
    rom[26584] = 25'b0000011110011010011101000;
    rom[26585] = 25'b0000011110011000110001011;
    rom[26586] = 25'b0000011110010111000101100;
    rom[26587] = 25'b0000011110010101011001010;
    rom[26588] = 25'b0000011110010011101101000;
    rom[26589] = 25'b0000011110010010000000100;
    rom[26590] = 25'b0000011110010000010011101;
    rom[26591] = 25'b0000011110001110100110110;
    rom[26592] = 25'b0000011110001100111001011;
    rom[26593] = 25'b0000011110001011001100001;
    rom[26594] = 25'b0000011110001001011110011;
    rom[26595] = 25'b0000011110000111110000100;
    rom[26596] = 25'b0000011110000110000010011;
    rom[26597] = 25'b0000011110000100010100000;
    rom[26598] = 25'b0000011110000010100101100;
    rom[26599] = 25'b0000011110000000110110110;
    rom[26600] = 25'b0000011101111111000111110;
    rom[26601] = 25'b0000011101111101011000100;
    rom[26602] = 25'b0000011101111011101001001;
    rom[26603] = 25'b0000011101111001111001100;
    rom[26604] = 25'b0000011101111000001001101;
    rom[26605] = 25'b0000011101110110011001101;
    rom[26606] = 25'b0000011101110100101001010;
    rom[26607] = 25'b0000011101110010111000110;
    rom[26608] = 25'b0000011101110001001000000;
    rom[26609] = 25'b0000011101101111010111000;
    rom[26610] = 25'b0000011101101101100101110;
    rom[26611] = 25'b0000011101101011110100011;
    rom[26612] = 25'b0000011101101010000010110;
    rom[26613] = 25'b0000011101101000010001000;
    rom[26614] = 25'b0000011101100110011110111;
    rom[26615] = 25'b0000011101100100101100101;
    rom[26616] = 25'b0000011101100010111010001;
    rom[26617] = 25'b0000011101100001000111011;
    rom[26618] = 25'b0000011101011111010100011;
    rom[26619] = 25'b0000011101011101100001010;
    rom[26620] = 25'b0000011101011011101101111;
    rom[26621] = 25'b0000011101011001111010010;
    rom[26622] = 25'b0000011101011000000110011;
    rom[26623] = 25'b0000011101010110010010011;
    rom[26624] = 25'b0000011101010100011110001;
    rom[26625] = 25'b0000011101010010101001101;
    rom[26626] = 25'b0000011101010000110101000;
    rom[26627] = 25'b0000011101001111000000000;
    rom[26628] = 25'b0000011101001101001010111;
    rom[26629] = 25'b0000011101001011010101100;
    rom[26630] = 25'b0000011101001001100000000;
    rom[26631] = 25'b0000011101000111101010001;
    rom[26632] = 25'b0000011101000101110100001;
    rom[26633] = 25'b0000011101000011111110000;
    rom[26634] = 25'b0000011101000010000111011;
    rom[26635] = 25'b0000011101000000010000111;
    rom[26636] = 25'b0000011100111110011001111;
    rom[26637] = 25'b0000011100111100100010110;
    rom[26638] = 25'b0000011100111010101011100;
    rom[26639] = 25'b0000011100111000110011111;
    rom[26640] = 25'b0000011100110110111100001;
    rom[26641] = 25'b0000011100110101000100001;
    rom[26642] = 25'b0000011100110011001100000;
    rom[26643] = 25'b0000011100110001010011100;
    rom[26644] = 25'b0000011100101111011010111;
    rom[26645] = 25'b0000011100101101100010000;
    rom[26646] = 25'b0000011100101011101001000;
    rom[26647] = 25'b0000011100101001101111101;
    rom[26648] = 25'b0000011100100111110110010;
    rom[26649] = 25'b0000011100100101111100011;
    rom[26650] = 25'b0000011100100100000010100;
    rom[26651] = 25'b0000011100100010001000010;
    rom[26652] = 25'b0000011100100000001110000;
    rom[26653] = 25'b0000011100011110010011011;
    rom[26654] = 25'b0000011100011100011000100;
    rom[26655] = 25'b0000011100011010011101100;
    rom[26656] = 25'b0000011100011000100010010;
    rom[26657] = 25'b0000011100010110100110111;
    rom[26658] = 25'b0000011100010100101011001;
    rom[26659] = 25'b0000011100010010101111001;
    rom[26660] = 25'b0000011100010000110011000;
    rom[26661] = 25'b0000011100001110110110110;
    rom[26662] = 25'b0000011100001100111010001;
    rom[26663] = 25'b0000011100001010111101011;
    rom[26664] = 25'b0000011100001001000000011;
    rom[26665] = 25'b0000011100000111000011010;
    rom[26666] = 25'b0000011100000101000101110;
    rom[26667] = 25'b0000011100000011001000001;
    rom[26668] = 25'b0000011100000001001010010;
    rom[26669] = 25'b0000011011111111001100001;
    rom[26670] = 25'b0000011011111101001101111;
    rom[26671] = 25'b0000011011111011001111011;
    rom[26672] = 25'b0000011011111001010000101;
    rom[26673] = 25'b0000011011110111010001110;
    rom[26674] = 25'b0000011011110101010010100;
    rom[26675] = 25'b0000011011110011010011001;
    rom[26676] = 25'b0000011011110001010011101;
    rom[26677] = 25'b0000011011101111010011110;
    rom[26678] = 25'b0000011011101101010011101;
    rom[26679] = 25'b0000011011101011010011100;
    rom[26680] = 25'b0000011011101001010011000;
    rom[26681] = 25'b0000011011100111010010011;
    rom[26682] = 25'b0000011011100101010001100;
    rom[26683] = 25'b0000011011100011010000011;
    rom[26684] = 25'b0000011011100001001111000;
    rom[26685] = 25'b0000011011011111001101100;
    rom[26686] = 25'b0000011011011101001011110;
    rom[26687] = 25'b0000011011011011001001110;
    rom[26688] = 25'b0000011011011001000111101;
    rom[26689] = 25'b0000011011010111000101010;
    rom[26690] = 25'b0000011011010101000010101;
    rom[26691] = 25'b0000011011010010111111110;
    rom[26692] = 25'b0000011011010000111100110;
    rom[26693] = 25'b0000011011001110111001011;
    rom[26694] = 25'b0000011011001100110101111;
    rom[26695] = 25'b0000011011001010110010010;
    rom[26696] = 25'b0000011011001000101110011;
    rom[26697] = 25'b0000011011000110101010010;
    rom[26698] = 25'b0000011011000100100101111;
    rom[26699] = 25'b0000011011000010100001010;
    rom[26700] = 25'b0000011011000000011100101;
    rom[26701] = 25'b0000011010111110010111101;
    rom[26702] = 25'b0000011010111100010010011;
    rom[26703] = 25'b0000011010111010001101000;
    rom[26704] = 25'b0000011010111000000111011;
    rom[26705] = 25'b0000011010110110000001100;
    rom[26706] = 25'b0000011010110011111011011;
    rom[26707] = 25'b0000011010110001110101010;
    rom[26708] = 25'b0000011010101111101110110;
    rom[26709] = 25'b0000011010101101101000000;
    rom[26710] = 25'b0000011010101011100001001;
    rom[26711] = 25'b0000011010101001011010000;
    rom[26712] = 25'b0000011010100111010010101;
    rom[26713] = 25'b0000011010100101001011001;
    rom[26714] = 25'b0000011010100011000011011;
    rom[26715] = 25'b0000011010100000111011011;
    rom[26716] = 25'b0000011010011110110011001;
    rom[26717] = 25'b0000011010011100101010110;
    rom[26718] = 25'b0000011010011010100010001;
    rom[26719] = 25'b0000011010011000011001010;
    rom[26720] = 25'b0000011010010110010000010;
    rom[26721] = 25'b0000011010010100000111000;
    rom[26722] = 25'b0000011010010001111101100;
    rom[26723] = 25'b0000011010001111110011111;
    rom[26724] = 25'b0000011010001101101001111;
    rom[26725] = 25'b0000011010001011011111111;
    rom[26726] = 25'b0000011010001001010101100;
    rom[26727] = 25'b0000011010000111001011000;
    rom[26728] = 25'b0000011010000101000000010;
    rom[26729] = 25'b0000011010000010110101010;
    rom[26730] = 25'b0000011010000000101010001;
    rom[26731] = 25'b0000011001111110011110101;
    rom[26732] = 25'b0000011001111100010011000;
    rom[26733] = 25'b0000011001111010000111010;
    rom[26734] = 25'b0000011001110111111011010;
    rom[26735] = 25'b0000011001110101101111000;
    rom[26736] = 25'b0000011001110011100010100;
    rom[26737] = 25'b0000011001110001010101111;
    rom[26738] = 25'b0000011001101111001001001;
    rom[26739] = 25'b0000011001101100111100000;
    rom[26740] = 25'b0000011001101010101110101;
    rom[26741] = 25'b0000011001101000100001010;
    rom[26742] = 25'b0000011001100110010011011;
    rom[26743] = 25'b0000011001100100000101100;
    rom[26744] = 25'b0000011001100001110111011;
    rom[26745] = 25'b0000011001011111101001000;
    rom[26746] = 25'b0000011001011101011010011;
    rom[26747] = 25'b0000011001011011001011110;
    rom[26748] = 25'b0000011001011000111100101;
    rom[26749] = 25'b0000011001010110101101100;
    rom[26750] = 25'b0000011001010100011110001;
    rom[26751] = 25'b0000011001010010001110100;
    rom[26752] = 25'b0000011001001111111110110;
    rom[26753] = 25'b0000011001001101101110101;
    rom[26754] = 25'b0000011001001011011110011;
    rom[26755] = 25'b0000011001001001001110000;
    rom[26756] = 25'b0000011001000110111101010;
    rom[26757] = 25'b0000011001000100101100011;
    rom[26758] = 25'b0000011001000010011011011;
    rom[26759] = 25'b0000011001000000001010000;
    rom[26760] = 25'b0000011000111101111000100;
    rom[26761] = 25'b0000011000111011100110110;
    rom[26762] = 25'b0000011000111001010100111;
    rom[26763] = 25'b0000011000110111000010110;
    rom[26764] = 25'b0000011000110100110000011;
    rom[26765] = 25'b0000011000110010011101110;
    rom[26766] = 25'b0000011000110000001011000;
    rom[26767] = 25'b0000011000101101111000000;
    rom[26768] = 25'b0000011000101011100100111;
    rom[26769] = 25'b0000011000101001010001011;
    rom[26770] = 25'b0000011000100110111101111;
    rom[26771] = 25'b0000011000100100101010000;
    rom[26772] = 25'b0000011000100010010110000;
    rom[26773] = 25'b0000011000100000000001111;
    rom[26774] = 25'b0000011000011101101101011;
    rom[26775] = 25'b0000011000011011011000110;
    rom[26776] = 25'b0000011000011001000011111;
    rom[26777] = 25'b0000011000010110101110111;
    rom[26778] = 25'b0000011000010100011001100;
    rom[26779] = 25'b0000011000010010000100001;
    rom[26780] = 25'b0000011000001111101110011;
    rom[26781] = 25'b0000011000001101011000100;
    rom[26782] = 25'b0000011000001011000010011;
    rom[26783] = 25'b0000011000001000101100001;
    rom[26784] = 25'b0000011000000110010101100;
    rom[26785] = 25'b0000011000000011111110111;
    rom[26786] = 25'b0000011000000001100111111;
    rom[26787] = 25'b0000010111111111010000110;
    rom[26788] = 25'b0000010111111100111001011;
    rom[26789] = 25'b0000010111111010100001111;
    rom[26790] = 25'b0000010111111000001010001;
    rom[26791] = 25'b0000010111110101110010001;
    rom[26792] = 25'b0000010111110011011010000;
    rom[26793] = 25'b0000010111110001000001100;
    rom[26794] = 25'b0000010111101110101001000;
    rom[26795] = 25'b0000010111101100010000001;
    rom[26796] = 25'b0000010111101001110111010;
    rom[26797] = 25'b0000010111100111011110000;
    rom[26798] = 25'b0000010111100101000100101;
    rom[26799] = 25'b0000010111100010101011000;
    rom[26800] = 25'b0000010111100000010001001;
    rom[26801] = 25'b0000010111011101110111001;
    rom[26802] = 25'b0000010111011011011100111;
    rom[26803] = 25'b0000010111011001000010100;
    rom[26804] = 25'b0000010111010110100111110;
    rom[26805] = 25'b0000010111010100001101000;
    rom[26806] = 25'b0000010111010001110001111;
    rom[26807] = 25'b0000010111001111010110101;
    rom[26808] = 25'b0000010111001100111011001;
    rom[26809] = 25'b0000010111001010011111100;
    rom[26810] = 25'b0000010111001000000011101;
    rom[26811] = 25'b0000010111000101100111100;
    rom[26812] = 25'b0000010111000011001011010;
    rom[26813] = 25'b0000010111000000101110110;
    rom[26814] = 25'b0000010110111110010010000;
    rom[26815] = 25'b0000010110111011110101001;
    rom[26816] = 25'b0000010110111001011000000;
    rom[26817] = 25'b0000010110110110111010101;
    rom[26818] = 25'b0000010110110100011101010;
    rom[26819] = 25'b0000010110110001111111100;
    rom[26820] = 25'b0000010110101111100001101;
    rom[26821] = 25'b0000010110101101000011011;
    rom[26822] = 25'b0000010110101010100101001;
    rom[26823] = 25'b0000010110101000000110101;
    rom[26824] = 25'b0000010110100101100111111;
    rom[26825] = 25'b0000010110100011001000111;
    rom[26826] = 25'b0000010110100000101001110;
    rom[26827] = 25'b0000010110011110001010011;
    rom[26828] = 25'b0000010110011011101010111;
    rom[26829] = 25'b0000010110011001001011001;
    rom[26830] = 25'b0000010110010110101011010;
    rom[26831] = 25'b0000010110010100001011000;
    rom[26832] = 25'b0000010110010001101010101;
    rom[26833] = 25'b0000010110001111001010001;
    rom[26834] = 25'b0000010110001100101001011;
    rom[26835] = 25'b0000010110001010001000011;
    rom[26836] = 25'b0000010110000111100111001;
    rom[26837] = 25'b0000010110000101000101110;
    rom[26838] = 25'b0000010110000010100100010;
    rom[26839] = 25'b0000010110000000000010100;
    rom[26840] = 25'b0000010101111101100000100;
    rom[26841] = 25'b0000010101111010111110011;
    rom[26842] = 25'b0000010101111000011100000;
    rom[26843] = 25'b0000010101110101111001011;
    rom[26844] = 25'b0000010101110011010110101;
    rom[26845] = 25'b0000010101110000110011101;
    rom[26846] = 25'b0000010101101110010000011;
    rom[26847] = 25'b0000010101101011101101000;
    rom[26848] = 25'b0000010101101001001001011;
    rom[26849] = 25'b0000010101100110100101110;
    rom[26850] = 25'b0000010101100100000001110;
    rom[26851] = 25'b0000010101100001011101100;
    rom[26852] = 25'b0000010101011110111001001;
    rom[26853] = 25'b0000010101011100010100100;
    rom[26854] = 25'b0000010101011001101111110;
    rom[26855] = 25'b0000010101010111001010110;
    rom[26856] = 25'b0000010101010100100101101;
    rom[26857] = 25'b0000010101010010000000010;
    rom[26858] = 25'b0000010101001111011010101;
    rom[26859] = 25'b0000010101001100110100111;
    rom[26860] = 25'b0000010101001010001110111;
    rom[26861] = 25'b0000010101000111101000110;
    rom[26862] = 25'b0000010101000101000010010;
    rom[26863] = 25'b0000010101000010011011110;
    rom[26864] = 25'b0000010100111111110101000;
    rom[26865] = 25'b0000010100111101001110000;
    rom[26866] = 25'b0000010100111010100110111;
    rom[26867] = 25'b0000010100110111111111011;
    rom[26868] = 25'b0000010100110101010111111;
    rom[26869] = 25'b0000010100110010110000000;
    rom[26870] = 25'b0000010100110000001000001;
    rom[26871] = 25'b0000010100101101100000000;
    rom[26872] = 25'b0000010100101010110111101;
    rom[26873] = 25'b0000010100101000001111000;
    rom[26874] = 25'b0000010100100101100110010;
    rom[26875] = 25'b0000010100100010111101011;
    rom[26876] = 25'b0000010100100000010100010;
    rom[26877] = 25'b0000010100011101101010110;
    rom[26878] = 25'b0000010100011011000001010;
    rom[26879] = 25'b0000010100011000010111100;
    rom[26880] = 25'b0000010100010101101101101;
    rom[26881] = 25'b0000010100010011000011100;
    rom[26882] = 25'b0000010100010000011001001;
    rom[26883] = 25'b0000010100001101101110101;
    rom[26884] = 25'b0000010100001011000011111;
    rom[26885] = 25'b0000010100001000011001000;
    rom[26886] = 25'b0000010100000101101101111;
    rom[26887] = 25'b0000010100000011000010101;
    rom[26888] = 25'b0000010100000000010111000;
    rom[26889] = 25'b0000010011111101101011011;
    rom[26890] = 25'b0000010011111010111111100;
    rom[26891] = 25'b0000010011111000010011011;
    rom[26892] = 25'b0000010011110101100111000;
    rom[26893] = 25'b0000010011110010111010101;
    rom[26894] = 25'b0000010011110000001101111;
    rom[26895] = 25'b0000010011101101100001000;
    rom[26896] = 25'b0000010011101010110100000;
    rom[26897] = 25'b0000010011101000000110110;
    rom[26898] = 25'b0000010011100101011001010;
    rom[26899] = 25'b0000010011100010101011101;
    rom[26900] = 25'b0000010011011111111101110;
    rom[26901] = 25'b0000010011011101001111110;
    rom[26902] = 25'b0000010011011010100001100;
    rom[26903] = 25'b0000010011010111110011000;
    rom[26904] = 25'b0000010011010101000100011;
    rom[26905] = 25'b0000010011010010010101101;
    rom[26906] = 25'b0000010011001111100110101;
    rom[26907] = 25'b0000010011001100110111011;
    rom[26908] = 25'b0000010011001010001000000;
    rom[26909] = 25'b0000010011000111011000100;
    rom[26910] = 25'b0000010011000100101000110;
    rom[26911] = 25'b0000010011000001111000110;
    rom[26912] = 25'b0000010010111111001000100;
    rom[26913] = 25'b0000010010111100011000010;
    rom[26914] = 25'b0000010010111001100111101;
    rom[26915] = 25'b0000010010110110110111000;
    rom[26916] = 25'b0000010010110100000110000;
    rom[26917] = 25'b0000010010110001010100111;
    rom[26918] = 25'b0000010010101110100011101;
    rom[26919] = 25'b0000010010101011110010000;
    rom[26920] = 25'b0000010010101001000000011;
    rom[26921] = 25'b0000010010100110001110100;
    rom[26922] = 25'b0000010010100011011100011;
    rom[26923] = 25'b0000010010100000101010001;
    rom[26924] = 25'b0000010010011101110111101;
    rom[26925] = 25'b0000010010011011000101000;
    rom[26926] = 25'b0000010010011000010010010;
    rom[26927] = 25'b0000010010010101011111001;
    rom[26928] = 25'b0000010010010010101100000;
    rom[26929] = 25'b0000010010001111111000101;
    rom[26930] = 25'b0000010010001101000100111;
    rom[26931] = 25'b0000010010001010010001001;
    rom[26932] = 25'b0000010010000111011101001;
    rom[26933] = 25'b0000010010000100101001000;
    rom[26934] = 25'b0000010010000001110100101;
    rom[26935] = 25'b0000010001111111000000001;
    rom[26936] = 25'b0000010001111100001011011;
    rom[26937] = 25'b0000010001111001010110011;
    rom[26938] = 25'b0000010001110110100001011;
    rom[26939] = 25'b0000010001110011101100000;
    rom[26940] = 25'b0000010001110000110110100;
    rom[26941] = 25'b0000010001101110000000111;
    rom[26942] = 25'b0000010001101011001011000;
    rom[26943] = 25'b0000010001101000010101000;
    rom[26944] = 25'b0000010001100101011110101;
    rom[26945] = 25'b0000010001100010101000010;
    rom[26946] = 25'b0000010001011111110001101;
    rom[26947] = 25'b0000010001011100111010111;
    rom[26948] = 25'b0000010001011010000011110;
    rom[26949] = 25'b0000010001010111001100101;
    rom[26950] = 25'b0000010001010100010101010;
    rom[26951] = 25'b0000010001010001011101110;
    rom[26952] = 25'b0000010001001110100110000;
    rom[26953] = 25'b0000010001001011101110001;
    rom[26954] = 25'b0000010001001000110101111;
    rom[26955] = 25'b0000010001000101111101101;
    rom[26956] = 25'b0000010001000011000101001;
    rom[26957] = 25'b0000010001000000001100100;
    rom[26958] = 25'b0000010000111101010011110;
    rom[26959] = 25'b0000010000111010011010101;
    rom[26960] = 25'b0000010000110111100001011;
    rom[26961] = 25'b0000010000110100101000000;
    rom[26962] = 25'b0000010000110001101110011;
    rom[26963] = 25'b0000010000101110110100101;
    rom[26964] = 25'b0000010000101011111010101;
    rom[26965] = 25'b0000010000101001000000100;
    rom[26966] = 25'b0000010000100110000110010;
    rom[26967] = 25'b0000010000100011001011101;
    rom[26968] = 25'b0000010000100000010000111;
    rom[26969] = 25'b0000010000011101010110001;
    rom[26970] = 25'b0000010000011010011011000;
    rom[26971] = 25'b0000010000010111011111110;
    rom[26972] = 25'b0000010000010100100100010;
    rom[26973] = 25'b0000010000010001101000101;
    rom[26974] = 25'b0000010000001110101100111;
    rom[26975] = 25'b0000010000001011110000111;
    rom[26976] = 25'b0000010000001000110100101;
    rom[26977] = 25'b0000010000000101111000010;
    rom[26978] = 25'b0000010000000010111011111;
    rom[26979] = 25'b0000001111111111111111001;
    rom[26980] = 25'b0000001111111101000010010;
    rom[26981] = 25'b0000001111111010000101001;
    rom[26982] = 25'b0000001111110111000111111;
    rom[26983] = 25'b0000001111110100001010011;
    rom[26984] = 25'b0000001111110001001100110;
    rom[26985] = 25'b0000001111101110001111000;
    rom[26986] = 25'b0000001111101011010001000;
    rom[26987] = 25'b0000001111101000010010110;
    rom[26988] = 25'b0000001111100101010100100;
    rom[26989] = 25'b0000001111100010010110000;
    rom[26990] = 25'b0000001111011111010111001;
    rom[26991] = 25'b0000001111011100011000010;
    rom[26992] = 25'b0000001111011001011001010;
    rom[26993] = 25'b0000001111010110011010000;
    rom[26994] = 25'b0000001111010011011010100;
    rom[26995] = 25'b0000001111010000011011000;
    rom[26996] = 25'b0000001111001101011011001;
    rom[26997] = 25'b0000001111001010011011001;
    rom[26998] = 25'b0000001111000111011011001;
    rom[26999] = 25'b0000001111000100011010101;
    rom[27000] = 25'b0000001111000001011010010;
    rom[27001] = 25'b0000001110111110011001100;
    rom[27002] = 25'b0000001110111011011000101;
    rom[27003] = 25'b0000001110111000010111101;
    rom[27004] = 25'b0000001110110101010110011;
    rom[27005] = 25'b0000001110110010010101000;
    rom[27006] = 25'b0000001110101111010011011;
    rom[27007] = 25'b0000001110101100010001101;
    rom[27008] = 25'b0000001110101001001111101;
    rom[27009] = 25'b0000001110100110001101101;
    rom[27010] = 25'b0000001110100011001011010;
    rom[27011] = 25'b0000001110100000001000110;
    rom[27012] = 25'b0000001110011101000110001;
    rom[27013] = 25'b0000001110011010000011010;
    rom[27014] = 25'b0000001110010111000000010;
    rom[27015] = 25'b0000001110010011111101001;
    rom[27016] = 25'b0000001110010000111001111;
    rom[27017] = 25'b0000001110001101110110010;
    rom[27018] = 25'b0000001110001010110010100;
    rom[27019] = 25'b0000001110000111101110110;
    rom[27020] = 25'b0000001110000100101010101;
    rom[27021] = 25'b0000001110000001100110011;
    rom[27022] = 25'b0000001101111110100010000;
    rom[27023] = 25'b0000001101111011011101011;
    rom[27024] = 25'b0000001101111000011000101;
    rom[27025] = 25'b0000001101110101010011110;
    rom[27026] = 25'b0000001101110010001110101;
    rom[27027] = 25'b0000001101101111001001011;
    rom[27028] = 25'b0000001101101100000011111;
    rom[27029] = 25'b0000001101101000111110010;
    rom[27030] = 25'b0000001101100101111000100;
    rom[27031] = 25'b0000001101100010110010100;
    rom[27032] = 25'b0000001101011111101100011;
    rom[27033] = 25'b0000001101011100100110000;
    rom[27034] = 25'b0000001101011001011111101;
    rom[27035] = 25'b0000001101010110011000111;
    rom[27036] = 25'b0000001101010011010010000;
    rom[27037] = 25'b0000001101010000001011000;
    rom[27038] = 25'b0000001101001101000011111;
    rom[27039] = 25'b0000001101001001111100100;
    rom[27040] = 25'b0000001101000110110101000;
    rom[27041] = 25'b0000001101000011101101010;
    rom[27042] = 25'b0000001101000000100101011;
    rom[27043] = 25'b0000001100111101011101011;
    rom[27044] = 25'b0000001100111010010101001;
    rom[27045] = 25'b0000001100110111001100110;
    rom[27046] = 25'b0000001100110100000100010;
    rom[27047] = 25'b0000001100110000111011100;
    rom[27048] = 25'b0000001100101101110010100;
    rom[27049] = 25'b0000001100101010101001100;
    rom[27050] = 25'b0000001100100111100000010;
    rom[27051] = 25'b0000001100100100010110111;
    rom[27052] = 25'b0000001100100001001101010;
    rom[27053] = 25'b0000001100011110000011100;
    rom[27054] = 25'b0000001100011010111001100;
    rom[27055] = 25'b0000001100010111101111100;
    rom[27056] = 25'b0000001100010100100101010;
    rom[27057] = 25'b0000001100010001011010110;
    rom[27058] = 25'b0000001100001110010000010;
    rom[27059] = 25'b0000001100001011000101011;
    rom[27060] = 25'b0000001100000111111010100;
    rom[27061] = 25'b0000001100000100101111100;
    rom[27062] = 25'b0000001100000001100100001;
    rom[27063] = 25'b0000001011111110011000110;
    rom[27064] = 25'b0000001011111011001101001;
    rom[27065] = 25'b0000001011111000000001011;
    rom[27066] = 25'b0000001011110100110101100;
    rom[27067] = 25'b0000001011110001101001010;
    rom[27068] = 25'b0000001011101110011101001;
    rom[27069] = 25'b0000001011101011010000100;
    rom[27070] = 25'b0000001011101000000100000;
    rom[27071] = 25'b0000001011100100110111010;
    rom[27072] = 25'b0000001011100001101010010;
    rom[27073] = 25'b0000001011011110011101001;
    rom[27074] = 25'b0000001011011011001111111;
    rom[27075] = 25'b0000001011011000000010100;
    rom[27076] = 25'b0000001011010100110100111;
    rom[27077] = 25'b0000001011010001100111001;
    rom[27078] = 25'b0000001011001110011001001;
    rom[27079] = 25'b0000001011001011001011001;
    rom[27080] = 25'b0000001011000111111100110;
    rom[27081] = 25'b0000001011000100101110011;
    rom[27082] = 25'b0000001011000001011111111;
    rom[27083] = 25'b0000001010111110010001000;
    rom[27084] = 25'b0000001010111011000010001;
    rom[27085] = 25'b0000001010110111110011000;
    rom[27086] = 25'b0000001010110100100011110;
    rom[27087] = 25'b0000001010110001010100011;
    rom[27088] = 25'b0000001010101110000100111;
    rom[27089] = 25'b0000001010101010110101000;
    rom[27090] = 25'b0000001010100111100101001;
    rom[27091] = 25'b0000001010100100010101001;
    rom[27092] = 25'b0000001010100001000100111;
    rom[27093] = 25'b0000001010011101110100100;
    rom[27094] = 25'b0000001010011010100100000;
    rom[27095] = 25'b0000001010010111010011010;
    rom[27096] = 25'b0000001010010100000010011;
    rom[27097] = 25'b0000001010010000110001011;
    rom[27098] = 25'b0000001010001101100000001;
    rom[27099] = 25'b0000001010001010001110110;
    rom[27100] = 25'b0000001010000110111101011;
    rom[27101] = 25'b0000001010000011101011101;
    rom[27102] = 25'b0000001010000000011001110;
    rom[27103] = 25'b0000001001111101000111110;
    rom[27104] = 25'b0000001001111001110101101;
    rom[27105] = 25'b0000001001110110100011010;
    rom[27106] = 25'b0000001001110011010000110;
    rom[27107] = 25'b0000001001101111111110010;
    rom[27108] = 25'b0000001001101100101011011;
    rom[27109] = 25'b0000001001101001011000100;
    rom[27110] = 25'b0000001001100110000101010;
    rom[27111] = 25'b0000001001100010110010001;
    rom[27112] = 25'b0000001001011111011110101;
    rom[27113] = 25'b0000001001011100001011000;
    rom[27114] = 25'b0000001001011000110111010;
    rom[27115] = 25'b0000001001010101100011011;
    rom[27116] = 25'b0000001001010010001111011;
    rom[27117] = 25'b0000001001001110111011001;
    rom[27118] = 25'b0000001001001011100110110;
    rom[27119] = 25'b0000001001001000010010001;
    rom[27120] = 25'b0000001001000100111101100;
    rom[27121] = 25'b0000001001000001101000101;
    rom[27122] = 25'b0000001000111110010011101;
    rom[27123] = 25'b0000001000111010111110100;
    rom[27124] = 25'b0000001000110111101001001;
    rom[27125] = 25'b0000001000110100010011101;
    rom[27126] = 25'b0000001000110000111110001;
    rom[27127] = 25'b0000001000101101101000011;
    rom[27128] = 25'b0000001000101010010010011;
    rom[27129] = 25'b0000001000100110111100010;
    rom[27130] = 25'b0000001000100011100110000;
    rom[27131] = 25'b0000001000100000001111101;
    rom[27132] = 25'b0000001000011100111001001;
    rom[27133] = 25'b0000001000011001100010011;
    rom[27134] = 25'b0000001000010110001011100;
    rom[27135] = 25'b0000001000010010110100100;
    rom[27136] = 25'b0000001000001111011101010;
    rom[27137] = 25'b0000001000001100000110000;
    rom[27138] = 25'b0000001000001000101110100;
    rom[27139] = 25'b0000001000000101010110111;
    rom[27140] = 25'b0000001000000001111111000;
    rom[27141] = 25'b0000000111111110100111001;
    rom[27142] = 25'b0000000111111011001111000;
    rom[27143] = 25'b0000000111110111110110111;
    rom[27144] = 25'b0000000111110100011110100;
    rom[27145] = 25'b0000000111110001000101111;
    rom[27146] = 25'b0000000111101101101101001;
    rom[27147] = 25'b0000000111101010010100010;
    rom[27148] = 25'b0000000111100110111011011;
    rom[27149] = 25'b0000000111100011100010010;
    rom[27150] = 25'b0000000111100000001000111;
    rom[27151] = 25'b0000000111011100101111100;
    rom[27152] = 25'b0000000111011001010101111;
    rom[27153] = 25'b0000000111010101111100001;
    rom[27154] = 25'b0000000111010010100010010;
    rom[27155] = 25'b0000000111001111001000001;
    rom[27156] = 25'b0000000111001011101110000;
    rom[27157] = 25'b0000000111001000010011101;
    rom[27158] = 25'b0000000111000100111001001;
    rom[27159] = 25'b0000000111000001011110100;
    rom[27160] = 25'b0000000110111110000011110;
    rom[27161] = 25'b0000000110111010101000110;
    rom[27162] = 25'b0000000110110111001101101;
    rom[27163] = 25'b0000000110110011110010100;
    rom[27164] = 25'b0000000110110000010111001;
    rom[27165] = 25'b0000000110101100111011100;
    rom[27166] = 25'b0000000110101001011111110;
    rom[27167] = 25'b0000000110100110000100000;
    rom[27168] = 25'b0000000110100010101000000;
    rom[27169] = 25'b0000000110011111001011111;
    rom[27170] = 25'b0000000110011011101111101;
    rom[27171] = 25'b0000000110011000010011010;
    rom[27172] = 25'b0000000110010100110110101;
    rom[27173] = 25'b0000000110010001011010000;
    rom[27174] = 25'b0000000110001101111101001;
    rom[27175] = 25'b0000000110001010100000001;
    rom[27176] = 25'b0000000110000111000011000;
    rom[27177] = 25'b0000000110000011100101101;
    rom[27178] = 25'b0000000110000000001000010;
    rom[27179] = 25'b0000000101111100101010101;
    rom[27180] = 25'b0000000101111001001101000;
    rom[27181] = 25'b0000000101110101101111001;
    rom[27182] = 25'b0000000101110010010001001;
    rom[27183] = 25'b0000000101101110110010111;
    rom[27184] = 25'b0000000101101011010100101;
    rom[27185] = 25'b0000000101100111110110010;
    rom[27186] = 25'b0000000101100100010111101;
    rom[27187] = 25'b0000000101100000111000111;
    rom[27188] = 25'b0000000101011101011010001;
    rom[27189] = 25'b0000000101011001111011001;
    rom[27190] = 25'b0000000101010110011011111;
    rom[27191] = 25'b0000000101010010111100101;
    rom[27192] = 25'b0000000101001111011101010;
    rom[27193] = 25'b0000000101001011111101101;
    rom[27194] = 25'b0000000101001000011101111;
    rom[27195] = 25'b0000000101000100111110001;
    rom[27196] = 25'b0000000101000001011110000;
    rom[27197] = 25'b0000000100111101111101111;
    rom[27198] = 25'b0000000100111010011101101;
    rom[27199] = 25'b0000000100110110111101010;
    rom[27200] = 25'b0000000100110011011100101;
    rom[27201] = 25'b0000000100101111111100000;
    rom[27202] = 25'b0000000100101100011011010;
    rom[27203] = 25'b0000000100101000111010010;
    rom[27204] = 25'b0000000100100101011001001;
    rom[27205] = 25'b0000000100100001110111111;
    rom[27206] = 25'b0000000100011110010110100;
    rom[27207] = 25'b0000000100011010110101000;
    rom[27208] = 25'b0000000100010111010011010;
    rom[27209] = 25'b0000000100010011110001011;
    rom[27210] = 25'b0000000100010000001111100;
    rom[27211] = 25'b0000000100001100101101011;
    rom[27212] = 25'b0000000100001001001011010;
    rom[27213] = 25'b0000000100000101101000111;
    rom[27214] = 25'b0000000100000010000110011;
    rom[27215] = 25'b0000000011111110100011110;
    rom[27216] = 25'b0000000011111011000001000;
    rom[27217] = 25'b0000000011110111011110001;
    rom[27218] = 25'b0000000011110011111011001;
    rom[27219] = 25'b0000000011110000011000000;
    rom[27220] = 25'b0000000011101100110100101;
    rom[27221] = 25'b0000000011101001010001001;
    rom[27222] = 25'b0000000011100101101101101;
    rom[27223] = 25'b0000000011100010001001111;
    rom[27224] = 25'b0000000011011110100110001;
    rom[27225] = 25'b0000000011011011000010001;
    rom[27226] = 25'b0000000011010111011110000;
    rom[27227] = 25'b0000000011010011111001110;
    rom[27228] = 25'b0000000011010000010101011;
    rom[27229] = 25'b0000000011001100110001000;
    rom[27230] = 25'b0000000011001001001100010;
    rom[27231] = 25'b0000000011000101100111100;
    rom[27232] = 25'b0000000011000010000010100;
    rom[27233] = 25'b0000000010111110011101100;
    rom[27234] = 25'b0000000010111010111000011;
    rom[27235] = 25'b0000000010110111010011001;
    rom[27236] = 25'b0000000010110011101101101;
    rom[27237] = 25'b0000000010110000001000001;
    rom[27238] = 25'b0000000010101100100010011;
    rom[27239] = 25'b0000000010101000111100101;
    rom[27240] = 25'b0000000010100101010110101;
    rom[27241] = 25'b0000000010100001110000100;
    rom[27242] = 25'b0000000010011110001010011;
    rom[27243] = 25'b0000000010011010100100000;
    rom[27244] = 25'b0000000010010110111101100;
    rom[27245] = 25'b0000000010010011010110111;
    rom[27246] = 25'b0000000010001111110000001;
    rom[27247] = 25'b0000000010001100001001010;
    rom[27248] = 25'b0000000010001000100010011;
    rom[27249] = 25'b0000000010000100111011010;
    rom[27250] = 25'b0000000010000001010100000;
    rom[27251] = 25'b0000000001111101101100101;
    rom[27252] = 25'b0000000001111010000101001;
    rom[27253] = 25'b0000000001110110011101100;
    rom[27254] = 25'b0000000001110010110101110;
    rom[27255] = 25'b0000000001101111001101111;
    rom[27256] = 25'b0000000001101011100101111;
    rom[27257] = 25'b0000000001100111111101101;
    rom[27258] = 25'b0000000001100100010101011;
    rom[27259] = 25'b0000000001100000101101001;
    rom[27260] = 25'b0000000001011101000100100;
    rom[27261] = 25'b0000000001011001011011111;
    rom[27262] = 25'b0000000001010101110011010;
    rom[27263] = 25'b0000000001010010001010010;
    rom[27264] = 25'b0000000001001110100001010;
    rom[27265] = 25'b0000000001001010111000001;
    rom[27266] = 25'b0000000001000111001110111;
    rom[27267] = 25'b0000000001000011100101011;
    rom[27268] = 25'b0000000000111111111100000;
    rom[27269] = 25'b0000000000111100010010011;
    rom[27270] = 25'b0000000000111000101000101;
    rom[27271] = 25'b0000000000110100111110110;
    rom[27272] = 25'b0000000000110001010100110;
    rom[27273] = 25'b0000000000101101101010101;
    rom[27274] = 25'b0000000000101010000000011;
    rom[27275] = 25'b0000000000100110010110000;
    rom[27276] = 25'b0000000000100010101011100;
    rom[27277] = 25'b0000000000011111000000111;
    rom[27278] = 25'b0000000000011011010110010;
    rom[27279] = 25'b0000000000010111101011011;
    rom[27280] = 25'b0000000000010100000000011;
    rom[27281] = 25'b0000000000010000010101010;
    rom[27282] = 25'b0000000000001100101010001;
    rom[27283] = 25'b0000000000001000111110110;
    rom[27284] = 25'b0000000000000101010011010;
    rom[27285] = 25'b0000000000000001100111110;
    rom[27286] = 25'b1111111111111101111100001;
    rom[27287] = 25'b1111111111111010010000010;
    rom[27288] = 25'b1111111111110110100100011;
    rom[27289] = 25'b1111111111110010111000010;
    rom[27290] = 25'b1111111111101111001100001;
    rom[27291] = 25'b1111111111101011011111111;
    rom[27292] = 25'b1111111111100111110011011;
    rom[27293] = 25'b1111111111100100000111000;
    rom[27294] = 25'b1111111111100000011010010;
    rom[27295] = 25'b1111111111011100101101100;
    rom[27296] = 25'b1111111111011001000000101;
    rom[27297] = 25'b1111111111010101010011110;
    rom[27298] = 25'b1111111111010001100110101;
    rom[27299] = 25'b1111111111001101111001010;
    rom[27300] = 25'b1111111111001010001100000;
    rom[27301] = 25'b1111111111000110011110100;
    rom[27302] = 25'b1111111111000010110001000;
    rom[27303] = 25'b1111111110111111000011010;
    rom[27304] = 25'b1111111110111011010101100;
    rom[27305] = 25'b1111111110110111100111101;
    rom[27306] = 25'b1111111110110011111001101;
    rom[27307] = 25'b1111111110110000001011100;
    rom[27308] = 25'b1111111110101100011101010;
    rom[27309] = 25'b1111111110101000101110111;
    rom[27310] = 25'b1111111110100101000000011;
    rom[27311] = 25'b1111111110100001010001111;
    rom[27312] = 25'b1111111110011101100011001;
    rom[27313] = 25'b1111111110011001110100010;
    rom[27314] = 25'b1111111110010110000101011;
    rom[27315] = 25'b1111111110010010010110010;
    rom[27316] = 25'b1111111110001110100111001;
    rom[27317] = 25'b1111111110001010110111111;
    rom[27318] = 25'b1111111110000111001000100;
    rom[27319] = 25'b1111111110000011011001000;
    rom[27320] = 25'b1111111101111111101001011;
    rom[27321] = 25'b1111111101111011111001110;
    rom[27322] = 25'b1111111101111000001001111;
    rom[27323] = 25'b1111111101110100011010000;
    rom[27324] = 25'b1111111101110000101010000;
    rom[27325] = 25'b1111111101101100111001110;
    rom[27326] = 25'b1111111101101001001001101;
    rom[27327] = 25'b1111111101100101011001010;
    rom[27328] = 25'b1111111101100001101000110;
    rom[27329] = 25'b1111111101011101111000001;
    rom[27330] = 25'b1111111101011010000111011;
    rom[27331] = 25'b1111111101010110010110101;
    rom[27332] = 25'b1111111101010010100101110;
    rom[27333] = 25'b1111111101001110110100110;
    rom[27334] = 25'b1111111101001011000011101;
    rom[27335] = 25'b1111111101000111010010100;
    rom[27336] = 25'b1111111101000011100001001;
    rom[27337] = 25'b1111111100111111101111101;
    rom[27338] = 25'b1111111100111011111110001;
    rom[27339] = 25'b1111111100111000001100100;
    rom[27340] = 25'b1111111100110100011010110;
    rom[27341] = 25'b1111111100110000101000111;
    rom[27342] = 25'b1111111100101100110110111;
    rom[27343] = 25'b1111111100101001000100111;
    rom[27344] = 25'b1111111100100101010010110;
    rom[27345] = 25'b1111111100100001100000011;
    rom[27346] = 25'b1111111100011101101110000;
    rom[27347] = 25'b1111111100011001111011100;
    rom[27348] = 25'b1111111100010110001001000;
    rom[27349] = 25'b1111111100010010010110010;
    rom[27350] = 25'b1111111100001110100011100;
    rom[27351] = 25'b1111111100001010110000101;
    rom[27352] = 25'b1111111100000110111101101;
    rom[27353] = 25'b1111111100000011001010100;
    rom[27354] = 25'b1111111011111111010111010;
    rom[27355] = 25'b1111111011111011100100000;
    rom[27356] = 25'b1111111011110111110000101;
    rom[27357] = 25'b1111111011110011111101001;
    rom[27358] = 25'b1111111011110000001001100;
    rom[27359] = 25'b1111111011101100010101111;
    rom[27360] = 25'b1111111011101000100010000;
    rom[27361] = 25'b1111111011100100101110000;
    rom[27362] = 25'b1111111011100000111010001;
    rom[27363] = 25'b1111111011011101000110000;
    rom[27364] = 25'b1111111011011001010001111;
    rom[27365] = 25'b1111111011010101011101100;
    rom[27366] = 25'b1111111011010001101001001;
    rom[27367] = 25'b1111111011001101110100101;
    rom[27368] = 25'b1111111011001010000000000;
    rom[27369] = 25'b1111111011000110001011010;
    rom[27370] = 25'b1111111011000010010110100;
    rom[27371] = 25'b1111111010111110100001101;
    rom[27372] = 25'b1111111010111010101100110;
    rom[27373] = 25'b1111111010110110110111100;
    rom[27374] = 25'b1111111010110011000010011;
    rom[27375] = 25'b1111111010101111001101001;
    rom[27376] = 25'b1111111010101011010111110;
    rom[27377] = 25'b1111111010100111100010011;
    rom[27378] = 25'b1111111010100011101100110;
    rom[27379] = 25'b1111111010011111110111001;
    rom[27380] = 25'b1111111010011100000001011;
    rom[27381] = 25'b1111111010011000001011100;
    rom[27382] = 25'b1111111010010100010101100;
    rom[27383] = 25'b1111111010010000011111101;
    rom[27384] = 25'b1111111010001100101001011;
    rom[27385] = 25'b1111111010001000110011010;
    rom[27386] = 25'b1111111010000100111100111;
    rom[27387] = 25'b1111111010000001000110100;
    rom[27388] = 25'b1111111001111101010000001;
    rom[27389] = 25'b1111111001111001011001100;
    rom[27390] = 25'b1111111001110101100010110;
    rom[27391] = 25'b1111111001110001101100000;
    rom[27392] = 25'b1111111001101101110101001;
    rom[27393] = 25'b1111111001101001111110001;
    rom[27394] = 25'b1111111001100110000111001;
    rom[27395] = 25'b1111111001100010010000000;
    rom[27396] = 25'b1111111001011110011000111;
    rom[27397] = 25'b1111111001011010100001100;
    rom[27398] = 25'b1111111001010110101010001;
    rom[27399] = 25'b1111111001010010110010101;
    rom[27400] = 25'b1111111001001110111011000;
    rom[27401] = 25'b1111111001001011000011011;
    rom[27402] = 25'b1111111001000111001011101;
    rom[27403] = 25'b1111111001000011010011110;
    rom[27404] = 25'b1111111000111111011011111;
    rom[27405] = 25'b1111111000111011100011110;
    rom[27406] = 25'b1111111000110111101011101;
    rom[27407] = 25'b1111111000110011110011100;
    rom[27408] = 25'b1111111000101111111011010;
    rom[27409] = 25'b1111111000101100000010111;
    rom[27410] = 25'b1111111000101000001010011;
    rom[27411] = 25'b1111111000100100010001111;
    rom[27412] = 25'b1111111000100000011001010;
    rom[27413] = 25'b1111111000011100100000100;
    rom[27414] = 25'b1111111000011000100111110;
    rom[27415] = 25'b1111111000010100101110111;
    rom[27416] = 25'b1111111000010000110101111;
    rom[27417] = 25'b1111111000001100111100111;
    rom[27418] = 25'b1111111000001001000011101;
    rom[27419] = 25'b1111111000000101001010100;
    rom[27420] = 25'b1111111000000001010001001;
    rom[27421] = 25'b1111110111111101010111111;
    rom[27422] = 25'b1111110111111001011110011;
    rom[27423] = 25'b1111110111110101100100110;
    rom[27424] = 25'b1111110111110001101011001;
    rom[27425] = 25'b1111110111101101110001011;
    rom[27426] = 25'b1111110111101001110111101;
    rom[27427] = 25'b1111110111100101111101110;
    rom[27428] = 25'b1111110111100010000011110;
    rom[27429] = 25'b1111110111011110001001111;
    rom[27430] = 25'b1111110111011010001111110;
    rom[27431] = 25'b1111110111010110010101100;
    rom[27432] = 25'b1111110111010010011011001;
    rom[27433] = 25'b1111110111001110100000110;
    rom[27434] = 25'b1111110111001010100110011;
    rom[27435] = 25'b1111110111000110101011111;
    rom[27436] = 25'b1111110111000010110001011;
    rom[27437] = 25'b1111110110111110110110101;
    rom[27438] = 25'b1111110110111010111011111;
    rom[27439] = 25'b1111110110110111000001001;
    rom[27440] = 25'b1111110110110011000110001;
    rom[27441] = 25'b1111110110101111001011001;
    rom[27442] = 25'b1111110110101011010000001;
    rom[27443] = 25'b1111110110100111010101000;
    rom[27444] = 25'b1111110110100011011001110;
    rom[27445] = 25'b1111110110011111011110100;
    rom[27446] = 25'b1111110110011011100011001;
    rom[27447] = 25'b1111110110010111100111101;
    rom[27448] = 25'b1111110110010011101100001;
    rom[27449] = 25'b1111110110001111110000100;
    rom[27450] = 25'b1111110110001011110100111;
    rom[27451] = 25'b1111110110000111111001001;
    rom[27452] = 25'b1111110110000011111101010;
    rom[27453] = 25'b1111110110000000000001011;
    rom[27454] = 25'b1111110101111100000101100;
    rom[27455] = 25'b1111110101111000001001011;
    rom[27456] = 25'b1111110101110100001101010;
    rom[27457] = 25'b1111110101110000010001001;
    rom[27458] = 25'b1111110101101100010100111;
    rom[27459] = 25'b1111110101101000011000100;
    rom[27460] = 25'b1111110101100100011100001;
    rom[27461] = 25'b1111110101100000011111101;
    rom[27462] = 25'b1111110101011100100011001;
    rom[27463] = 25'b1111110101011000100110100;
    rom[27464] = 25'b1111110101010100101001110;
    rom[27465] = 25'b1111110101010000101101001;
    rom[27466] = 25'b1111110101001100110000010;
    rom[27467] = 25'b1111110101001000110011011;
    rom[27468] = 25'b1111110101000100110110011;
    rom[27469] = 25'b1111110101000000111001010;
    rom[27470] = 25'b1111110100111100111100010;
    rom[27471] = 25'b1111110100111000111111000;
    rom[27472] = 25'b1111110100110101000001110;
    rom[27473] = 25'b1111110100110001000100100;
    rom[27474] = 25'b1111110100101101000111001;
    rom[27475] = 25'b1111110100101001001001110;
    rom[27476] = 25'b1111110100100101001100001;
    rom[27477] = 25'b1111110100100001001110101;
    rom[27478] = 25'b1111110100011101010001000;
    rom[27479] = 25'b1111110100011001010011010;
    rom[27480] = 25'b1111110100010101010101100;
    rom[27481] = 25'b1111110100010001010111110;
    rom[27482] = 25'b1111110100001101011001110;
    rom[27483] = 25'b1111110100001001011011110;
    rom[27484] = 25'b1111110100000101011101110;
    rom[27485] = 25'b1111110100000001011111101;
    rom[27486] = 25'b1111110011111101100001100;
    rom[27487] = 25'b1111110011111001100011010;
    rom[27488] = 25'b1111110011110101100101000;
    rom[27489] = 25'b1111110011110001100110101;
    rom[27490] = 25'b1111110011101101101000001;
    rom[27491] = 25'b1111110011101001101001110;
    rom[27492] = 25'b1111110011100101101011010;
    rom[27493] = 25'b1111110011100001101100100;
    rom[27494] = 25'b1111110011011101101101111;
    rom[27495] = 25'b1111110011011001101111010;
    rom[27496] = 25'b1111110011010101110000011;
    rom[27497] = 25'b1111110011010001110001100;
    rom[27498] = 25'b1111110011001101110010101;
    rom[27499] = 25'b1111110011001001110011110;
    rom[27500] = 25'b1111110011000101110100101;
    rom[27501] = 25'b1111110011000001110101100;
    rom[27502] = 25'b1111110010111101110110011;
    rom[27503] = 25'b1111110010111001110111001;
    rom[27504] = 25'b1111110010110101111000000;
    rom[27505] = 25'b1111110010110001111000101;
    rom[27506] = 25'b1111110010101101111001010;
    rom[27507] = 25'b1111110010101001111001110;
    rom[27508] = 25'b1111110010100101111010010;
    rom[27509] = 25'b1111110010100001111010110;
    rom[27510] = 25'b1111110010011101111011001;
    rom[27511] = 25'b1111110010011001111011100;
    rom[27512] = 25'b1111110010010101111011110;
    rom[27513] = 25'b1111110010010001111100000;
    rom[27514] = 25'b1111110010001101111100001;
    rom[27515] = 25'b1111110010001001111100010;
    rom[27516] = 25'b1111110010000101111100010;
    rom[27517] = 25'b1111110010000001111100010;
    rom[27518] = 25'b1111110001111101111100010;
    rom[27519] = 25'b1111110001111001111100001;
    rom[27520] = 25'b1111110001110101111100000;
    rom[27521] = 25'b1111110001110001111011110;
    rom[27522] = 25'b1111110001101101111011100;
    rom[27523] = 25'b1111110001101001111011001;
    rom[27524] = 25'b1111110001100101111010111;
    rom[27525] = 25'b1111110001100001111010011;
    rom[27526] = 25'b1111110001011101111001111;
    rom[27527] = 25'b1111110001011001111001011;
    rom[27528] = 25'b1111110001010101111000110;
    rom[27529] = 25'b1111110001010001111000001;
    rom[27530] = 25'b1111110001001101110111100;
    rom[27531] = 25'b1111110001001001110110110;
    rom[27532] = 25'b1111110001000101110110000;
    rom[27533] = 25'b1111110001000001110101001;
    rom[27534] = 25'b1111110000111101110100010;
    rom[27535] = 25'b1111110000111001110011011;
    rom[27536] = 25'b1111110000110101110010011;
    rom[27537] = 25'b1111110000110001110001010;
    rom[27538] = 25'b1111110000101101110000010;
    rom[27539] = 25'b1111110000101001101111001;
    rom[27540] = 25'b1111110000100101101110000;
    rom[27541] = 25'b1111110000100001101100110;
    rom[27542] = 25'b1111110000011101101011011;
    rom[27543] = 25'b1111110000011001101010001;
    rom[27544] = 25'b1111110000010101101000110;
    rom[27545] = 25'b1111110000010001100111011;
    rom[27546] = 25'b1111110000001101100101111;
    rom[27547] = 25'b1111110000001001100100100;
    rom[27548] = 25'b1111110000000101100010111;
    rom[27549] = 25'b1111110000000001100001011;
    rom[27550] = 25'b1111101111111101011111101;
    rom[27551] = 25'b1111101111111001011110000;
    rom[27552] = 25'b1111101111110101011100010;
    rom[27553] = 25'b1111101111110001011010100;
    rom[27554] = 25'b1111101111101101011000101;
    rom[27555] = 25'b1111101111101001010110111;
    rom[27556] = 25'b1111101111100101010101000;
    rom[27557] = 25'b1111101111100001010011000;
    rom[27558] = 25'b1111101111011101010001000;
    rom[27559] = 25'b1111101111011001001111000;
    rom[27560] = 25'b1111101111010101001101000;
    rom[27561] = 25'b1111101111010001001010111;
    rom[27562] = 25'b1111101111001101001000110;
    rom[27563] = 25'b1111101111001001000110100;
    rom[27564] = 25'b1111101111000101000100010;
    rom[27565] = 25'b1111101111000001000010001;
    rom[27566] = 25'b1111101110111100111111110;
    rom[27567] = 25'b1111101110111000111101100;
    rom[27568] = 25'b1111101110110100111011000;
    rom[27569] = 25'b1111101110110000111000101;
    rom[27570] = 25'b1111101110101100110110001;
    rom[27571] = 25'b1111101110101000110011101;
    rom[27572] = 25'b1111101110100100110001001;
    rom[27573] = 25'b1111101110100000101110101;
    rom[27574] = 25'b1111101110011100101100000;
    rom[27575] = 25'b1111101110011000101001011;
    rom[27576] = 25'b1111101110010100100110110;
    rom[27577] = 25'b1111101110010000100100000;
    rom[27578] = 25'b1111101110001100100001010;
    rom[27579] = 25'b1111101110001000011110011;
    rom[27580] = 25'b1111101110000100011011101;
    rom[27581] = 25'b1111101110000000011000110;
    rom[27582] = 25'b1111101101111100010101111;
    rom[27583] = 25'b1111101101111000010011000;
    rom[27584] = 25'b1111101101110100010000000;
    rom[27585] = 25'b1111101101110000001101000;
    rom[27586] = 25'b1111101101101100001010000;
    rom[27587] = 25'b1111101101101000000111000;
    rom[27588] = 25'b1111101101100100000011111;
    rom[27589] = 25'b1111101101100000000000110;
    rom[27590] = 25'b1111101101011011111101101;
    rom[27591] = 25'b1111101101010111111010011;
    rom[27592] = 25'b1111101101010011110111010;
    rom[27593] = 25'b1111101101001111110100000;
    rom[27594] = 25'b1111101101001011110000101;
    rom[27595] = 25'b1111101101000111101101011;
    rom[27596] = 25'b1111101101000011101010001;
    rom[27597] = 25'b1111101100111111100110110;
    rom[27598] = 25'b1111101100111011100011011;
    rom[27599] = 25'b1111101100110111011111111;
    rom[27600] = 25'b1111101100110011011100100;
    rom[27601] = 25'b1111101100101111011000111;
    rom[27602] = 25'b1111101100101011010101100;
    rom[27603] = 25'b1111101100100111010001111;
    rom[27604] = 25'b1111101100100011001110011;
    rom[27605] = 25'b1111101100011111001010110;
    rom[27606] = 25'b1111101100011011000111001;
    rom[27607] = 25'b1111101100010111000011100;
    rom[27608] = 25'b1111101100010010111111111;
    rom[27609] = 25'b1111101100001110111100010;
    rom[27610] = 25'b1111101100001010111000100;
    rom[27611] = 25'b1111101100000110110100110;
    rom[27612] = 25'b1111101100000010110001000;
    rom[27613] = 25'b1111101011111110101101001;
    rom[27614] = 25'b1111101011111010101001011;
    rom[27615] = 25'b1111101011110110100101101;
    rom[27616] = 25'b1111101011110010100001101;
    rom[27617] = 25'b1111101011101110011101110;
    rom[27618] = 25'b1111101011101010011001111;
    rom[27619] = 25'b1111101011100110010110000;
    rom[27620] = 25'b1111101011100010010010000;
    rom[27621] = 25'b1111101011011110001110000;
    rom[27622] = 25'b1111101011011010001010000;
    rom[27623] = 25'b1111101011010110000110000;
    rom[27624] = 25'b1111101011010010000010000;
    rom[27625] = 25'b1111101011001101111110000;
    rom[27626] = 25'b1111101011001001111001111;
    rom[27627] = 25'b1111101011000101110101110;
    rom[27628] = 25'b1111101011000001110001110;
    rom[27629] = 25'b1111101010111101101101100;
    rom[27630] = 25'b1111101010111001101001011;
    rom[27631] = 25'b1111101010110101100101001;
    rom[27632] = 25'b1111101010110001100001000;
    rom[27633] = 25'b1111101010101101011100111;
    rom[27634] = 25'b1111101010101001011000100;
    rom[27635] = 25'b1111101010100101010100011;
    rom[27636] = 25'b1111101010100001010000001;
    rom[27637] = 25'b1111101010011101001011111;
    rom[27638] = 25'b1111101010011001000111101;
    rom[27639] = 25'b1111101010010101000011010;
    rom[27640] = 25'b1111101010010000111110111;
    rom[27641] = 25'b1111101010001100111010101;
    rom[27642] = 25'b1111101010001000110110010;
    rom[27643] = 25'b1111101010000100110001111;
    rom[27644] = 25'b1111101010000000101101100;
    rom[27645] = 25'b1111101001111100101001001;
    rom[27646] = 25'b1111101001111000100100101;
    rom[27647] = 25'b1111101001110100100000010;
    rom[27648] = 25'b1111101001110000011011111;
    rom[27649] = 25'b1111101001101100010111011;
    rom[27650] = 25'b1111101001101000010010111;
    rom[27651] = 25'b1111101001100100001110100;
    rom[27652] = 25'b1111101001100000001010000;
    rom[27653] = 25'b1111101001011100000101100;
    rom[27654] = 25'b1111101001011000000001000;
    rom[27655] = 25'b1111101001010011111100100;
    rom[27656] = 25'b1111101001001111111000000;
    rom[27657] = 25'b1111101001001011110011100;
    rom[27658] = 25'b1111101001000111101110111;
    rom[27659] = 25'b1111101001000011101010011;
    rom[27660] = 25'b1111101000111111100101110;
    rom[27661] = 25'b1111101000111011100001010;
    rom[27662] = 25'b1111101000110111011100110;
    rom[27663] = 25'b1111101000110011011000000;
    rom[27664] = 25'b1111101000101111010011100;
    rom[27665] = 25'b1111101000101011001110111;
    rom[27666] = 25'b1111101000100111001010011;
    rom[27667] = 25'b1111101000100011000101101;
    rom[27668] = 25'b1111101000011111000001000;
    rom[27669] = 25'b1111101000011010111100100;
    rom[27670] = 25'b1111101000010110110111111;
    rom[27671] = 25'b1111101000010010110011010;
    rom[27672] = 25'b1111101000001110101110100;
    rom[27673] = 25'b1111101000001010101001111;
    rom[27674] = 25'b1111101000000110100101010;
    rom[27675] = 25'b1111101000000010100000101;
    rom[27676] = 25'b1111100111111110011100000;
    rom[27677] = 25'b1111100111111010010111011;
    rom[27678] = 25'b1111100111110110010010110;
    rom[27679] = 25'b1111100111110010001110000;
    rom[27680] = 25'b1111100111101110001001011;
    rom[27681] = 25'b1111100111101010000100101;
    rom[27682] = 25'b1111100111100110000000000;
    rom[27683] = 25'b1111100111100001111011011;
    rom[27684] = 25'b1111100111011101110110110;
    rom[27685] = 25'b1111100111011001110010000;
    rom[27686] = 25'b1111100111010101101101011;
    rom[27687] = 25'b1111100111010001101000110;
    rom[27688] = 25'b1111100111001101100100001;
    rom[27689] = 25'b1111100111001001011111011;
    rom[27690] = 25'b1111100111000101011010110;
    rom[27691] = 25'b1111100111000001010110000;
    rom[27692] = 25'b1111100110111101010001011;
    rom[27693] = 25'b1111100110111001001100110;
    rom[27694] = 25'b1111100110110101001000001;
    rom[27695] = 25'b1111100110110001000011100;
    rom[27696] = 25'b1111100110101100111110111;
    rom[27697] = 25'b1111100110101000111010010;
    rom[27698] = 25'b1111100110100100110101100;
    rom[27699] = 25'b1111100110100000110000111;
    rom[27700] = 25'b1111100110011100101100010;
    rom[27701] = 25'b1111100110011000100111101;
    rom[27702] = 25'b1111100110010100100011001;
    rom[27703] = 25'b1111100110010000011110011;
    rom[27704] = 25'b1111100110001100011001110;
    rom[27705] = 25'b1111100110001000010101010;
    rom[27706] = 25'b1111100110000100010000101;
    rom[27707] = 25'b1111100110000000001100000;
    rom[27708] = 25'b1111100101111100000111100;
    rom[27709] = 25'b1111100101111000000010111;
    rom[27710] = 25'b1111100101110011111110010;
    rom[27711] = 25'b1111100101101111111001110;
    rom[27712] = 25'b1111100101101011110101010;
    rom[27713] = 25'b1111100101100111110000110;
    rom[27714] = 25'b1111100101100011101100010;
    rom[27715] = 25'b1111100101011111100111101;
    rom[27716] = 25'b1111100101011011100011010;
    rom[27717] = 25'b1111100101010111011110101;
    rom[27718] = 25'b1111100101010011011010001;
    rom[27719] = 25'b1111100101001111010101110;
    rom[27720] = 25'b1111100101001011010001010;
    rom[27721] = 25'b1111100101000111001100111;
    rom[27722] = 25'b1111100101000011001000011;
    rom[27723] = 25'b1111100100111111000100000;
    rom[27724] = 25'b1111100100111010111111100;
    rom[27725] = 25'b1111100100110110111011001;
    rom[27726] = 25'b1111100100110010110110110;
    rom[27727] = 25'b1111100100101110110010100;
    rom[27728] = 25'b1111100100101010101110001;
    rom[27729] = 25'b1111100100100110101001110;
    rom[27730] = 25'b1111100100100010100101011;
    rom[27731] = 25'b1111100100011110100001001;
    rom[27732] = 25'b1111100100011010011100111;
    rom[27733] = 25'b1111100100010110011000100;
    rom[27734] = 25'b1111100100010010010100010;
    rom[27735] = 25'b1111100100001110010000000;
    rom[27736] = 25'b1111100100001010001011111;
    rom[27737] = 25'b1111100100000110000111101;
    rom[27738] = 25'b1111100100000010000011011;
    rom[27739] = 25'b1111100011111101111111010;
    rom[27740] = 25'b1111100011111001111011001;
    rom[27741] = 25'b1111100011110101110111000;
    rom[27742] = 25'b1111100011110001110010111;
    rom[27743] = 25'b1111100011101101101110110;
    rom[27744] = 25'b1111100011101001101010110;
    rom[27745] = 25'b1111100011100101100110101;
    rom[27746] = 25'b1111100011100001100010101;
    rom[27747] = 25'b1111100011011101011110100;
    rom[27748] = 25'b1111100011011001011010100;
    rom[27749] = 25'b1111100011010101010110101;
    rom[27750] = 25'b1111100011010001010010101;
    rom[27751] = 25'b1111100011001101001110110;
    rom[27752] = 25'b1111100011001001001010111;
    rom[27753] = 25'b1111100011000101000111000;
    rom[27754] = 25'b1111100011000001000011001;
    rom[27755] = 25'b1111100010111100111111010;
    rom[27756] = 25'b1111100010111000111011100;
    rom[27757] = 25'b1111100010110100110111101;
    rom[27758] = 25'b1111100010110000110100000;
    rom[27759] = 25'b1111100010101100110000010;
    rom[27760] = 25'b1111100010101000101100100;
    rom[27761] = 25'b1111100010100100101000111;
    rom[27762] = 25'b1111100010100000100101010;
    rom[27763] = 25'b1111100010011100100001101;
    rom[27764] = 25'b1111100010011000011110000;
    rom[27765] = 25'b1111100010010100011010011;
    rom[27766] = 25'b1111100010010000010110111;
    rom[27767] = 25'b1111100010001100010011011;
    rom[27768] = 25'b1111100010001000001111111;
    rom[27769] = 25'b1111100010000100001100011;
    rom[27770] = 25'b1111100010000000001001000;
    rom[27771] = 25'b1111100001111100000101101;
    rom[27772] = 25'b1111100001111000000010010;
    rom[27773] = 25'b1111100001110011111110111;
    rom[27774] = 25'b1111100001101111111011101;
    rom[27775] = 25'b1111100001101011111000010;
    rom[27776] = 25'b1111100001100111110101000;
    rom[27777] = 25'b1111100001100011110001111;
    rom[27778] = 25'b1111100001011111101110101;
    rom[27779] = 25'b1111100001011011101011100;
    rom[27780] = 25'b1111100001010111101000100;
    rom[27781] = 25'b1111100001010011100101010;
    rom[27782] = 25'b1111100001001111100010010;
    rom[27783] = 25'b1111100001001011011111010;
    rom[27784] = 25'b1111100001000111011100010;
    rom[27785] = 25'b1111100001000011011001011;
    rom[27786] = 25'b1111100000111111010110011;
    rom[27787] = 25'b1111100000111011010011100;
    rom[27788] = 25'b1111100000110111010000101;
    rom[27789] = 25'b1111100000110011001101111;
    rom[27790] = 25'b1111100000101111001011001;
    rom[27791] = 25'b1111100000101011001000011;
    rom[27792] = 25'b1111100000100111000101101;
    rom[27793] = 25'b1111100000100011000011000;
    rom[27794] = 25'b1111100000011111000000011;
    rom[27795] = 25'b1111100000011010111101110;
    rom[27796] = 25'b1111100000010110111011010;
    rom[27797] = 25'b1111100000010010111000110;
    rom[27798] = 25'b1111100000001110110110010;
    rom[27799] = 25'b1111100000001010110011111;
    rom[27800] = 25'b1111100000000110110001100;
    rom[27801] = 25'b1111100000000010101111001;
    rom[27802] = 25'b1111011111111110101100111;
    rom[27803] = 25'b1111011111111010101010101;
    rom[27804] = 25'b1111011111110110101000011;
    rom[27805] = 25'b1111011111110010100110001;
    rom[27806] = 25'b1111011111101110100100000;
    rom[27807] = 25'b1111011111101010100001111;
    rom[27808] = 25'b1111011111100110011111111;
    rom[27809] = 25'b1111011111100010011101111;
    rom[27810] = 25'b1111011111011110011011111;
    rom[27811] = 25'b1111011111011010011010000;
    rom[27812] = 25'b1111011111010110011000001;
    rom[27813] = 25'b1111011111010010010110010;
    rom[27814] = 25'b1111011111001110010100100;
    rom[27815] = 25'b1111011111001010010010110;
    rom[27816] = 25'b1111011111000110010001000;
    rom[27817] = 25'b1111011111000010001111011;
    rom[27818] = 25'b1111011110111110001101110;
    rom[27819] = 25'b1111011110111010001100001;
    rom[27820] = 25'b1111011110110110001010110;
    rom[27821] = 25'b1111011110110010001001010;
    rom[27822] = 25'b1111011110101110000111110;
    rom[27823] = 25'b1111011110101010000110011;
    rom[27824] = 25'b1111011110100110000101001;
    rom[27825] = 25'b1111011110100010000011111;
    rom[27826] = 25'b1111011110011110000010100;
    rom[27827] = 25'b1111011110011010000001100;
    rom[27828] = 25'b1111011110010110000000010;
    rom[27829] = 25'b1111011110010001111111001;
    rom[27830] = 25'b1111011110001101111110001;
    rom[27831] = 25'b1111011110001001111101001;
    rom[27832] = 25'b1111011110000101111100010;
    rom[27833] = 25'b1111011110000001111011100;
    rom[27834] = 25'b1111011101111101111010101;
    rom[27835] = 25'b1111011101111001111001111;
    rom[27836] = 25'b1111011101110101111001001;
    rom[27837] = 25'b1111011101110001111000100;
    rom[27838] = 25'b1111011101101101110111111;
    rom[27839] = 25'b1111011101101001110111010;
    rom[27840] = 25'b1111011101100101110110110;
    rom[27841] = 25'b1111011101100001110110011;
    rom[27842] = 25'b1111011101011101110110000;
    rom[27843] = 25'b1111011101011001110101101;
    rom[27844] = 25'b1111011101010101110101011;
    rom[27845] = 25'b1111011101010001110101001;
    rom[27846] = 25'b1111011101001101110101000;
    rom[27847] = 25'b1111011101001001110100110;
    rom[27848] = 25'b1111011101000101110100111;
    rom[27849] = 25'b1111011101000001110100110;
    rom[27850] = 25'b1111011100111101110100111;
    rom[27851] = 25'b1111011100111001110101000;
    rom[27852] = 25'b1111011100110101110101001;
    rom[27853] = 25'b1111011100110001110101011;
    rom[27854] = 25'b1111011100101101110101110;
    rom[27855] = 25'b1111011100101001110110000;
    rom[27856] = 25'b1111011100100101110110100;
    rom[27857] = 25'b1111011100100001110110111;
    rom[27858] = 25'b1111011100011101110111100;
    rom[27859] = 25'b1111011100011001111000001;
    rom[27860] = 25'b1111011100010101111000110;
    rom[27861] = 25'b1111011100010001111001100;
    rom[27862] = 25'b1111011100001101111010010;
    rom[27863] = 25'b1111011100001001111011001;
    rom[27864] = 25'b1111011100000101111100001;
    rom[27865] = 25'b1111011100000001111101000;
    rom[27866] = 25'b1111011011111101111110001;
    rom[27867] = 25'b1111011011111001111111001;
    rom[27868] = 25'b1111011011110110000000010;
    rom[27869] = 25'b1111011011110010000001100;
    rom[27870] = 25'b1111011011101110000010111;
    rom[27871] = 25'b1111011011101010000100010;
    rom[27872] = 25'b1111011011100110000101101;
    rom[27873] = 25'b1111011011100010000111001;
    rom[27874] = 25'b1111011011011110001000101;
    rom[27875] = 25'b1111011011011010001010010;
    rom[27876] = 25'b1111011011010110001100000;
    rom[27877] = 25'b1111011011010010001101110;
    rom[27878] = 25'b1111011011001110001111101;
    rom[27879] = 25'b1111011011001010010001100;
    rom[27880] = 25'b1111011011000110010011100;
    rom[27881] = 25'b1111011011000010010101100;
    rom[27882] = 25'b1111011010111110010111101;
    rom[27883] = 25'b1111011010111010011001110;
    rom[27884] = 25'b1111011010110110011100001;
    rom[27885] = 25'b1111011010110010011110011;
    rom[27886] = 25'b1111011010101110100000110;
    rom[27887] = 25'b1111011010101010100011010;
    rom[27888] = 25'b1111011010100110100101110;
    rom[27889] = 25'b1111011010100010101000011;
    rom[27890] = 25'b1111011010011110101011000;
    rom[27891] = 25'b1111011010011010101101110;
    rom[27892] = 25'b1111011010010110110000100;
    rom[27893] = 25'b1111011010010010110011100;
    rom[27894] = 25'b1111011010001110110110100;
    rom[27895] = 25'b1111011010001010111001100;
    rom[27896] = 25'b1111011010000110111100101;
    rom[27897] = 25'b1111011010000010111111110;
    rom[27898] = 25'b1111011001111111000011001;
    rom[27899] = 25'b1111011001111011000110011;
    rom[27900] = 25'b1111011001110111001001111;
    rom[27901] = 25'b1111011001110011001101011;
    rom[27902] = 25'b1111011001101111010000111;
    rom[27903] = 25'b1111011001101011010100101;
    rom[27904] = 25'b1111011001100111011000010;
    rom[27905] = 25'b1111011001100011011100001;
    rom[27906] = 25'b1111011001011111100000000;
    rom[27907] = 25'b1111011001011011100011111;
    rom[27908] = 25'b1111011001010111101000000;
    rom[27909] = 25'b1111011001010011101100001;
    rom[27910] = 25'b1111011001001111110000011;
    rom[27911] = 25'b1111011001001011110100101;
    rom[27912] = 25'b1111011001000111111001000;
    rom[27913] = 25'b1111011001000011111101011;
    rom[27914] = 25'b1111011001000000000001111;
    rom[27915] = 25'b1111011000111100000110100;
    rom[27916] = 25'b1111011000111000001011010;
    rom[27917] = 25'b1111011000110100010000000;
    rom[27918] = 25'b1111011000110000010100111;
    rom[27919] = 25'b1111011000101100011001111;
    rom[27920] = 25'b1111011000101000011110111;
    rom[27921] = 25'b1111011000100100100011111;
    rom[27922] = 25'b1111011000100000101001001;
    rom[27923] = 25'b1111011000011100101110011;
    rom[27924] = 25'b1111011000011000110011110;
    rom[27925] = 25'b1111011000010100111001001;
    rom[27926] = 25'b1111011000010000111110110;
    rom[27927] = 25'b1111011000001101000100011;
    rom[27928] = 25'b1111011000001001001010001;
    rom[27929] = 25'b1111011000000101001111110;
    rom[27930] = 25'b1111011000000001010101110;
    rom[27931] = 25'b1111010111111101011011110;
    rom[27932] = 25'b1111010111111001100001110;
    rom[27933] = 25'b1111010111110101100111111;
    rom[27934] = 25'b1111010111110001101110001;
    rom[27935] = 25'b1111010111101101110100011;
    rom[27936] = 25'b1111010111101001111010111;
    rom[27937] = 25'b1111010111100110000001011;
    rom[27938] = 25'b1111010111100010000111111;
    rom[27939] = 25'b1111010111011110001110100;
    rom[27940] = 25'b1111010111011010010101011;
    rom[27941] = 25'b1111010111010110011100010;
    rom[27942] = 25'b1111010111010010100011001;
    rom[27943] = 25'b1111010111001110101010010;
    rom[27944] = 25'b1111010111001010110001010;
    rom[27945] = 25'b1111010111000110111000100;
    rom[27946] = 25'b1111010111000010111111111;
    rom[27947] = 25'b1111010110111111000111011;
    rom[27948] = 25'b1111010110111011001110111;
    rom[27949] = 25'b1111010110110111010110011;
    rom[27950] = 25'b1111010110110011011110001;
    rom[27951] = 25'b1111010110101111100101111;
    rom[27952] = 25'b1111010110101011101101111;
    rom[27953] = 25'b1111010110100111110101111;
    rom[27954] = 25'b1111010110100011111101111;
    rom[27955] = 25'b1111010110100000000110000;
    rom[27956] = 25'b1111010110011100001110011;
    rom[27957] = 25'b1111010110011000010110110;
    rom[27958] = 25'b1111010110010100011111001;
    rom[27959] = 25'b1111010110010000100111110;
    rom[27960] = 25'b1111010110001100110000011;
    rom[27961] = 25'b1111010110001000111001001;
    rom[27962] = 25'b1111010110000101000010001;
    rom[27963] = 25'b1111010110000001001011000;
    rom[27964] = 25'b1111010101111101010100000;
    rom[27965] = 25'b1111010101111001011101010;
    rom[27966] = 25'b1111010101110101100110100;
    rom[27967] = 25'b1111010101110001101111111;
    rom[27968] = 25'b1111010101101101111001011;
    rom[27969] = 25'b1111010101101010000010111;
    rom[27970] = 25'b1111010101100110001100100;
    rom[27971] = 25'b1111010101100010010110011;
    rom[27972] = 25'b1111010101011110100000001;
    rom[27973] = 25'b1111010101011010101010010;
    rom[27974] = 25'b1111010101010110110100011;
    rom[27975] = 25'b1111010101010010111110011;
    rom[27976] = 25'b1111010101001111001000110;
    rom[27977] = 25'b1111010101001011010011001;
    rom[27978] = 25'b1111010101000111011101110;
    rom[27979] = 25'b1111010101000011101000010;
    rom[27980] = 25'b1111010100111111110011000;
    rom[27981] = 25'b1111010100111011111101110;
    rom[27982] = 25'b1111010100111000001000101;
    rom[27983] = 25'b1111010100110100010011110;
    rom[27984] = 25'b1111010100110000011110111;
    rom[27985] = 25'b1111010100101100101010001;
    rom[27986] = 25'b1111010100101000110101100;
    rom[27987] = 25'b1111010100100101000000111;
    rom[27988] = 25'b1111010100100001001100100;
    rom[27989] = 25'b1111010100011101011000010;
    rom[27990] = 25'b1111010100011001100100000;
    rom[27991] = 25'b1111010100010101101111111;
    rom[27992] = 25'b1111010100010001111011111;
    rom[27993] = 25'b1111010100001110001000000;
    rom[27994] = 25'b1111010100001010010100010;
    rom[27995] = 25'b1111010100000110100000101;
    rom[27996] = 25'b1111010100000010101101001;
    rom[27997] = 25'b1111010011111110111001101;
    rom[27998] = 25'b1111010011111011000110010;
    rom[27999] = 25'b1111010011110111010011001;
    rom[28000] = 25'b1111010011110011100000000;
    rom[28001] = 25'b1111010011101111101101000;
    rom[28002] = 25'b1111010011101011111010010;
    rom[28003] = 25'b1111010011101000000111011;
    rom[28004] = 25'b1111010011100100010100110;
    rom[28005] = 25'b1111010011100000100010010;
    rom[28006] = 25'b1111010011011100101111111;
    rom[28007] = 25'b1111010011011000111101101;
    rom[28008] = 25'b1111010011010101001011011;
    rom[28009] = 25'b1111010011010001011001011;
    rom[28010] = 25'b1111010011001101100111011;
    rom[28011] = 25'b1111010011001001110101101;
    rom[28012] = 25'b1111010011000110000011111;
    rom[28013] = 25'b1111010011000010010010011;
    rom[28014] = 25'b1111010010111110100000111;
    rom[28015] = 25'b1111010010111010101111100;
    rom[28016] = 25'b1111010010110110111110010;
    rom[28017] = 25'b1111010010110011001101010;
    rom[28018] = 25'b1111010010101111011100001;
    rom[28019] = 25'b1111010010101011101011011;
    rom[28020] = 25'b1111010010100111111010101;
    rom[28021] = 25'b1111010010100100001001111;
    rom[28022] = 25'b1111010010100000011001100;
    rom[28023] = 25'b1111010010011100101001001;
    rom[28024] = 25'b1111010010011000111000110;
    rom[28025] = 25'b1111010010010101001000101;
    rom[28026] = 25'b1111010010010001011000101;
    rom[28027] = 25'b1111010010001101101000110;
    rom[28028] = 25'b1111010010001001111001000;
    rom[28029] = 25'b1111010010000110001001011;
    rom[28030] = 25'b1111010010000010011001111;
    rom[28031] = 25'b1111010001111110101010011;
    rom[28032] = 25'b1111010001111010111011001;
    rom[28033] = 25'b1111010001110111001100000;
    rom[28034] = 25'b1111010001110011011101000;
    rom[28035] = 25'b1111010001101111101110001;
    rom[28036] = 25'b1111010001101011111111011;
    rom[28037] = 25'b1111010001101000010000110;
    rom[28038] = 25'b1111010001100100100010010;
    rom[28039] = 25'b1111010001100000110011111;
    rom[28040] = 25'b1111010001011101000101101;
    rom[28041] = 25'b1111010001011001010111100;
    rom[28042] = 25'b1111010001010101101001100;
    rom[28043] = 25'b1111010001010001111011101;
    rom[28044] = 25'b1111010001001110001101111;
    rom[28045] = 25'b1111010001001010100000010;
    rom[28046] = 25'b1111010001000110110010111;
    rom[28047] = 25'b1111010001000011000101100;
    rom[28048] = 25'b1111010000111111011000011;
    rom[28049] = 25'b1111010000111011101011010;
    rom[28050] = 25'b1111010000110111111110010;
    rom[28051] = 25'b1111010000110100010001100;
    rom[28052] = 25'b1111010000110000100100111;
    rom[28053] = 25'b1111010000101100111000010;
    rom[28054] = 25'b1111010000101001001011111;
    rom[28055] = 25'b1111010000100101011111100;
    rom[28056] = 25'b1111010000100001110011011;
    rom[28057] = 25'b1111010000011110000111011;
    rom[28058] = 25'b1111010000011010011011100;
    rom[28059] = 25'b1111010000010110101111110;
    rom[28060] = 25'b1111010000010011000100001;
    rom[28061] = 25'b1111010000001111011000110;
    rom[28062] = 25'b1111010000001011101101011;
    rom[28063] = 25'b1111010000001000000010010;
    rom[28064] = 25'b1111010000000100010111010;
    rom[28065] = 25'b1111010000000000101100010;
    rom[28066] = 25'b1111001111111101000001100;
    rom[28067] = 25'b1111001111111001010110111;
    rom[28068] = 25'b1111001111110101101100010;
    rom[28069] = 25'b1111001111110010000010000;
    rom[28070] = 25'b1111001111101110010111110;
    rom[28071] = 25'b1111001111101010101101101;
    rom[28072] = 25'b1111001111100111000011110;
    rom[28073] = 25'b1111001111100011011010000;
    rom[28074] = 25'b1111001111011111110000010;
    rom[28075] = 25'b1111001111011100000110110;
    rom[28076] = 25'b1111001111011000011101011;
    rom[28077] = 25'b1111001111010100110100001;
    rom[28078] = 25'b1111001111010001001011001;
    rom[28079] = 25'b1111001111001101100010001;
    rom[28080] = 25'b1111001111001001111001010;
    rom[28081] = 25'b1111001111000110010000101;
    rom[28082] = 25'b1111001111000010101000001;
    rom[28083] = 25'b1111001110111110111111110;
    rom[28084] = 25'b1111001110111011010111100;
    rom[28085] = 25'b1111001110110111101111100;
    rom[28086] = 25'b1111001110110100000111100;
    rom[28087] = 25'b1111001110110000011111110;
    rom[28088] = 25'b1111001110101100111000001;
    rom[28089] = 25'b1111001110101001010000101;
    rom[28090] = 25'b1111001110100101101001010;
    rom[28091] = 25'b1111001110100010000010000;
    rom[28092] = 25'b1111001110011110011011000;
    rom[28093] = 25'b1111001110011010110100001;
    rom[28094] = 25'b1111001110010111001101011;
    rom[28095] = 25'b1111001110010011100110110;
    rom[28096] = 25'b1111001110010000000000011;
    rom[28097] = 25'b1111001110001100011010000;
    rom[28098] = 25'b1111001110001000110011111;
    rom[28099] = 25'b1111001110000101001101111;
    rom[28100] = 25'b1111001110000001101000000;
    rom[28101] = 25'b1111001101111110000010010;
    rom[28102] = 25'b1111001101111010011100110;
    rom[28103] = 25'b1111001101110110110111011;
    rom[28104] = 25'b1111001101110011010010001;
    rom[28105] = 25'b1111001101101111101101000;
    rom[28106] = 25'b1111001101101100001000000;
    rom[28107] = 25'b1111001101101000100011011;
    rom[28108] = 25'b1111001101100100111110101;
    rom[28109] = 25'b1111001101100001011010010;
    rom[28110] = 25'b1111001101011101110101111;
    rom[28111] = 25'b1111001101011010010001110;
    rom[28112] = 25'b1111001101010110101101101;
    rom[28113] = 25'b1111001101010011001001110;
    rom[28114] = 25'b1111001101001111100110001;
    rom[28115] = 25'b1111001101001100000010101;
    rom[28116] = 25'b1111001101001000011111010;
    rom[28117] = 25'b1111001101000100111100000;
    rom[28118] = 25'b1111001101000001011000111;
    rom[28119] = 25'b1111001100111101110110000;
    rom[28120] = 25'b1111001100111010010011010;
    rom[28121] = 25'b1111001100110110110000101;
    rom[28122] = 25'b1111001100110011001110010;
    rom[28123] = 25'b1111001100101111101100000;
    rom[28124] = 25'b1111001100101100001001111;
    rom[28125] = 25'b1111001100101000101000000;
    rom[28126] = 25'b1111001100100101000110001;
    rom[28127] = 25'b1111001100100001100100100;
    rom[28128] = 25'b1111001100011110000011000;
    rom[28129] = 25'b1111001100011010100001110;
    rom[28130] = 25'b1111001100010111000000101;
    rom[28131] = 25'b1111001100010011011111101;
    rom[28132] = 25'b1111001100001111111110111;
    rom[28133] = 25'b1111001100001100011110001;
    rom[28134] = 25'b1111001100001000111101101;
    rom[28135] = 25'b1111001100000101011101011;
    rom[28136] = 25'b1111001100000001111101010;
    rom[28137] = 25'b1111001011111110011101001;
    rom[28138] = 25'b1111001011111010111101010;
    rom[28139] = 25'b1111001011110111011101101;
    rom[28140] = 25'b1111001011110011111110001;
    rom[28141] = 25'b1111001011110000011110111;
    rom[28142] = 25'b1111001011101100111111110;
    rom[28143] = 25'b1111001011101001100000101;
    rom[28144] = 25'b1111001011100110000001111;
    rom[28145] = 25'b1111001011100010100011010;
    rom[28146] = 25'b1111001011011111000100101;
    rom[28147] = 25'b1111001011011011100110011;
    rom[28148] = 25'b1111001011011000001000010;
    rom[28149] = 25'b1111001011010100101010010;
    rom[28150] = 25'b1111001011010001001100100;
    rom[28151] = 25'b1111001011001101101110110;
    rom[28152] = 25'b1111001011001010010001011;
    rom[28153] = 25'b1111001011000110110100000;
    rom[28154] = 25'b1111001011000011010110111;
    rom[28155] = 25'b1111001010111111111001111;
    rom[28156] = 25'b1111001010111100011101001;
    rom[28157] = 25'b1111001010111001000000101;
    rom[28158] = 25'b1111001010110101100100001;
    rom[28159] = 25'b1111001010110010000111111;
    rom[28160] = 25'b1111001010101110101011110;
    rom[28161] = 25'b1111001010101011001111111;
    rom[28162] = 25'b1111001010100111110100001;
    rom[28163] = 25'b1111001010100100011000101;
    rom[28164] = 25'b1111001010100000111101001;
    rom[28165] = 25'b1111001010011101100001111;
    rom[28166] = 25'b1111001010011010000110111;
    rom[28167] = 25'b1111001010010110101100000;
    rom[28168] = 25'b1111001010010011010001011;
    rom[28169] = 25'b1111001010001111110110110;
    rom[28170] = 25'b1111001010001100011100100;
    rom[28171] = 25'b1111001010001001000010010;
    rom[28172] = 25'b1111001010000101101000011;
    rom[28173] = 25'b1111001010000010001110100;
    rom[28174] = 25'b1111001001111110110101000;
    rom[28175] = 25'b1111001001111011011011101;
    rom[28176] = 25'b1111001001111000000010010;
    rom[28177] = 25'b1111001001110100101001010;
    rom[28178] = 25'b1111001001110001010000010;
    rom[28179] = 25'b1111001001101101110111100;
    rom[28180] = 25'b1111001001101010011111000;
    rom[28181] = 25'b1111001001100111000110101;
    rom[28182] = 25'b1111001001100011101110100;
    rom[28183] = 25'b1111001001100000010110101;
    rom[28184] = 25'b1111001001011100111110110;
    rom[28185] = 25'b1111001001011001100111001;
    rom[28186] = 25'b1111001001010110001111110;
    rom[28187] = 25'b1111001001010010111000011;
    rom[28188] = 25'b1111001001001111100001011;
    rom[28189] = 25'b1111001001001100001010100;
    rom[28190] = 25'b1111001001001000110011110;
    rom[28191] = 25'b1111001001000101011101010;
    rom[28192] = 25'b1111001001000010000111000;
    rom[28193] = 25'b1111001000111110110000110;
    rom[28194] = 25'b1111001000111011011010111;
    rom[28195] = 25'b1111001000111000000101001;
    rom[28196] = 25'b1111001000110100101111100;
    rom[28197] = 25'b1111001000110001011010001;
    rom[28198] = 25'b1111001000101110000100111;
    rom[28199] = 25'b1111001000101010101111111;
    rom[28200] = 25'b1111001000100111011011001;
    rom[28201] = 25'b1111001000100100000110100;
    rom[28202] = 25'b1111001000100000110010000;
    rom[28203] = 25'b1111001000011101011101110;
    rom[28204] = 25'b1111001000011010001001101;
    rom[28205] = 25'b1111001000010110110101110;
    rom[28206] = 25'b1111001000010011100010001;
    rom[28207] = 25'b1111001000010000001110101;
    rom[28208] = 25'b1111001000001100111011010;
    rom[28209] = 25'b1111001000001001101000010;
    rom[28210] = 25'b1111001000000110010101010;
    rom[28211] = 25'b1111001000000011000010101;
    rom[28212] = 25'b1111000111111111110000000;
    rom[28213] = 25'b1111000111111100011101101;
    rom[28214] = 25'b1111000111111001001011100;
    rom[28215] = 25'b1111000111110101111001101;
    rom[28216] = 25'b1111000111110010100111111;
    rom[28217] = 25'b1111000111101111010110011;
    rom[28218] = 25'b1111000111101100000101000;
    rom[28219] = 25'b1111000111101000110011110;
    rom[28220] = 25'b1111000111100101100010111;
    rom[28221] = 25'b1111000111100010010010000;
    rom[28222] = 25'b1111000111011111000001100;
    rom[28223] = 25'b1111000111011011110001001;
    rom[28224] = 25'b1111000111011000100000111;
    rom[28225] = 25'b1111000111010101010000111;
    rom[28226] = 25'b1111000111010010000001001;
    rom[28227] = 25'b1111000111001110110001100;
    rom[28228] = 25'b1111000111001011100010010;
    rom[28229] = 25'b1111000111001000010011000;
    rom[28230] = 25'b1111000111000101000100000;
    rom[28231] = 25'b1111000111000001110101010;
    rom[28232] = 25'b1111000110111110100110110;
    rom[28233] = 25'b1111000110111011011000011;
    rom[28234] = 25'b1111000110111000001010001;
    rom[28235] = 25'b1111000110110100111100001;
    rom[28236] = 25'b1111000110110001101110011;
    rom[28237] = 25'b1111000110101110100000111;
    rom[28238] = 25'b1111000110101011010011100;
    rom[28239] = 25'b1111000110101000000110011;
    rom[28240] = 25'b1111000110100100111001011;
    rom[28241] = 25'b1111000110100001101100101;
    rom[28242] = 25'b1111000110011110100000000;
    rom[28243] = 25'b1111000110011011010011110;
    rom[28244] = 25'b1111000110011000000111100;
    rom[28245] = 25'b1111000110010100111011101;
    rom[28246] = 25'b1111000110010001101111111;
    rom[28247] = 25'b1111000110001110100100011;
    rom[28248] = 25'b1111000110001011011001001;
    rom[28249] = 25'b1111000110001000001110000;
    rom[28250] = 25'b1111000110000101000011001;
    rom[28251] = 25'b1111000110000001111000011;
    rom[28252] = 25'b1111000101111110101110000;
    rom[28253] = 25'b1111000101111011100011101;
    rom[28254] = 25'b1111000101111000011001101;
    rom[28255] = 25'b1111000101110101001111110;
    rom[28256] = 25'b1111000101110010000110001;
    rom[28257] = 25'b1111000101101110111100110;
    rom[28258] = 25'b1111000101101011110011100;
    rom[28259] = 25'b1111000101101000101010100;
    rom[28260] = 25'b1111000101100101100001110;
    rom[28261] = 25'b1111000101100010011001001;
    rom[28262] = 25'b1111000101011111010000110;
    rom[28263] = 25'b1111000101011100001000101;
    rom[28264] = 25'b1111000101011001000000101;
    rom[28265] = 25'b1111000101010101111000111;
    rom[28266] = 25'b1111000101010010110001011;
    rom[28267] = 25'b1111000101001111101010001;
    rom[28268] = 25'b1111000101001100100011000;
    rom[28269] = 25'b1111000101001001011100001;
    rom[28270] = 25'b1111000101000110010101100;
    rom[28271] = 25'b1111000101000011001111000;
    rom[28272] = 25'b1111000101000000001000110;
    rom[28273] = 25'b1111000100111101000010110;
    rom[28274] = 25'b1111000100111001111101000;
    rom[28275] = 25'b1111000100110110110111011;
    rom[28276] = 25'b1111000100110011110010001;
    rom[28277] = 25'b1111000100110000101100111;
    rom[28278] = 25'b1111000100101101101000000;
    rom[28279] = 25'b1111000100101010100011010;
    rom[28280] = 25'b1111000100100111011110111;
    rom[28281] = 25'b1111000100100100011010101;
    rom[28282] = 25'b1111000100100001010110100;
    rom[28283] = 25'b1111000100011110010010101;
    rom[28284] = 25'b1111000100011011001111001;
    rom[28285] = 25'b1111000100011000001011110;
    rom[28286] = 25'b1111000100010101001000101;
    rom[28287] = 25'b1111000100010010000101101;
    rom[28288] = 25'b1111000100001111000010111;
    rom[28289] = 25'b1111000100001100000000011;
    rom[28290] = 25'b1111000100001000111110001;
    rom[28291] = 25'b1111000100000101111100001;
    rom[28292] = 25'b1111000100000010111010010;
    rom[28293] = 25'b1111000011111111111000101;
    rom[28294] = 25'b1111000011111100110111010;
    rom[28295] = 25'b1111000011111001110110001;
    rom[28296] = 25'b1111000011110110110101010;
    rom[28297] = 25'b1111000011110011110100100;
    rom[28298] = 25'b1111000011110000110100001;
    rom[28299] = 25'b1111000011101101110011110;
    rom[28300] = 25'b1111000011101010110011110;
    rom[28301] = 25'b1111000011100111110100000;
    rom[28302] = 25'b1111000011100100110100011;
    rom[28303] = 25'b1111000011100001110101001;
    rom[28304] = 25'b1111000011011110110101111;
    rom[28305] = 25'b1111000011011011110111000;
    rom[28306] = 25'b1111000011011000111000011;
    rom[28307] = 25'b1111000011010101111010000;
    rom[28308] = 25'b1111000011010010111011110;
    rom[28309] = 25'b1111000011001111111101111;
    rom[28310] = 25'b1111000011001101000000001;
    rom[28311] = 25'b1111000011001010000010101;
    rom[28312] = 25'b1111000011000111000101010;
    rom[28313] = 25'b1111000011000100001000010;
    rom[28314] = 25'b1111000011000001001011100;
    rom[28315] = 25'b1111000010111110001110111;
    rom[28316] = 25'b1111000010111011010010100;
    rom[28317] = 25'b1111000010111000010110100;
    rom[28318] = 25'b1111000010110101011010101;
    rom[28319] = 25'b1111000010110010011111000;
    rom[28320] = 25'b1111000010101111100011100;
    rom[28321] = 25'b1111000010101100101000010;
    rom[28322] = 25'b1111000010101001101101011;
    rom[28323] = 25'b1111000010100110110010101;
    rom[28324] = 25'b1111000010100011111000010;
    rom[28325] = 25'b1111000010100000111101111;
    rom[28326] = 25'b1111000010011110000100000;
    rom[28327] = 25'b1111000010011011001010010;
    rom[28328] = 25'b1111000010011000010000110;
    rom[28329] = 25'b1111000010010101010111011;
    rom[28330] = 25'b1111000010010010011110011;
    rom[28331] = 25'b1111000010001111100101100;
    rom[28332] = 25'b1111000010001100101101000;
    rom[28333] = 25'b1111000010001001110100101;
    rom[28334] = 25'b1111000010000110111100101;
    rom[28335] = 25'b1111000010000100000100101;
    rom[28336] = 25'b1111000010000001001101001;
    rom[28337] = 25'b1111000001111110010101101;
    rom[28338] = 25'b1111000001111011011110100;
    rom[28339] = 25'b1111000001111000100111110;
    rom[28340] = 25'b1111000001110101110001000;
    rom[28341] = 25'b1111000001110010111010101;
    rom[28342] = 25'b1111000001110000000100100;
    rom[28343] = 25'b1111000001101101001110100;
    rom[28344] = 25'b1111000001101010011000110;
    rom[28345] = 25'b1111000001100111100011011;
    rom[28346] = 25'b1111000001100100101110001;
    rom[28347] = 25'b1111000001100001111001010;
    rom[28348] = 25'b1111000001011111000100101;
    rom[28349] = 25'b1111000001011100010000000;
    rom[28350] = 25'b1111000001011001011011111;
    rom[28351] = 25'b1111000001010110100111111;
    rom[28352] = 25'b1111000001010011110100010;
    rom[28353] = 25'b1111000001010001000000110;
    rom[28354] = 25'b1111000001001110001101100;
    rom[28355] = 25'b1111000001001011011010100;
    rom[28356] = 25'b1111000001001000100111110;
    rom[28357] = 25'b1111000001000101110101010;
    rom[28358] = 25'b1111000001000011000011000;
    rom[28359] = 25'b1111000001000000010001000;
    rom[28360] = 25'b1111000000111101011111010;
    rom[28361] = 25'b1111000000111010101101110;
    rom[28362] = 25'b1111000000110111111100100;
    rom[28363] = 25'b1111000000110101001011100;
    rom[28364] = 25'b1111000000110010011010110;
    rom[28365] = 25'b1111000000101111101010010;
    rom[28366] = 25'b1111000000101100111010000;
    rom[28367] = 25'b1111000000101010001010000;
    rom[28368] = 25'b1111000000100111011010011;
    rom[28369] = 25'b1111000000100100101010110;
    rom[28370] = 25'b1111000000100001111011101;
    rom[28371] = 25'b1111000000011111001100100;
    rom[28372] = 25'b1111000000011100011101111;
    rom[28373] = 25'b1111000000011001101111011;
    rom[28374] = 25'b1111000000010111000001001;
    rom[28375] = 25'b1111000000010100010011001;
    rom[28376] = 25'b1111000000010001100101100;
    rom[28377] = 25'b1111000000001110111000000;
    rom[28378] = 25'b1111000000001100001010110;
    rom[28379] = 25'b1111000000001001011101111;
    rom[28380] = 25'b1111000000000110110001001;
    rom[28381] = 25'b1111000000000100000100110;
    rom[28382] = 25'b1111000000000001011000101;
    rom[28383] = 25'b1110111111111110101100101;
    rom[28384] = 25'b1110111111111100000001000;
    rom[28385] = 25'b1110111111111001010101100;
    rom[28386] = 25'b1110111111110110101010100;
    rom[28387] = 25'b1110111111110011111111100;
    rom[28388] = 25'b1110111111110001010101000;
    rom[28389] = 25'b1110111111101110101010100;
    rom[28390] = 25'b1110111111101100000000100;
    rom[28391] = 25'b1110111111101001010110101;
    rom[28392] = 25'b1110111111100110101101000;
    rom[28393] = 25'b1110111111100100000011101;
    rom[28394] = 25'b1110111111100001011010101;
    rom[28395] = 25'b1110111111011110110001110;
    rom[28396] = 25'b1110111111011100001001010;
    rom[28397] = 25'b1110111111011001100001000;
    rom[28398] = 25'b1110111111010110111001000;
    rom[28399] = 25'b1110111111010100010001010;
    rom[28400] = 25'b1110111111010001101001110;
    rom[28401] = 25'b1110111111001111000010100;
    rom[28402] = 25'b1110111111001100011011100;
    rom[28403] = 25'b1110111111001001110100111;
    rom[28404] = 25'b1110111111000111001110100;
    rom[28405] = 25'b1110111111000100101000010;
    rom[28406] = 25'b1110111111000010000010011;
    rom[28407] = 25'b1110111110111111011100110;
    rom[28408] = 25'b1110111110111100110111010;
    rom[28409] = 25'b1110111110111010010010010;
    rom[28410] = 25'b1110111110110111101101011;
    rom[28411] = 25'b1110111110110101001000111;
    rom[28412] = 25'b1110111110110010100100100;
    rom[28413] = 25'b1110111110110000000000100;
    rom[28414] = 25'b1110111110101101011100110;
    rom[28415] = 25'b1110111110101010111001010;
    rom[28416] = 25'b1110111110101000010110000;
    rom[28417] = 25'b1110111110100101110011000;
    rom[28418] = 25'b1110111110100011010000011;
    rom[28419] = 25'b1110111110100000101110000;
    rom[28420] = 25'b1110111110011110001011111;
    rom[28421] = 25'b1110111110011011101001111;
    rom[28422] = 25'b1110111110011001001000011;
    rom[28423] = 25'b1110111110010110100111000;
    rom[28424] = 25'b1110111110010100000110000;
    rom[28425] = 25'b1110111110010001100101001;
    rom[28426] = 25'b1110111110001111000100101;
    rom[28427] = 25'b1110111110001100100100011;
    rom[28428] = 25'b1110111110001010000100011;
    rom[28429] = 25'b1110111110000111100100110;
    rom[28430] = 25'b1110111110000101000101010;
    rom[28431] = 25'b1110111110000010100110001;
    rom[28432] = 25'b1110111110000000000111011;
    rom[28433] = 25'b1110111101111101101000110;
    rom[28434] = 25'b1110111101111011001010100;
    rom[28435] = 25'b1110111101111000101100011;
    rom[28436] = 25'b1110111101110110001110101;
    rom[28437] = 25'b1110111101110011110001001;
    rom[28438] = 25'b1110111101110001010011111;
    rom[28439] = 25'b1110111101101110110111000;
    rom[28440] = 25'b1110111101101100011010011;
    rom[28441] = 25'b1110111101101001111110000;
    rom[28442] = 25'b1110111101100111100001111;
    rom[28443] = 25'b1110111101100101000110001;
    rom[28444] = 25'b1110111101100010101010100;
    rom[28445] = 25'b1110111101100000001111010;
    rom[28446] = 25'b1110111101011101110100010;
    rom[28447] = 25'b1110111101011011011001100;
    rom[28448] = 25'b1110111101011000111111001;
    rom[28449] = 25'b1110111101010110100101000;
    rom[28450] = 25'b1110111101010100001011001;
    rom[28451] = 25'b1110111101010001110001100;
    rom[28452] = 25'b1110111101001111011000010;
    rom[28453] = 25'b1110111101001100111111011;
    rom[28454] = 25'b1110111101001010100110100;
    rom[28455] = 25'b1110111101001000001110001;
    rom[28456] = 25'b1110111101000101110101111;
    rom[28457] = 25'b1110111101000011011110000;
    rom[28458] = 25'b1110111101000001000110100;
    rom[28459] = 25'b1110111100111110101111010;
    rom[28460] = 25'b1110111100111100011000010;
    rom[28461] = 25'b1110111100111010000001011;
    rom[28462] = 25'b1110111100110111101010111;
    rom[28463] = 25'b1110111100110101010100110;
    rom[28464] = 25'b1110111100110010111111000;
    rom[28465] = 25'b1110111100110000101001011;
    rom[28466] = 25'b1110111100101110010100000;
    rom[28467] = 25'b1110111100101011111111000;
    rom[28468] = 25'b1110111100101001101010011;
    rom[28469] = 25'b1110111100100111010101111;
    rom[28470] = 25'b1110111100100101000001110;
    rom[28471] = 25'b1110111100100010101101110;
    rom[28472] = 25'b1110111100100000011010010;
    rom[28473] = 25'b1110111100011110000111000;
    rom[28474] = 25'b1110111100011011110100000;
    rom[28475] = 25'b1110111100011001100001010;
    rom[28476] = 25'b1110111100010111001110111;
    rom[28477] = 25'b1110111100010100111100110;
    rom[28478] = 25'b1110111100010010101010111;
    rom[28479] = 25'b1110111100010000011001011;
    rom[28480] = 25'b1110111100001110001000001;
    rom[28481] = 25'b1110111100001011110111001;
    rom[28482] = 25'b1110111100001001100110100;
    rom[28483] = 25'b1110111100000111010110001;
    rom[28484] = 25'b1110111100000101000110001;
    rom[28485] = 25'b1110111100000010110110011;
    rom[28486] = 25'b1110111100000000100110111;
    rom[28487] = 25'b1110111011111110010111101;
    rom[28488] = 25'b1110111011111100001000110;
    rom[28489] = 25'b1110111011111001111010001;
    rom[28490] = 25'b1110111011110111101011111;
    rom[28491] = 25'b1110111011110101011101111;
    rom[28492] = 25'b1110111011110011010000001;
    rom[28493] = 25'b1110111011110001000010110;
    rom[28494] = 25'b1110111011101110110101101;
    rom[28495] = 25'b1110111011101100101000110;
    rom[28496] = 25'b1110111011101010011100010;
    rom[28497] = 25'b1110111011101000010000001;
    rom[28498] = 25'b1110111011100110000100001;
    rom[28499] = 25'b1110111011100011111000100;
    rom[28500] = 25'b1110111011100001101101001;
    rom[28501] = 25'b1110111011011111100010001;
    rom[28502] = 25'b1110111011011101010111011;
    rom[28503] = 25'b1110111011011011001101000;
    rom[28504] = 25'b1110111011011001000010111;
    rom[28505] = 25'b1110111011010110111001000;
    rom[28506] = 25'b1110111011010100101111100;
    rom[28507] = 25'b1110111011010010100110010;
    rom[28508] = 25'b1110111011010000011101011;
    rom[28509] = 25'b1110111011001110010100110;
    rom[28510] = 25'b1110111011001100001100011;
    rom[28511] = 25'b1110111011001010000100100;
    rom[28512] = 25'b1110111011000111111100101;
    rom[28513] = 25'b1110111011000101110101010;
    rom[28514] = 25'b1110111011000011101110010;
    rom[28515] = 25'b1110111011000001100111011;
    rom[28516] = 25'b1110111010111111100000111;
    rom[28517] = 25'b1110111010111101011010110;
    rom[28518] = 25'b1110111010111011010100111;
    rom[28519] = 25'b1110111010111001001111010;
    rom[28520] = 25'b1110111010110111001010000;
    rom[28521] = 25'b1110111010110101000101000;
    rom[28522] = 25'b1110111010110011000000011;
    rom[28523] = 25'b1110111010110000111100000;
    rom[28524] = 25'b1110111010101110111000000;
    rom[28525] = 25'b1110111010101100110100010;
    rom[28526] = 25'b1110111010101010110000111;
    rom[28527] = 25'b1110111010101000101101110;
    rom[28528] = 25'b1110111010100110101010111;
    rom[28529] = 25'b1110111010100100101000011;
    rom[28530] = 25'b1110111010100010100110001;
    rom[28531] = 25'b1110111010100000100100011;
    rom[28532] = 25'b1110111010011110100010110;
    rom[28533] = 25'b1110111010011100100001100;
    rom[28534] = 25'b1110111010011010100000100;
    rom[28535] = 25'b1110111010011000011111111;
    rom[28536] = 25'b1110111010010110011111101;
    rom[28537] = 25'b1110111010010100011111100;
    rom[28538] = 25'b1110111010010010011111111;
    rom[28539] = 25'b1110111010010000100000011;
    rom[28540] = 25'b1110111010001110100001011;
    rom[28541] = 25'b1110111010001100100010101;
    rom[28542] = 25'b1110111010001010100100001;
    rom[28543] = 25'b1110111010001000100110001;
    rom[28544] = 25'b1110111010000110101000010;
    rom[28545] = 25'b1110111010000100101010101;
    rom[28546] = 25'b1110111010000010101101100;
    rom[28547] = 25'b1110111010000000110000101;
    rom[28548] = 25'b1110111001111110110100001;
    rom[28549] = 25'b1110111001111100110111111;
    rom[28550] = 25'b1110111001111010111100000;
    rom[28551] = 25'b1110111001111001000000011;
    rom[28552] = 25'b1110111001110111000101000;
    rom[28553] = 25'b1110111001110101001010001;
    rom[28554] = 25'b1110111001110011001111011;
    rom[28555] = 25'b1110111001110001010101000;
    rom[28556] = 25'b1110111001101111011011000;
    rom[28557] = 25'b1110111001101101100001011;
    rom[28558] = 25'b1110111001101011101000000;
    rom[28559] = 25'b1110111001101001101111000;
    rom[28560] = 25'b1110111001100111110110010;
    rom[28561] = 25'b1110111001100101111101110;
    rom[28562] = 25'b1110111001100100000101101;
    rom[28563] = 25'b1110111001100010001101111;
    rom[28564] = 25'b1110111001100000010110011;
    rom[28565] = 25'b1110111001011110011111010;
    rom[28566] = 25'b1110111001011100101000011;
    rom[28567] = 25'b1110111001011010110001111;
    rom[28568] = 25'b1110111001011000111011110;
    rom[28569] = 25'b1110111001010111000101111;
    rom[28570] = 25'b1110111001010101010000100;
    rom[28571] = 25'b1110111001010011011011010;
    rom[28572] = 25'b1110111001010001100110011;
    rom[28573] = 25'b1110111001001111110001110;
    rom[28574] = 25'b1110111001001101111101100;
    rom[28575] = 25'b1110111001001100001001101;
    rom[28576] = 25'b1110111001001010010110001;
    rom[28577] = 25'b1110111001001000100010111;
    rom[28578] = 25'b1110111001000110101111111;
    rom[28579] = 25'b1110111001000100111101010;
    rom[28580] = 25'b1110111001000011001011000;
    rom[28581] = 25'b1110111001000001011001001;
    rom[28582] = 25'b1110111000111111100111011;
    rom[28583] = 25'b1110111000111101110110001;
    rom[28584] = 25'b1110111000111100000101001;
    rom[28585] = 25'b1110111000111010010100100;
    rom[28586] = 25'b1110111000111000100100010;
    rom[28587] = 25'b1110111000110110110100010;
    rom[28588] = 25'b1110111000110101000100101;
    rom[28589] = 25'b1110111000110011010101010;
    rom[28590] = 25'b1110111000110001100110011;
    rom[28591] = 25'b1110111000101111110111101;
    rom[28592] = 25'b1110111000101110001001010;
    rom[28593] = 25'b1110111000101100011011010;
    rom[28594] = 25'b1110111000101010101101101;
    rom[28595] = 25'b1110111000101001000000010;
    rom[28596] = 25'b1110111000100111010011011;
    rom[28597] = 25'b1110111000100101100110101;
    rom[28598] = 25'b1110111000100011111010010;
    rom[28599] = 25'b1110111000100010001110011;
    rom[28600] = 25'b1110111000100000100010101;
    rom[28601] = 25'b1110111000011110110111010;
    rom[28602] = 25'b1110111000011101001100011;
    rom[28603] = 25'b1110111000011011100001101;
    rom[28604] = 25'b1110111000011001110111011;
    rom[28605] = 25'b1110111000011000001101011;
    rom[28606] = 25'b1110111000010110100011101;
    rom[28607] = 25'b1110111000010100111010010;
    rom[28608] = 25'b1110111000010011010001010;
    rom[28609] = 25'b1110111000010001101000101;
    rom[28610] = 25'b1110111000010000000000010;
    rom[28611] = 25'b1110111000001110011000011;
    rom[28612] = 25'b1110111000001100110000110;
    rom[28613] = 25'b1110111000001011001001011;
    rom[28614] = 25'b1110111000001001100010011;
    rom[28615] = 25'b1110111000000111111011110;
    rom[28616] = 25'b1110111000000110010101100;
    rom[28617] = 25'b1110111000000100101111100;
    rom[28618] = 25'b1110111000000011001001111;
    rom[28619] = 25'b1110111000000001100100101;
    rom[28620] = 25'b1110110111111111111111110;
    rom[28621] = 25'b1110110111111110011011001;
    rom[28622] = 25'b1110110111111100110110111;
    rom[28623] = 25'b1110110111111011010011000;
    rom[28624] = 25'b1110110111111001101111011;
    rom[28625] = 25'b1110110111111000001100001;
    rom[28626] = 25'b1110110111110110101001010;
    rom[28627] = 25'b1110110111110101000110110;
    rom[28628] = 25'b1110110111110011100100100;
    rom[28629] = 25'b1110110111110010000010101;
    rom[28630] = 25'b1110110111110000100001001;
    rom[28631] = 25'b1110110111101111000000000;
    rom[28632] = 25'b1110110111101101011111001;
    rom[28633] = 25'b1110110111101011111110101;
    rom[28634] = 25'b1110110111101010011110100;
    rom[28635] = 25'b1110110111101000111110101;
    rom[28636] = 25'b1110110111100111011111010;
    rom[28637] = 25'b1110110111100110000000001;
    rom[28638] = 25'b1110110111100100100001011;
    rom[28639] = 25'b1110110111100011000011000;
    rom[28640] = 25'b1110110111100001100100111;
    rom[28641] = 25'b1110110111100000000111001;
    rom[28642] = 25'b1110110111011110101001110;
    rom[28643] = 25'b1110110111011101001100110;
    rom[28644] = 25'b1110110111011011110000001;
    rom[28645] = 25'b1110110111011010010011110;
    rom[28646] = 25'b1110110111011000110111110;
    rom[28647] = 25'b1110110111010111011100001;
    rom[28648] = 25'b1110110111010110000000111;
    rom[28649] = 25'b1110110111010100100101111;
    rom[28650] = 25'b1110110111010011001011010;
    rom[28651] = 25'b1110110111010001110001000;
    rom[28652] = 25'b1110110111010000010111001;
    rom[28653] = 25'b1110110111001110111101101;
    rom[28654] = 25'b1110110111001101100100100;
    rom[28655] = 25'b1110110111001100001011101;
    rom[28656] = 25'b1110110111001010110011001;
    rom[28657] = 25'b1110110111001001011011000;
    rom[28658] = 25'b1110110111001000000011010;
    rom[28659] = 25'b1110110111000110101011110;
    rom[28660] = 25'b1110110111000101010100110;
    rom[28661] = 25'b1110110111000011111110000;
    rom[28662] = 25'b1110110111000010100111101;
    rom[28663] = 25'b1110110111000001010001101;
    rom[28664] = 25'b1110110110111111111100000;
    rom[28665] = 25'b1110110110111110100110101;
    rom[28666] = 25'b1110110110111101010001110;
    rom[28667] = 25'b1110110110111011111101001;
    rom[28668] = 25'b1110110110111010101000111;
    rom[28669] = 25'b1110110110111001010100111;
    rom[28670] = 25'b1110110110111000000001011;
    rom[28671] = 25'b1110110110110110101110010;
    rom[28672] = 25'b1110110110110101011011100;
    rom[28673] = 25'b1110110110110100001001000;
    rom[28674] = 25'b1110110110110010110110111;
    rom[28675] = 25'b1110110110110001100101001;
    rom[28676] = 25'b1110110110110000010011110;
    rom[28677] = 25'b1110110110101111000010110;
    rom[28678] = 25'b1110110110101101110010000;
    rom[28679] = 25'b1110110110101100100001110;
    rom[28680] = 25'b1110110110101011010001110;
    rom[28681] = 25'b1110110110101010000010010;
    rom[28682] = 25'b1110110110101000110011000;
    rom[28683] = 25'b1110110110100111100100001;
    rom[28684] = 25'b1110110110100110010101101;
    rom[28685] = 25'b1110110110100101000111011;
    rom[28686] = 25'b1110110110100011111001101;
    rom[28687] = 25'b1110110110100010101100010;
    rom[28688] = 25'b1110110110100001011111001;
    rom[28689] = 25'b1110110110100000010010011;
    rom[28690] = 25'b1110110110011111000110001;
    rom[28691] = 25'b1110110110011101111010001;
    rom[28692] = 25'b1110110110011100101110100;
    rom[28693] = 25'b1110110110011011100011010;
    rom[28694] = 25'b1110110110011010011000011;
    rom[28695] = 25'b1110110110011001001101111;
    rom[28696] = 25'b1110110110011000000011110;
    rom[28697] = 25'b1110110110010110111001111;
    rom[28698] = 25'b1110110110010101110000011;
    rom[28699] = 25'b1110110110010100100111011;
    rom[28700] = 25'b1110110110010011011110101;
    rom[28701] = 25'b1110110110010010010110010;
    rom[28702] = 25'b1110110110010001001110011;
    rom[28703] = 25'b1110110110010000000110110;
    rom[28704] = 25'b1110110110001110111111100;
    rom[28705] = 25'b1110110110001101111000101;
    rom[28706] = 25'b1110110110001100110010001;
    rom[28707] = 25'b1110110110001011101100000;
    rom[28708] = 25'b1110110110001010100110010;
    rom[28709] = 25'b1110110110001001100000111;
    rom[28710] = 25'b1110110110001000011011110;
    rom[28711] = 25'b1110110110000111010111001;
    rom[28712] = 25'b1110110110000110010010110;
    rom[28713] = 25'b1110110110000101001110111;
    rom[28714] = 25'b1110110110000100001011010;
    rom[28715] = 25'b1110110110000011001000001;
    rom[28716] = 25'b1110110110000010000101010;
    rom[28717] = 25'b1110110110000001000010111;
    rom[28718] = 25'b1110110110000000000000110;
    rom[28719] = 25'b1110110101111110111111001;
    rom[28720] = 25'b1110110101111101111101110;
    rom[28721] = 25'b1110110101111100111100111;
    rom[28722] = 25'b1110110101111011111100010;
    rom[28723] = 25'b1110110101111010111100000;
    rom[28724] = 25'b1110110101111001111100010;
    rom[28725] = 25'b1110110101111000111100101;
    rom[28726] = 25'b1110110101110111111101100;
    rom[28727] = 25'b1110110101110110111110111;
    rom[28728] = 25'b1110110101110110000000100;
    rom[28729] = 25'b1110110101110101000010100;
    rom[28730] = 25'b1110110101110100000101000;
    rom[28731] = 25'b1110110101110011000111110;
    rom[28732] = 25'b1110110101110010001010111;
    rom[28733] = 25'b1110110101110001001110011;
    rom[28734] = 25'b1110110101110000010010010;
    rom[28735] = 25'b1110110101101111010110101;
    rom[28736] = 25'b1110110101101110011011001;
    rom[28737] = 25'b1110110101101101100000010;
    rom[28738] = 25'b1110110101101100100101110;
    rom[28739] = 25'b1110110101101011101011011;
    rom[28740] = 25'b1110110101101010110001101;
    rom[28741] = 25'b1110110101101001111000001;
    rom[28742] = 25'b1110110101101000111111000;
    rom[28743] = 25'b1110110101101000000110011;
    rom[28744] = 25'b1110110101100111001110000;
    rom[28745] = 25'b1110110101100110010110001;
    rom[28746] = 25'b1110110101100101011110100;
    rom[28747] = 25'b1110110101100100100111011;
    rom[28748] = 25'b1110110101100011110000100;
    rom[28749] = 25'b1110110101100010111010001;
    rom[28750] = 25'b1110110101100010000100000;
    rom[28751] = 25'b1110110101100001001110011;
    rom[28752] = 25'b1110110101100000011001001;
    rom[28753] = 25'b1110110101011111100100010;
    rom[28754] = 25'b1110110101011110101111101;
    rom[28755] = 25'b1110110101011101111011100;
    rom[28756] = 25'b1110110101011101000111110;
    rom[28757] = 25'b1110110101011100010100011;
    rom[28758] = 25'b1110110101011011100001100;
    rom[28759] = 25'b1110110101011010101110111;
    rom[28760] = 25'b1110110101011001111100101;
    rom[28761] = 25'b1110110101011001001010110;
    rom[28762] = 25'b1110110101011000011001010;
    rom[28763] = 25'b1110110101010111101000010;
    rom[28764] = 25'b1110110101010110110111100;
    rom[28765] = 25'b1110110101010110000111001;
    rom[28766] = 25'b1110110101010101010111010;
    rom[28767] = 25'b1110110101010100100111110;
    rom[28768] = 25'b1110110101010011111000100;
    rom[28769] = 25'b1110110101010011001001111;
    rom[28770] = 25'b1110110101010010011011100;
    rom[28771] = 25'b1110110101010001101101100;
    rom[28772] = 25'b1110110101010000111111111;
    rom[28773] = 25'b1110110101010000010010101;
    rom[28774] = 25'b1110110101001111100101111;
    rom[28775] = 25'b1110110101001110111001011;
    rom[28776] = 25'b1110110101001110001101011;
    rom[28777] = 25'b1110110101001101100001101;
    rom[28778] = 25'b1110110101001100110110011;
    rom[28779] = 25'b1110110101001100001011100;
    rom[28780] = 25'b1110110101001011100001000;
    rom[28781] = 25'b1110110101001010110110111;
    rom[28782] = 25'b1110110101001010001101010;
    rom[28783] = 25'b1110110101001001100011111;
    rom[28784] = 25'b1110110101001000111011000;
    rom[28785] = 25'b1110110101001000010010011;
    rom[28786] = 25'b1110110101000111101010010;
    rom[28787] = 25'b1110110101000111000010100;
    rom[28788] = 25'b1110110101000110011011001;
    rom[28789] = 25'b1110110101000101110100001;
    rom[28790] = 25'b1110110101000101001101100;
    rom[28791] = 25'b1110110101000100100111011;
    rom[28792] = 25'b1110110101000100000001100;
    rom[28793] = 25'b1110110101000011011100001;
    rom[28794] = 25'b1110110101000010110111001;
    rom[28795] = 25'b1110110101000010010010100;
    rom[28796] = 25'b1110110101000001101110010;
    rom[28797] = 25'b1110110101000001001010011;
    rom[28798] = 25'b1110110101000000100111000;
    rom[28799] = 25'b1110110101000000000011111;
    rom[28800] = 25'b1110110100111111100001010;
    rom[28801] = 25'b1110110100111110111111001;
    rom[28802] = 25'b1110110100111110011101001;
    rom[28803] = 25'b1110110100111101111011110;
    rom[28804] = 25'b1110110100111101011010101;
    rom[28805] = 25'b1110110100111100111010000;
    rom[28806] = 25'b1110110100111100011001101;
    rom[28807] = 25'b1110110100111011111001111;
    rom[28808] = 25'b1110110100111011011010011;
    rom[28809] = 25'b1110110100111010111011010;
    rom[28810] = 25'b1110110100111010011100100;
    rom[28811] = 25'b1110110100111001111110010;
    rom[28812] = 25'b1110110100111001100000011;
    rom[28813] = 25'b1110110100111001000010111;
    rom[28814] = 25'b1110110100111000100101111;
    rom[28815] = 25'b1110110100111000001001001;
    rom[28816] = 25'b1110110100110111101100110;
    rom[28817] = 25'b1110110100110111010001000;
    rom[28818] = 25'b1110110100110110110101011;
    rom[28819] = 25'b1110110100110110011010011;
    rom[28820] = 25'b1110110100110101111111101;
    rom[28821] = 25'b1110110100110101100101011;
    rom[28822] = 25'b1110110100110101001011100;
    rom[28823] = 25'b1110110100110100110010000;
    rom[28824] = 25'b1110110100110100011000111;
    rom[28825] = 25'b1110110100110100000000010;
    rom[28826] = 25'b1110110100110011101000000;
    rom[28827] = 25'b1110110100110011010000000;
    rom[28828] = 25'b1110110100110010111000101;
    rom[28829] = 25'b1110110100110010100001100;
    rom[28830] = 25'b1110110100110010001010111;
    rom[28831] = 25'b1110110100110001110100100;
    rom[28832] = 25'b1110110100110001011110101;
    rom[28833] = 25'b1110110100110001001001010;
    rom[28834] = 25'b1110110100110000110100010;
    rom[28835] = 25'b1110110100110000011111100;
    rom[28836] = 25'b1110110100110000001011010;
    rom[28837] = 25'b1110110100101111110111100;
    rom[28838] = 25'b1110110100101111100100000;
    rom[28839] = 25'b1110110100101111010001000;
    rom[28840] = 25'b1110110100101110111110011;
    rom[28841] = 25'b1110110100101110101100001;
    rom[28842] = 25'b1110110100101110011010010;
    rom[28843] = 25'b1110110100101110001000111;
    rom[28844] = 25'b1110110100101101110111111;
    rom[28845] = 25'b1110110100101101100111010;
    rom[28846] = 25'b1110110100101101010111001;
    rom[28847] = 25'b1110110100101101000111011;
    rom[28848] = 25'b1110110100101100111000000;
    rom[28849] = 25'b1110110100101100101001001;
    rom[28850] = 25'b1110110100101100011010100;
    rom[28851] = 25'b1110110100101100001100011;
    rom[28852] = 25'b1110110100101011111110101;
    rom[28853] = 25'b1110110100101011110001011;
    rom[28854] = 25'b1110110100101011100100100;
    rom[28855] = 25'b1110110100101011011000000;
    rom[28856] = 25'b1110110100101011001011110;
    rom[28857] = 25'b1110110100101011000000001;
    rom[28858] = 25'b1110110100101010110100111;
    rom[28859] = 25'b1110110100101010101010000;
    rom[28860] = 25'b1110110100101010011111100;
    rom[28861] = 25'b1110110100101010010101100;
    rom[28862] = 25'b1110110100101010001011111;
    rom[28863] = 25'b1110110100101010000010110;
    rom[28864] = 25'b1110110100101001111001111;
    rom[28865] = 25'b1110110100101001110001100;
    rom[28866] = 25'b1110110100101001101001101;
    rom[28867] = 25'b1110110100101001100010000;
    rom[28868] = 25'b1110110100101001011010111;
    rom[28869] = 25'b1110110100101001010100001;
    rom[28870] = 25'b1110110100101001001101111;
    rom[28871] = 25'b1110110100101001001000000;
    rom[28872] = 25'b1110110100101001000010100;
    rom[28873] = 25'b1110110100101000111101010;
    rom[28874] = 25'b1110110100101000111000110;
    rom[28875] = 25'b1110110100101000110100011;
    rom[28876] = 25'b1110110100101000110000101;
    rom[28877] = 25'b1110110100101000101101010;
    rom[28878] = 25'b1110110100101000101010010;
    rom[28879] = 25'b1110110100101000100111101;
    rom[28880] = 25'b1110110100101000100101100;
    rom[28881] = 25'b1110110100101000100011110;
    rom[28882] = 25'b1110110100101000100010011;
    rom[28883] = 25'b1110110100101000100001100;
    rom[28884] = 25'b1110110100101000100001000;
    rom[28885] = 25'b1110110100101000100000111;
    rom[28886] = 25'b1110110100101000100001010;
    rom[28887] = 25'b1110110100101000100010000;
    rom[28888] = 25'b1110110100101000100011001;
    rom[28889] = 25'b1110110100101000100100111;
    rom[28890] = 25'b1110110100101000100110110;
    rom[28891] = 25'b1110110100101000101001010;
    rom[28892] = 25'b1110110100101000101100001;
    rom[28893] = 25'b1110110100101000101111011;
    rom[28894] = 25'b1110110100101000110011001;
    rom[28895] = 25'b1110110100101000110111010;
    rom[28896] = 25'b1110110100101000111011110;
    rom[28897] = 25'b1110110100101001000000101;
    rom[28898] = 25'b1110110100101001000110001;
    rom[28899] = 25'b1110110100101001001011111;
    rom[28900] = 25'b1110110100101001010010001;
    rom[28901] = 25'b1110110100101001011000110;
    rom[28902] = 25'b1110110100101001011111111;
    rom[28903] = 25'b1110110100101001100111011;
    rom[28904] = 25'b1110110100101001101111001;
    rom[28905] = 25'b1110110100101001110111101;
    rom[28906] = 25'b1110110100101010000000011;
    rom[28907] = 25'b1110110100101010001001100;
    rom[28908] = 25'b1110110100101010010011001;
    rom[28909] = 25'b1110110100101010011101001;
    rom[28910] = 25'b1110110100101010100111101;
    rom[28911] = 25'b1110110100101010110010100;
    rom[28912] = 25'b1110110100101010111101110;
    rom[28913] = 25'b1110110100101011001001100;
    rom[28914] = 25'b1110110100101011010101101;
    rom[28915] = 25'b1110110100101011100010010;
    rom[28916] = 25'b1110110100101011101111010;
    rom[28917] = 25'b1110110100101011111100101;
    rom[28918] = 25'b1110110100101100001010101;
    rom[28919] = 25'b1110110100101100011000110;
    rom[28920] = 25'b1110110100101100100111100;
    rom[28921] = 25'b1110110100101100110110101;
    rom[28922] = 25'b1110110100101101000110010;
    rom[28923] = 25'b1110110100101101010110010;
    rom[28924] = 25'b1110110100101101100110101;
    rom[28925] = 25'b1110110100101101110111100;
    rom[28926] = 25'b1110110100101110001000110;
    rom[28927] = 25'b1110110100101110011010100;
    rom[28928] = 25'b1110110100101110101100101;
    rom[28929] = 25'b1110110100101110111111001;
    rom[28930] = 25'b1110110100101111010010001;
    rom[28931] = 25'b1110110100101111100101100;
    rom[28932] = 25'b1110110100101111111001100;
    rom[28933] = 25'b1110110100110000001101110;
    rom[28934] = 25'b1110110100110000100010100;
    rom[28935] = 25'b1110110100110000110111100;
    rom[28936] = 25'b1110110100110001001101001;
    rom[28937] = 25'b1110110100110001100011001;
    rom[28938] = 25'b1110110100110001111001101;
    rom[28939] = 25'b1110110100110010010000100;
    rom[28940] = 25'b1110110100110010100111110;
    rom[28941] = 25'b1110110100110010111111011;
    rom[28942] = 25'b1110110100110011010111101;
    rom[28943] = 25'b1110110100110011110000001;
    rom[28944] = 25'b1110110100110100001001010;
    rom[28945] = 25'b1110110100110100100010110;
    rom[28946] = 25'b1110110100110100111100101;
    rom[28947] = 25'b1110110100110101010110111;
    rom[28948] = 25'b1110110100110101110001101;
    rom[28949] = 25'b1110110100110110001100110;
    rom[28950] = 25'b1110110100110110101000011;
    rom[28951] = 25'b1110110100110111000100100;
    rom[28952] = 25'b1110110100110111100001000;
    rom[28953] = 25'b1110110100110111111110000;
    rom[28954] = 25'b1110110100111000011011010;
    rom[28955] = 25'b1110110100111000111001001;
    rom[28956] = 25'b1110110100111001010111011;
    rom[28957] = 25'b1110110100111001110110000;
    rom[28958] = 25'b1110110100111010010101001;
    rom[28959] = 25'b1110110100111010110100101;
    rom[28960] = 25'b1110110100111011010100101;
    rom[28961] = 25'b1110110100111011110101000;
    rom[28962] = 25'b1110110100111100010101111;
    rom[28963] = 25'b1110110100111100110111010;
    rom[28964] = 25'b1110110100111101011000111;
    rom[28965] = 25'b1110110100111101111011001;
    rom[28966] = 25'b1110110100111110011101101;
    rom[28967] = 25'b1110110100111111000000101;
    rom[28968] = 25'b1110110100111111100100001;
    rom[28969] = 25'b1110110101000000001000001;
    rom[28970] = 25'b1110110101000000101100011;
    rom[28971] = 25'b1110110101000001010001010;
    rom[28972] = 25'b1110110101000001110110011;
    rom[28973] = 25'b1110110101000010011100001;
    rom[28974] = 25'b1110110101000011000010010;
    rom[28975] = 25'b1110110101000011101000110;
    rom[28976] = 25'b1110110101000100001111110;
    rom[28977] = 25'b1110110101000100110111001;
    rom[28978] = 25'b1110110101000101011111000;
    rom[28979] = 25'b1110110101000110000111011;
    rom[28980] = 25'b1110110101000110110000001;
    rom[28981] = 25'b1110110101000111011001010;
    rom[28982] = 25'b1110110101001000000010111;
    rom[28983] = 25'b1110110101001000101101000;
    rom[28984] = 25'b1110110101001001010111100;
    rom[28985] = 25'b1110110101001010000010100;
    rom[28986] = 25'b1110110101001010101101111;
    rom[28987] = 25'b1110110101001011011001110;
    rom[28988] = 25'b1110110101001100000110000;
    rom[28989] = 25'b1110110101001100110010110;
    rom[28990] = 25'b1110110101001101011111111;
    rom[28991] = 25'b1110110101001110001101100;
    rom[28992] = 25'b1110110101001110111011100;
    rom[28993] = 25'b1110110101001111101010000;
    rom[28994] = 25'b1110110101010000011001000;
    rom[28995] = 25'b1110110101010001001000011;
    rom[28996] = 25'b1110110101010001111000010;
    rom[28997] = 25'b1110110101010010101000100;
    rom[28998] = 25'b1110110101010011011001001;
    rom[28999] = 25'b1110110101010100001010011;
    rom[29000] = 25'b1110110101010100111100000;
    rom[29001] = 25'b1110110101010101101110000;
    rom[29002] = 25'b1110110101010110100000101;
    rom[29003] = 25'b1110110101010111010011100;
    rom[29004] = 25'b1110110101011000000110111;
    rom[29005] = 25'b1110110101011000111010110;
    rom[29006] = 25'b1110110101011001101111000;
    rom[29007] = 25'b1110110101011010100011110;
    rom[29008] = 25'b1110110101011011011001000;
    rom[29009] = 25'b1110110101011100001110100;
    rom[29010] = 25'b1110110101011101000100101;
    rom[29011] = 25'b1110110101011101111011001;
    rom[29012] = 25'b1110110101011110110010001;
    rom[29013] = 25'b1110110101011111101001100;
    rom[29014] = 25'b1110110101100000100001100;
    rom[29015] = 25'b1110110101100001011001110;
    rom[29016] = 25'b1110110101100010010010101;
    rom[29017] = 25'b1110110101100011001011110;
    rom[29018] = 25'b1110110101100100000101100;
    rom[29019] = 25'b1110110101100100111111100;
    rom[29020] = 25'b1110110101100101111010001;
    rom[29021] = 25'b1110110101100110110101001;
    rom[29022] = 25'b1110110101100111110000101;
    rom[29023] = 25'b1110110101101000101100100;
    rom[29024] = 25'b1110110101101001101000111;
    rom[29025] = 25'b1110110101101010100101101;
    rom[29026] = 25'b1110110101101011100010111;
    rom[29027] = 25'b1110110101101100100000101;
    rom[29028] = 25'b1110110101101101011110110;
    rom[29029] = 25'b1110110101101110011101011;
    rom[29030] = 25'b1110110101101111011100100;
    rom[29031] = 25'b1110110101110000011100000;
    rom[29032] = 25'b1110110101110001011011111;
    rom[29033] = 25'b1110110101110010011100011;
    rom[29034] = 25'b1110110101110011011101010;
    rom[29035] = 25'b1110110101110100011110101;
    rom[29036] = 25'b1110110101110101100000011;
    rom[29037] = 25'b1110110101110110100010101;
    rom[29038] = 25'b1110110101110111100101010;
    rom[29039] = 25'b1110110101111000101000011;
    rom[29040] = 25'b1110110101111001101100000;
    rom[29041] = 25'b1110110101111010110000001;
    rom[29042] = 25'b1110110101111011110100101;
    rom[29043] = 25'b1110110101111100111001101;
    rom[29044] = 25'b1110110101111101111111000;
    rom[29045] = 25'b1110110101111111000100111;
    rom[29046] = 25'b1110110110000000001011001;
    rom[29047] = 25'b1110110110000001010001111;
    rom[29048] = 25'b1110110110000010011001001;
    rom[29049] = 25'b1110110110000011100000111;
    rom[29050] = 25'b1110110110000100101001000;
    rom[29051] = 25'b1110110110000101110001101;
    rom[29052] = 25'b1110110110000110111010101;
    rom[29053] = 25'b1110110110001000000100001;
    rom[29054] = 25'b1110110110001001001110001;
    rom[29055] = 25'b1110110110001010011000101;
    rom[29056] = 25'b1110110110001011100011100;
    rom[29057] = 25'b1110110110001100101110111;
    rom[29058] = 25'b1110110110001101111010101;
    rom[29059] = 25'b1110110110001111000110111;
    rom[29060] = 25'b1110110110010000010011100;
    rom[29061] = 25'b1110110110010001100000110;
    rom[29062] = 25'b1110110110010010101110011;
    rom[29063] = 25'b1110110110010011111100100;
    rom[29064] = 25'b1110110110010101001011000;
    rom[29065] = 25'b1110110110010110011010000;
    rom[29066] = 25'b1110110110010111101001100;
    rom[29067] = 25'b1110110110011000111001011;
    rom[29068] = 25'b1110110110011010001001110;
    rom[29069] = 25'b1110110110011011011010101;
    rom[29070] = 25'b1110110110011100101011111;
    rom[29071] = 25'b1110110110011101111101101;
    rom[29072] = 25'b1110110110011111001111111;
    rom[29073] = 25'b1110110110100000100010100;
    rom[29074] = 25'b1110110110100001110101101;
    rom[29075] = 25'b1110110110100011001001010;
    rom[29076] = 25'b1110110110100100011101010;
    rom[29077] = 25'b1110110110100101110001111;
    rom[29078] = 25'b1110110110100111000110111;
    rom[29079] = 25'b1110110110101000011100010;
    rom[29080] = 25'b1110110110101001110010001;
    rom[29081] = 25'b1110110110101011001000100;
    rom[29082] = 25'b1110110110101100011111011;
    rom[29083] = 25'b1110110110101101110110110;
    rom[29084] = 25'b1110110110101111001110011;
    rom[29085] = 25'b1110110110110000100110101;
    rom[29086] = 25'b1110110110110001111111011;
    rom[29087] = 25'b1110110110110011011000100;
    rom[29088] = 25'b1110110110110100110010001;
    rom[29089] = 25'b1110110110110110001100001;
    rom[29090] = 25'b1110110110110111100110101;
    rom[29091] = 25'b1110110110111001000001101;
    rom[29092] = 25'b1110110110111010011101001;
    rom[29093] = 25'b1110110110111011111001000;
    rom[29094] = 25'b1110110110111101010101100;
    rom[29095] = 25'b1110110110111110110010010;
    rom[29096] = 25'b1110110111000000001111101;
    rom[29097] = 25'b1110110111000001101101011;
    rom[29098] = 25'b1110110111000011001011101;
    rom[29099] = 25'b1110110111000100101010011;
    rom[29100] = 25'b1110110111000110001001100;
    rom[29101] = 25'b1110110111000111101001001;
    rom[29102] = 25'b1110110111001001001001010;
    rom[29103] = 25'b1110110111001010101001110;
    rom[29104] = 25'b1110110111001100001010111;
    rom[29105] = 25'b1110110111001101101100011;
    rom[29106] = 25'b1110110111001111001110010;
    rom[29107] = 25'b1110110111010000110000110;
    rom[29108] = 25'b1110110111010010010011101;
    rom[29109] = 25'b1110110111010011110111000;
    rom[29110] = 25'b1110110111010101011010111;
    rom[29111] = 25'b1110110111010110111111010;
    rom[29112] = 25'b1110110111011000100100000;
    rom[29113] = 25'b1110110111011010001001010;
    rom[29114] = 25'b1110110111011011101110111;
    rom[29115] = 25'b1110110111011101010101000;
    rom[29116] = 25'b1110110111011110111011110;
    rom[29117] = 25'b1110110111100000100010110;
    rom[29118] = 25'b1110110111100010001010011;
    rom[29119] = 25'b1110110111100011110010011;
    rom[29120] = 25'b1110110111100101011010111;
    rom[29121] = 25'b1110110111100111000100000;
    rom[29122] = 25'b1110110111101000101101011;
    rom[29123] = 25'b1110110111101010010111010;
    rom[29124] = 25'b1110110111101100000001101;
    rom[29125] = 25'b1110110111101101101100101;
    rom[29126] = 25'b1110110111101111010111111;
    rom[29127] = 25'b1110110111110001000011101;
    rom[29128] = 25'b1110110111110010110000000;
    rom[29129] = 25'b1110110111110100011100101;
    rom[29130] = 25'b1110110111110110001001111;
    rom[29131] = 25'b1110110111110111110111101;
    rom[29132] = 25'b1110110111111001100101101;
    rom[29133] = 25'b1110110111111011010100011;
    rom[29134] = 25'b1110110111111101000011100;
    rom[29135] = 25'b1110110111111110110011000;
    rom[29136] = 25'b1110111000000000100011000;
    rom[29137] = 25'b1110111000000010010011101;
    rom[29138] = 25'b1110111000000100000100100;
    rom[29139] = 25'b1110111000000101110110000;
    rom[29140] = 25'b1110111000000111100111111;
    rom[29141] = 25'b1110111000001001011010010;
    rom[29142] = 25'b1110111000001011001101001;
    rom[29143] = 25'b1110111000001101000000100;
    rom[29144] = 25'b1110111000001110110100010;
    rom[29145] = 25'b1110111000010000101000101;
    rom[29146] = 25'b1110111000010010011101011;
    rom[29147] = 25'b1110111000010100010010101;
    rom[29148] = 25'b1110111000010110001000011;
    rom[29149] = 25'b1110111000010111111110100;
    rom[29150] = 25'b1110111000011001110101001;
    rom[29151] = 25'b1110111000011011101100010;
    rom[29152] = 25'b1110111000011101100011111;
    rom[29153] = 25'b1110111000011111011100000;
    rom[29154] = 25'b1110111000100001010100100;
    rom[29155] = 25'b1110111000100011001101100;
    rom[29156] = 25'b1110111000100101000111000;
    rom[29157] = 25'b1110111000100111000001000;
    rom[29158] = 25'b1110111000101000111011100;
    rom[29159] = 25'b1110111000101010110110011;
    rom[29160] = 25'b1110111000101100110001110;
    rom[29161] = 25'b1110111000101110101101101;
    rom[29162] = 25'b1110111000110000101001111;
    rom[29163] = 25'b1110111000110010100110110;
    rom[29164] = 25'b1110111000110100100100001;
    rom[29165] = 25'b1110111000110110100001111;
    rom[29166] = 25'b1110111000111000100000001;
    rom[29167] = 25'b1110111000111010011110111;
    rom[29168] = 25'b1110111000111100011110001;
    rom[29169] = 25'b1110111000111110011101110;
    rom[29170] = 25'b1110111001000000011101111;
    rom[29171] = 25'b1110111001000010011110100;
    rom[29172] = 25'b1110111001000100011111101;
    rom[29173] = 25'b1110111001000110100001010;
    rom[29174] = 25'b1110111001001000100011011;
    rom[29175] = 25'b1110111001001010100101111;
    rom[29176] = 25'b1110111001001100101000111;
    rom[29177] = 25'b1110111001001110101100011;
    rom[29178] = 25'b1110111001010000110000011;
    rom[29179] = 25'b1110111001010010110100110;
    rom[29180] = 25'b1110111001010100111001110;
    rom[29181] = 25'b1110111001010110111111010;
    rom[29182] = 25'b1110111001011001000101000;
    rom[29183] = 25'b1110111001011011001011011;
    rom[29184] = 25'b1110111001011101010010010;
    rom[29185] = 25'b1110111001011111011001101;
    rom[29186] = 25'b1110111001100001100001100;
    rom[29187] = 25'b1110111001100011101001110;
    rom[29188] = 25'b1110111001100101110010011;
    rom[29189] = 25'b1110111001100111111011110;
    rom[29190] = 25'b1110111001101010000101100;
    rom[29191] = 25'b1110111001101100001111101;
    rom[29192] = 25'b1110111001101110011010011;
    rom[29193] = 25'b1110111001110000100101100;
    rom[29194] = 25'b1110111001110010110001001;
    rom[29195] = 25'b1110111001110100111101010;
    rom[29196] = 25'b1110111001110111001001111;
    rom[29197] = 25'b1110111001111001010110111;
    rom[29198] = 25'b1110111001111011100100100;
    rom[29199] = 25'b1110111001111101110010100;
    rom[29200] = 25'b1110111010000000000001001;
    rom[29201] = 25'b1110111010000010010000001;
    rom[29202] = 25'b1110111010000100011111101;
    rom[29203] = 25'b1110111010000110101111101;
    rom[29204] = 25'b1110111010001001000000000;
    rom[29205] = 25'b1110111010001011010001000;
    rom[29206] = 25'b1110111010001101100010011;
    rom[29207] = 25'b1110111010001111110100011;
    rom[29208] = 25'b1110111010010010000110101;
    rom[29209] = 25'b1110111010010100011001101;
    rom[29210] = 25'b1110111010010110101101000;
    rom[29211] = 25'b1110111010011001000000110;
    rom[29212] = 25'b1110111010011011010101001;
    rom[29213] = 25'b1110111010011101101001111;
    rom[29214] = 25'b1110111010011111111111001;
    rom[29215] = 25'b1110111010100010010101000;
    rom[29216] = 25'b1110111010100100101011001;
    rom[29217] = 25'b1110111010100111000001111;
    rom[29218] = 25'b1110111010101001011001001;
    rom[29219] = 25'b1110111010101011110000110;
    rom[29220] = 25'b1110111010101110001001000;
    rom[29221] = 25'b1110111010110000100001110;
    rom[29222] = 25'b1110111010110010111010110;
    rom[29223] = 25'b1110111010110101010100100;
    rom[29224] = 25'b1110111010110111101110101;
    rom[29225] = 25'b1110111010111010001001001;
    rom[29226] = 25'b1110111010111100100100010;
    rom[29227] = 25'b1110111010111110111111111;
    rom[29228] = 25'b1110111011000001011011111;
    rom[29229] = 25'b1110111011000011111000011;
    rom[29230] = 25'b1110111011000110010101100;
    rom[29231] = 25'b1110111011001000110011000;
    rom[29232] = 25'b1110111011001011010001000;
    rom[29233] = 25'b1110111011001101101111100;
    rom[29234] = 25'b1110111011010000001110100;
    rom[29235] = 25'b1110111011010010101101111;
    rom[29236] = 25'b1110111011010101001101111;
    rom[29237] = 25'b1110111011010111101110010;
    rom[29238] = 25'b1110111011011010001111001;
    rom[29239] = 25'b1110111011011100110000100;
    rom[29240] = 25'b1110111011011111010010100;
    rom[29241] = 25'b1110111011100001110100111;
    rom[29242] = 25'b1110111011100100010111101;
    rom[29243] = 25'b1110111011100110111011001;
    rom[29244] = 25'b1110111011101001011110111;
    rom[29245] = 25'b1110111011101100000011010;
    rom[29246] = 25'b1110111011101110101000000;
    rom[29247] = 25'b1110111011110001001101010;
    rom[29248] = 25'b1110111011110011110011001;
    rom[29249] = 25'b1110111011110110011001011;
    rom[29250] = 25'b1110111011111001000000001;
    rom[29251] = 25'b1110111011111011100111011;
    rom[29252] = 25'b1110111011111110001111001;
    rom[29253] = 25'b1110111100000000110111011;
    rom[29254] = 25'b1110111100000011100000001;
    rom[29255] = 25'b1110111100000110001001010;
    rom[29256] = 25'b1110111100001000110010111;
    rom[29257] = 25'b1110111100001011011101001;
    rom[29258] = 25'b1110111100001110000111110;
    rom[29259] = 25'b1110111100010000110010111;
    rom[29260] = 25'b1110111100010011011110101;
    rom[29261] = 25'b1110111100010110001010101;
    rom[29262] = 25'b1110111100011000110111010;
    rom[29263] = 25'b1110111100011011100100011;
    rom[29264] = 25'b1110111100011110010010000;
    rom[29265] = 25'b1110111100100001000000001;
    rom[29266] = 25'b1110111100100011101110101;
    rom[29267] = 25'b1110111100100110011101110;
    rom[29268] = 25'b1110111100101001001101010;
    rom[29269] = 25'b1110111100101011111101011;
    rom[29270] = 25'b1110111100101110101101111;
    rom[29271] = 25'b1110111100110001011110111;
    rom[29272] = 25'b1110111100110100010000011;
    rom[29273] = 25'b1110111100110111000010011;
    rom[29274] = 25'b1110111100111001110100111;
    rom[29275] = 25'b1110111100111100100111111;
    rom[29276] = 25'b1110111100111111011011011;
    rom[29277] = 25'b1110111101000010001111011;
    rom[29278] = 25'b1110111101000101000011110;
    rom[29279] = 25'b1110111101000111111000110;
    rom[29280] = 25'b1110111101001010101110010;
    rom[29281] = 25'b1110111101001101100100001;
    rom[29282] = 25'b1110111101010000011010100;
    rom[29283] = 25'b1110111101010011010001100;
    rom[29284] = 25'b1110111101010110001000111;
    rom[29285] = 25'b1110111101011001000000110;
    rom[29286] = 25'b1110111101011011111001001;
    rom[29287] = 25'b1110111101011110110010000;
    rom[29288] = 25'b1110111101100001101011011;
    rom[29289] = 25'b1110111101100100100101010;
    rom[29290] = 25'b1110111101100111011111101;
    rom[29291] = 25'b1110111101101010011010011;
    rom[29292] = 25'b1110111101101101010101110;
    rom[29293] = 25'b1110111101110000010001101;
    rom[29294] = 25'b1110111101110011001101111;
    rom[29295] = 25'b1110111101110110001010110;
    rom[29296] = 25'b1110111101111001001000000;
    rom[29297] = 25'b1110111101111100000101111;
    rom[29298] = 25'b1110111101111111000100001;
    rom[29299] = 25'b1110111110000010000010111;
    rom[29300] = 25'b1110111110000101000010001;
    rom[29301] = 25'b1110111110001000000010000;
    rom[29302] = 25'b1110111110001011000010010;
    rom[29303] = 25'b1110111110001110000011000;
    rom[29304] = 25'b1110111110010001000100010;
    rom[29305] = 25'b1110111110010100000110000;
    rom[29306] = 25'b1110111110010111001000010;
    rom[29307] = 25'b1110111110011010001010111;
    rom[29308] = 25'b1110111110011101001110010;
    rom[29309] = 25'b1110111110100000010001111;
    rom[29310] = 25'b1110111110100011010110000;
    rom[29311] = 25'b1110111110100110011010111;
    rom[29312] = 25'b1110111110101001100000000;
    rom[29313] = 25'b1110111110101100100101101;
    rom[29314] = 25'b1110111110101111101011111;
    rom[29315] = 25'b1110111110110010110010100;
    rom[29316] = 25'b1110111110110101111001110;
    rom[29317] = 25'b1110111110111001000001011;
    rom[29318] = 25'b1110111110111100001001100;
    rom[29319] = 25'b1110111110111111010010010;
    rom[29320] = 25'b1110111111000010011011011;
    rom[29321] = 25'b1110111111000101100101000;
    rom[29322] = 25'b1110111111001000101111010;
    rom[29323] = 25'b1110111111001011111001111;
    rom[29324] = 25'b1110111111001111000101000;
    rom[29325] = 25'b1110111111010010010000101;
    rom[29326] = 25'b1110111111010101011100110;
    rom[29327] = 25'b1110111111011000101001011;
    rom[29328] = 25'b1110111111011011110110100;
    rom[29329] = 25'b1110111111011111000100001;
    rom[29330] = 25'b1110111111100010010010010;
    rom[29331] = 25'b1110111111100101100000110;
    rom[29332] = 25'b1110111111101000101111111;
    rom[29333] = 25'b1110111111101011111111100;
    rom[29334] = 25'b1110111111101111001111101;
    rom[29335] = 25'b1110111111110010100000010;
    rom[29336] = 25'b1110111111110101110001010;
    rom[29337] = 25'b1110111111111001000010111;
    rom[29338] = 25'b1110111111111100010100111;
    rom[29339] = 25'b1110111111111111100111100;
    rom[29340] = 25'b1111000000000010111010100;
    rom[29341] = 25'b1111000000000110001110001;
    rom[29342] = 25'b1111000000001001100010010;
    rom[29343] = 25'b1111000000001100110110110;
    rom[29344] = 25'b1111000000010000001011110;
    rom[29345] = 25'b1111000000010011100001011;
    rom[29346] = 25'b1111000000010110110111011;
    rom[29347] = 25'b1111000000011010001101111;
    rom[29348] = 25'b1111000000011101100101000;
    rom[29349] = 25'b1111000000100000111100100;
    rom[29350] = 25'b1111000000100100010100101;
    rom[29351] = 25'b1111000000100111101101001;
    rom[29352] = 25'b1111000000101011000110001;
    rom[29353] = 25'b1111000000101110011111110;
    rom[29354] = 25'b1111000000110001111001110;
    rom[29355] = 25'b1111000000110101010100010;
    rom[29356] = 25'b1111000000111000101111010;
    rom[29357] = 25'b1111000000111100001010110;
    rom[29358] = 25'b1111000000111111100110110;
    rom[29359] = 25'b1111000001000011000011011;
    rom[29360] = 25'b1111000001000110100000011;
    rom[29361] = 25'b1111000001001001111101111;
    rom[29362] = 25'b1111000001001101011011111;
    rom[29363] = 25'b1111000001010000111010011;
    rom[29364] = 25'b1111000001010100011001011;
    rom[29365] = 25'b1111000001010111111000111;
    rom[29366] = 25'b1111000001011011011000111;
    rom[29367] = 25'b1111000001011110111001011;
    rom[29368] = 25'b1111000001100010011010011;
    rom[29369] = 25'b1111000001100101111011111;
    rom[29370] = 25'b1111000001101001011101111;
    rom[29371] = 25'b1111000001101101000000011;
    rom[29372] = 25'b1111000001110000100011011;
    rom[29373] = 25'b1111000001110100000110111;
    rom[29374] = 25'b1111000001110111101010111;
    rom[29375] = 25'b1111000001111011001111011;
    rom[29376] = 25'b1111000001111110110100010;
    rom[29377] = 25'b1111000010000010011001111;
    rom[29378] = 25'b1111000010000101111111110;
    rom[29379] = 25'b1111000010001001100110010;
    rom[29380] = 25'b1111000010001101001101010;
    rom[29381] = 25'b1111000010010000110100110;
    rom[29382] = 25'b1111000010010100011100110;
    rom[29383] = 25'b1111000010011000000101010;
    rom[29384] = 25'b1111000010011011101110010;
    rom[29385] = 25'b1111000010011111010111101;
    rom[29386] = 25'b1111000010100011000001110;
    rom[29387] = 25'b1111000010100110101100010;
    rom[29388] = 25'b1111000010101010010111001;
    rom[29389] = 25'b1111000010101110000010101;
    rom[29390] = 25'b1111000010110001101110101;
    rom[29391] = 25'b1111000010110101011011001;
    rom[29392] = 25'b1111000010111001001000000;
    rom[29393] = 25'b1111000010111100110101100;
    rom[29394] = 25'b1111000011000000100011100;
    rom[29395] = 25'b1111000011000100010010000;
    rom[29396] = 25'b1111000011001000000001000;
    rom[29397] = 25'b1111000011001011110000100;
    rom[29398] = 25'b1111000011001111100000011;
    rom[29399] = 25'b1111000011010011010000111;
    rom[29400] = 25'b1111000011010111000001111;
    rom[29401] = 25'b1111000011011010110011011;
    rom[29402] = 25'b1111000011011110100101011;
    rom[29403] = 25'b1111000011100010010111111;
    rom[29404] = 25'b1111000011100110001010111;
    rom[29405] = 25'b1111000011101001111110010;
    rom[29406] = 25'b1111000011101101110010010;
    rom[29407] = 25'b1111000011110001100110110;
    rom[29408] = 25'b1111000011110101011011110;
    rom[29409] = 25'b1111000011111001010001010;
    rom[29410] = 25'b1111000011111101000111010;
    rom[29411] = 25'b1111000100000000111101110;
    rom[29412] = 25'b1111000100000100110100110;
    rom[29413] = 25'b1111000100001000101100001;
    rom[29414] = 25'b1111000100001100100100010;
    rom[29415] = 25'b1111000100010000011100110;
    rom[29416] = 25'b1111000100010100010101101;
    rom[29417] = 25'b1111000100011000001111010;
    rom[29418] = 25'b1111000100011100001001010;
    rom[29419] = 25'b1111000100100000000011101;
    rom[29420] = 25'b1111000100100011111110110;
    rom[29421] = 25'b1111000100100111111010001;
    rom[29422] = 25'b1111000100101011110110001;
    rom[29423] = 25'b1111000100101111110010101;
    rom[29424] = 25'b1111000100110011101111101;
    rom[29425] = 25'b1111000100110111101101001;
    rom[29426] = 25'b1111000100111011101011010;
    rom[29427] = 25'b1111000100111111101001101;
    rom[29428] = 25'b1111000101000011101000110;
    rom[29429] = 25'b1111000101000111101000010;
    rom[29430] = 25'b1111000101001011101000010;
    rom[29431] = 25'b1111000101001111101000110;
    rom[29432] = 25'b1111000101010011101001110;
    rom[29433] = 25'b1111000101010111101011010;
    rom[29434] = 25'b1111000101011011101101010;
    rom[29435] = 25'b1111000101011111101111111;
    rom[29436] = 25'b1111000101100011110010110;
    rom[29437] = 25'b1111000101100111110110010;
    rom[29438] = 25'b1111000101101011111010011;
    rom[29439] = 25'b1111000101101111111110111;
    rom[29440] = 25'b1111000101110100000011111;
    rom[29441] = 25'b1111000101111000001001100;
    rom[29442] = 25'b1111000101111100001111100;
    rom[29443] = 25'b1111000110000000010110000;
    rom[29444] = 25'b1111000110000100011101001;
    rom[29445] = 25'b1111000110001000100100101;
    rom[29446] = 25'b1111000110001100101100101;
    rom[29447] = 25'b1111000110010000110101001;
    rom[29448] = 25'b1111000110010100111110010;
    rom[29449] = 25'b1111000110011001000111110;
    rom[29450] = 25'b1111000110011101010001110;
    rom[29451] = 25'b1111000110100001011100011;
    rom[29452] = 25'b1111000110100101100111011;
    rom[29453] = 25'b1111000110101001110010111;
    rom[29454] = 25'b1111000110101101111111000;
    rom[29455] = 25'b1111000110110010001011100;
    rom[29456] = 25'b1111000110110110011000101;
    rom[29457] = 25'b1111000110111010100110010;
    rom[29458] = 25'b1111000110111110110100010;
    rom[29459] = 25'b1111000111000011000010110;
    rom[29460] = 25'b1111000111000111010001111;
    rom[29461] = 25'b1111000111001011100001100;
    rom[29462] = 25'b1111000111001111110001100;
    rom[29463] = 25'b1111000111010100000010001;
    rom[29464] = 25'b1111000111011000010011001;
    rom[29465] = 25'b1111000111011100100100110;
    rom[29466] = 25'b1111000111100000110110111;
    rom[29467] = 25'b1111000111100101001001100;
    rom[29468] = 25'b1111000111101001011100101;
    rom[29469] = 25'b1111000111101101110000001;
    rom[29470] = 25'b1111000111110010000100010;
    rom[29471] = 25'b1111000111110110011000111;
    rom[29472] = 25'b1111000111111010101110000;
    rom[29473] = 25'b1111000111111111000011100;
    rom[29474] = 25'b1111001000000011011001101;
    rom[29475] = 25'b1111001000000111110000010;
    rom[29476] = 25'b1111001000001100000111100;
    rom[29477] = 25'b1111001000010000011111000;
    rom[29478] = 25'b1111001000010100110111001;
    rom[29479] = 25'b1111001000011001001111110;
    rom[29480] = 25'b1111001000011101101000111;
    rom[29481] = 25'b1111001000100010000010100;
    rom[29482] = 25'b1111001000100110011100101;
    rom[29483] = 25'b1111001000101010110111010;
    rom[29484] = 25'b1111001000101111010010100;
    rom[29485] = 25'b1111001000110011101110000;
    rom[29486] = 25'b1111001000111000001010010;
    rom[29487] = 25'b1111001000111100100110111;
    rom[29488] = 25'b1111001001000001000100000;
    rom[29489] = 25'b1111001001000101100001101;
    rom[29490] = 25'b1111001001001001111111110;
    rom[29491] = 25'b1111001001001110011110100;
    rom[29492] = 25'b1111001001010010111101101;
    rom[29493] = 25'b1111001001010111011101010;
    rom[29494] = 25'b1111001001011011111101100;
    rom[29495] = 25'b1111001001100000011110001;
    rom[29496] = 25'b1111001001100100111111010;
    rom[29497] = 25'b1111001001101001100001000;
    rom[29498] = 25'b1111001001101110000011001;
    rom[29499] = 25'b1111001001110010100101111;
    rom[29500] = 25'b1111001001110111001001000;
    rom[29501] = 25'b1111001001111011101100101;
    rom[29502] = 25'b1111001010000000010000111;
    rom[29503] = 25'b1111001010000100110101100;
    rom[29504] = 25'b1111001010001001011010110;
    rom[29505] = 25'b1111001010001110000000100;
    rom[29506] = 25'b1111001010010010100110101;
    rom[29507] = 25'b1111001010010111001101011;
    rom[29508] = 25'b1111001010011011110100101;
    rom[29509] = 25'b1111001010100000011100010;
    rom[29510] = 25'b1111001010100101000100100;
    rom[29511] = 25'b1111001010101001101101010;
    rom[29512] = 25'b1111001010101110010110011;
    rom[29513] = 25'b1111001010110011000000001;
    rom[29514] = 25'b1111001010110111101010011;
    rom[29515] = 25'b1111001010111100010101000;
    rom[29516] = 25'b1111001011000001000000011;
    rom[29517] = 25'b1111001011000101101100000;
    rom[29518] = 25'b1111001011001010011000010;
    rom[29519] = 25'b1111001011001111000101001;
    rom[29520] = 25'b1111001011010011110010010;
    rom[29521] = 25'b1111001011011000100000000;
    rom[29522] = 25'b1111001011011101001110010;
    rom[29523] = 25'b1111001011100001111101000;
    rom[29524] = 25'b1111001011100110101100010;
    rom[29525] = 25'b1111001011101011011100000;
    rom[29526] = 25'b1111001011110000001100010;
    rom[29527] = 25'b1111001011110100111101000;
    rom[29528] = 25'b1111001011111001101110010;
    rom[29529] = 25'b1111001011111110100000000;
    rom[29530] = 25'b1111001100000011010010011;
    rom[29531] = 25'b1111001100001000000101001;
    rom[29532] = 25'b1111001100001100111000011;
    rom[29533] = 25'b1111001100010001101100001;
    rom[29534] = 25'b1111001100010110100000100;
    rom[29535] = 25'b1111001100011011010101010;
    rom[29536] = 25'b1111001100100000001010100;
    rom[29537] = 25'b1111001100100101000000011;
    rom[29538] = 25'b1111001100101001110110101;
    rom[29539] = 25'b1111001100101110101101011;
    rom[29540] = 25'b1111001100110011100100110;
    rom[29541] = 25'b1111001100111000011100100;
    rom[29542] = 25'b1111001100111101010100111;
    rom[29543] = 25'b1111001101000010001101101;
    rom[29544] = 25'b1111001101000111000110111;
    rom[29545] = 25'b1111001101001100000000101;
    rom[29546] = 25'b1111001101010000111011000;
    rom[29547] = 25'b1111001101010101110101111;
    rom[29548] = 25'b1111001101011010110001010;
    rom[29549] = 25'b1111001101011111101101000;
    rom[29550] = 25'b1111001101100100101001011;
    rom[29551] = 25'b1111001101101001100110001;
    rom[29552] = 25'b1111001101101110100011011;
    rom[29553] = 25'b1111001101110011100001011;
    rom[29554] = 25'b1111001101111000011111101;
    rom[29555] = 25'b1111001101111101011110100;
    rom[29556] = 25'b1111001110000010011101110;
    rom[29557] = 25'b1111001110000111011101101;
    rom[29558] = 25'b1111001110001100011110000;
    rom[29559] = 25'b1111001110010001011110111;
    rom[29560] = 25'b1111001110010110100000001;
    rom[29561] = 25'b1111001110011011100010000;
    rom[29562] = 25'b1111001110100000100100011;
    rom[29563] = 25'b1111001110100101100111010;
    rom[29564] = 25'b1111001110101010101010101;
    rom[29565] = 25'b1111001110101111101110100;
    rom[29566] = 25'b1111001110110100110010110;
    rom[29567] = 25'b1111001110111001110111110;
    rom[29568] = 25'b1111001110111110111101000;
    rom[29569] = 25'b1111001111000100000010111;
    rom[29570] = 25'b1111001111001001001001010;
    rom[29571] = 25'b1111001111001110010000001;
    rom[29572] = 25'b1111001111010011010111100;
    rom[29573] = 25'b1111001111011000011111011;
    rom[29574] = 25'b1111001111011101100111110;
    rom[29575] = 25'b1111001111100010110000101;
    rom[29576] = 25'b1111001111100111111010000;
    rom[29577] = 25'b1111001111101101000011111;
    rom[29578] = 25'b1111001111110010001110010;
    rom[29579] = 25'b1111001111110111011001001;
    rom[29580] = 25'b1111001111111100100100100;
    rom[29581] = 25'b1111010000000001110000011;
    rom[29582] = 25'b1111010000000110111100110;
    rom[29583] = 25'b1111010000001100001001110;
    rom[29584] = 25'b1111010000010001010111001;
    rom[29585] = 25'b1111010000010110100101000;
    rom[29586] = 25'b1111010000011011110011011;
    rom[29587] = 25'b1111010000100001000010010;
    rom[29588] = 25'b1111010000100110010001110;
    rom[29589] = 25'b1111010000101011100001101;
    rom[29590] = 25'b1111010000110000110010000;
    rom[29591] = 25'b1111010000110110000010111;
    rom[29592] = 25'b1111010000111011010100010;
    rom[29593] = 25'b1111010001000000100110010;
    rom[29594] = 25'b1111010001000101111000100;
    rom[29595] = 25'b1111010001001011001011100;
    rom[29596] = 25'b1111010001010000011110111;
    rom[29597] = 25'b1111010001010101110010110;
    rom[29598] = 25'b1111010001011011000111010;
    rom[29599] = 25'b1111010001100000011100001;
    rom[29600] = 25'b1111010001100101110001100;
    rom[29601] = 25'b1111010001101011000111011;
    rom[29602] = 25'b1111010001110000011101111;
    rom[29603] = 25'b1111010001110101110100110;
    rom[29604] = 25'b1111010001111011001100001;
    rom[29605] = 25'b1111010010000000100100001;
    rom[29606] = 25'b1111010010000101111100100;
    rom[29607] = 25'b1111010010001011010101011;
    rom[29608] = 25'b1111010010010000101110111;
    rom[29609] = 25'b1111010010010110001000110;
    rom[29610] = 25'b1111010010011011100011001;
    rom[29611] = 25'b1111010010100000111110000;
    rom[29612] = 25'b1111010010100110011001100;
    rom[29613] = 25'b1111010010101011110101011;
    rom[29614] = 25'b1111010010110001010001111;
    rom[29615] = 25'b1111010010110110101110110;
    rom[29616] = 25'b1111010010111100001100001;
    rom[29617] = 25'b1111010011000001101010000;
    rom[29618] = 25'b1111010011000111001000100;
    rom[29619] = 25'b1111010011001100100111011;
    rom[29620] = 25'b1111010011010010000110110;
    rom[29621] = 25'b1111010011010111100110110;
    rom[29622] = 25'b1111010011011101000111001;
    rom[29623] = 25'b1111010011100010101000000;
    rom[29624] = 25'b1111010011101000001001100;
    rom[29625] = 25'b1111010011101101101011010;
    rom[29626] = 25'b1111010011110011001101110;
    rom[29627] = 25'b1111010011111000110000101;
    rom[29628] = 25'b1111010011111110010100001;
    rom[29629] = 25'b1111010100000011111000000;
    rom[29630] = 25'b1111010100001001011100011;
    rom[29631] = 25'b1111010100001111000001010;
    rom[29632] = 25'b1111010100010100100110110;
    rom[29633] = 25'b1111010100011010001100101;
    rom[29634] = 25'b1111010100011111110011000;
    rom[29635] = 25'b1111010100100101011010000;
    rom[29636] = 25'b1111010100101011000001010;
    rom[29637] = 25'b1111010100110000101001010;
    rom[29638] = 25'b1111010100110110010001101;
    rom[29639] = 25'b1111010100111011111010100;
    rom[29640] = 25'b1111010101000001100100000;
    rom[29641] = 25'b1111010101000111001101111;
    rom[29642] = 25'b1111010101001100111000010;
    rom[29643] = 25'b1111010101010010100011001;
    rom[29644] = 25'b1111010101011000001110100;
    rom[29645] = 25'b1111010101011101111010011;
    rom[29646] = 25'b1111010101100011100110110;
    rom[29647] = 25'b1111010101101001010011110;
    rom[29648] = 25'b1111010101101111000001000;
    rom[29649] = 25'b1111010101110100101110111;
    rom[29650] = 25'b1111010101111010011101010;
    rom[29651] = 25'b1111010110000000001100010;
    rom[29652] = 25'b1111010110000101111011101;
    rom[29653] = 25'b1111010110001011101011100;
    rom[29654] = 25'b1111010110010001011011111;
    rom[29655] = 25'b1111010110010111001100101;
    rom[29656] = 25'b1111010110011100111110001;
    rom[29657] = 25'b1111010110100010101111111;
    rom[29658] = 25'b1111010110101000100010010;
    rom[29659] = 25'b1111010110101110010101001;
    rom[29660] = 25'b1111010110110100001000100;
    rom[29661] = 25'b1111010110111001111100011;
    rom[29662] = 25'b1111010110111111110000110;
    rom[29663] = 25'b1111010111000101100101100;
    rom[29664] = 25'b1111010111001011011010111;
    rom[29665] = 25'b1111010111010001010000110;
    rom[29666] = 25'b1111010111010111000111000;
    rom[29667] = 25'b1111010111011100111101111;
    rom[29668] = 25'b1111010111100010110101001;
    rom[29669] = 25'b1111010111101000101101000;
    rom[29670] = 25'b1111010111101110100101010;
    rom[29671] = 25'b1111010111110100011110001;
    rom[29672] = 25'b1111010111111010010111100;
    rom[29673] = 25'b1111011000000000010001010;
    rom[29674] = 25'b1111011000000110001011101;
    rom[29675] = 25'b1111011000001100000110011;
    rom[29676] = 25'b1111011000010010000001101;
    rom[29677] = 25'b1111011000010111111101100;
    rom[29678] = 25'b1111011000011101111001110;
    rom[29679] = 25'b1111011000100011110110101;
    rom[29680] = 25'b1111011000101001110011110;
    rom[29681] = 25'b1111011000101111110001101;
    rom[29682] = 25'b1111011000110101101111111;
    rom[29683] = 25'b1111011000111011101110101;
    rom[29684] = 25'b1111011001000001101110000;
    rom[29685] = 25'b1111011001000111101101101;
    rom[29686] = 25'b1111011001001101101110000;
    rom[29687] = 25'b1111011001010011101110110;
    rom[29688] = 25'b1111011001011001101111111;
    rom[29689] = 25'b1111011001011111110001101;
    rom[29690] = 25'b1111011001100101110011111;
    rom[29691] = 25'b1111011001101011110110101;
    rom[29692] = 25'b1111011001110001111001111;
    rom[29693] = 25'b1111011001110111111101100;
    rom[29694] = 25'b1111011001111110000001110;
    rom[29695] = 25'b1111011010000100000110100;
    rom[29696] = 25'b1111011010001010001011101;
    rom[29697] = 25'b1111011010010000010001011;
    rom[29698] = 25'b1111011010010110010111100;
    rom[29699] = 25'b1111011010011100011110010;
    rom[29700] = 25'b1111011010100010100101011;
    rom[29701] = 25'b1111011010101000101101000;
    rom[29702] = 25'b1111011010101110110101010;
    rom[29703] = 25'b1111011010110100111101111;
    rom[29704] = 25'b1111011010111011000111000;
    rom[29705] = 25'b1111011011000001010000101;
    rom[29706] = 25'b1111011011000111011010110;
    rom[29707] = 25'b1111011011001101100101011;
    rom[29708] = 25'b1111011011010011110000100;
    rom[29709] = 25'b1111011011011001111100001;
    rom[29710] = 25'b1111011011100000001000010;
    rom[29711] = 25'b1111011011100110010100111;
    rom[29712] = 25'b1111011011101100100001111;
    rom[29713] = 25'b1111011011110010101111100;
    rom[29714] = 25'b1111011011111000111101101;
    rom[29715] = 25'b1111011011111111001100001;
    rom[29716] = 25'b1111011100000101011011010;
    rom[29717] = 25'b1111011100001011101010110;
    rom[29718] = 25'b1111011100010001111010110;
    rom[29719] = 25'b1111011100011000001011010;
    rom[29720] = 25'b1111011100011110011100011;
    rom[29721] = 25'b1111011100100100101101111;
    rom[29722] = 25'b1111011100101010111111111;
    rom[29723] = 25'b1111011100110001010010011;
    rom[29724] = 25'b1111011100110111100101011;
    rom[29725] = 25'b1111011100111101111000110;
    rom[29726] = 25'b1111011101000100001100110;
    rom[29727] = 25'b1111011101001010100001010;
    rom[29728] = 25'b1111011101010000110110010;
    rom[29729] = 25'b1111011101010111001011101;
    rom[29730] = 25'b1111011101011101100001101;
    rom[29731] = 25'b1111011101100011111000000;
    rom[29732] = 25'b1111011101101010001110111;
    rom[29733] = 25'b1111011101110000100110011;
    rom[29734] = 25'b1111011101110110111110010;
    rom[29735] = 25'b1111011101111101010110101;
    rom[29736] = 25'b1111011110000011101111100;
    rom[29737] = 25'b1111011110001010001000111;
    rom[29738] = 25'b1111011110010000100010110;
    rom[29739] = 25'b1111011110010110111101001;
    rom[29740] = 25'b1111011110011101011000000;
    rom[29741] = 25'b1111011110100011110011010;
    rom[29742] = 25'b1111011110101010001111001;
    rom[29743] = 25'b1111011110110000101011011;
    rom[29744] = 25'b1111011110110111001000001;
    rom[29745] = 25'b1111011110111101100101100;
    rom[29746] = 25'b1111011111000100000011010;
    rom[29747] = 25'b1111011111001010100001100;
    rom[29748] = 25'b1111011111010001000000010;
    rom[29749] = 25'b1111011111010111011111100;
    rom[29750] = 25'b1111011111011101111111010;
    rom[29751] = 25'b1111011111100100011111100;
    rom[29752] = 25'b1111011111101011000000001;
    rom[29753] = 25'b1111011111110001100001010;
    rom[29754] = 25'b1111011111111000000011000;
    rom[29755] = 25'b1111011111111110100101001;
    rom[29756] = 25'b1111100000000101000111110;
    rom[29757] = 25'b1111100000001011101010111;
    rom[29758] = 25'b1111100000010010001110101;
    rom[29759] = 25'b1111100000011000110010110;
    rom[29760] = 25'b1111100000011111010111010;
    rom[29761] = 25'b1111100000100101111100011;
    rom[29762] = 25'b1111100000101100100010000;
    rom[29763] = 25'b1111100000110011001000000;
    rom[29764] = 25'b1111100000111001101110101;
    rom[29765] = 25'b1111100001000000010101101;
    rom[29766] = 25'b1111100001000110111101001;
    rom[29767] = 25'b1111100001001101100101001;
    rom[29768] = 25'b1111100001010100001101101;
    rom[29769] = 25'b1111100001011010110110101;
    rom[29770] = 25'b1111100001100001100000000;
    rom[29771] = 25'b1111100001101000001010000;
    rom[29772] = 25'b1111100001101110110100100;
    rom[29773] = 25'b1111100001110101011111011;
    rom[29774] = 25'b1111100001111100001010110;
    rom[29775] = 25'b1111100010000010110110101;
    rom[29776] = 25'b1111100010001001100011000;
    rom[29777] = 25'b1111100010010000010000000;
    rom[29778] = 25'b1111100010010110111101010;
    rom[29779] = 25'b1111100010011101101011001;
    rom[29780] = 25'b1111100010100100011001011;
    rom[29781] = 25'b1111100010101011001000010;
    rom[29782] = 25'b1111100010110001110111100;
    rom[29783] = 25'b1111100010111000100111010;
    rom[29784] = 25'b1111100010111111010111100;
    rom[29785] = 25'b1111100011000110001000010;
    rom[29786] = 25'b1111100011001100111001100;
    rom[29787] = 25'b1111100011010011101011001;
    rom[29788] = 25'b1111100011011010011101011;
    rom[29789] = 25'b1111100011100001010000000;
    rom[29790] = 25'b1111100011101000000011001;
    rom[29791] = 25'b1111100011101110110110110;
    rom[29792] = 25'b1111100011110101101010111;
    rom[29793] = 25'b1111100011111100011111100;
    rom[29794] = 25'b1111100100000011010100101;
    rom[29795] = 25'b1111100100001010001010001;
    rom[29796] = 25'b1111100100010001000000010;
    rom[29797] = 25'b1111100100010111110110110;
    rom[29798] = 25'b1111100100011110101101110;
    rom[29799] = 25'b1111100100100101100101010;
    rom[29800] = 25'b1111100100101100011101010;
    rom[29801] = 25'b1111100100110011010101110;
    rom[29802] = 25'b1111100100111010001110101;
    rom[29803] = 25'b1111100101000001001000000;
    rom[29804] = 25'b1111100101001000000010000;
    rom[29805] = 25'b1111100101001110111100011;
    rom[29806] = 25'b1111100101010101110111001;
    rom[29807] = 25'b1111100101011100110010101;
    rom[29808] = 25'b1111100101100011101110011;
    rom[29809] = 25'b1111100101101010101010101;
    rom[29810] = 25'b1111100101110001100111100;
    rom[29811] = 25'b1111100101111000100100110;
    rom[29812] = 25'b1111100101111111100010100;
    rom[29813] = 25'b1111100110000110100000110;
    rom[29814] = 25'b1111100110001101011111011;
    rom[29815] = 25'b1111100110010100011110101;
    rom[29816] = 25'b1111100110011011011110010;
    rom[29817] = 25'b1111100110100010011110011;
    rom[29818] = 25'b1111100110101001011111000;
    rom[29819] = 25'b1111100110110000100000001;
    rom[29820] = 25'b1111100110110111100001101;
    rom[29821] = 25'b1111100110111110100011110;
    rom[29822] = 25'b1111100111000101100110010;
    rom[29823] = 25'b1111100111001100101001010;
    rom[29824] = 25'b1111100111010011101100110;
    rom[29825] = 25'b1111100111011010110000110;
    rom[29826] = 25'b1111100111100001110101010;
    rom[29827] = 25'b1111100111101000111010001;
    rom[29828] = 25'b1111100111101111111111100;
    rom[29829] = 25'b1111100111110111000101011;
    rom[29830] = 25'b1111100111111110001011110;
    rom[29831] = 25'b1111101000000101010010101;
    rom[29832] = 25'b1111101000001100011001111;
    rom[29833] = 25'b1111101000010011100001110;
    rom[29834] = 25'b1111101000011010101001111;
    rom[29835] = 25'b1111101000100001110010101;
    rom[29836] = 25'b1111101000101000111011111;
    rom[29837] = 25'b1111101000110000000101101;
    rom[29838] = 25'b1111101000110111001111110;
    rom[29839] = 25'b1111101000111110011010011;
    rom[29840] = 25'b1111101001000101100101100;
    rom[29841] = 25'b1111101001001100110001001;
    rom[29842] = 25'b1111101001010011111101010;
    rom[29843] = 25'b1111101001011011001001110;
    rom[29844] = 25'b1111101001100010010110110;
    rom[29845] = 25'b1111101001101001100100001;
    rom[29846] = 25'b1111101001110000110010001;
    rom[29847] = 25'b1111101001111000000000101;
    rom[29848] = 25'b1111101001111111001111100;
    rom[29849] = 25'b1111101010000110011110111;
    rom[29850] = 25'b1111101010001101101110110;
    rom[29851] = 25'b1111101010010100111111001;
    rom[29852] = 25'b1111101010011100010000000;
    rom[29853] = 25'b1111101010100011100001010;
    rom[29854] = 25'b1111101010101010110011000;
    rom[29855] = 25'b1111101010110010000101010;
    rom[29856] = 25'b1111101010111001010111111;
    rom[29857] = 25'b1111101011000000101011001;
    rom[29858] = 25'b1111101011000111111110110;
    rom[29859] = 25'b1111101011001111010010111;
    rom[29860] = 25'b1111101011010110100111100;
    rom[29861] = 25'b1111101011011101111100100;
    rom[29862] = 25'b1111101011100101010010000;
    rom[29863] = 25'b1111101011101100101000000;
    rom[29864] = 25'b1111101011110011111110100;
    rom[29865] = 25'b1111101011111011010101100;
    rom[29866] = 25'b1111101100000010101100111;
    rom[29867] = 25'b1111101100001010000100110;
    rom[29868] = 25'b1111101100010001011101001;
    rom[29869] = 25'b1111101100011000110101111;
    rom[29870] = 25'b1111101100100000001111010;
    rom[29871] = 25'b1111101100100111101001000;
    rom[29872] = 25'b1111101100101111000011010;
    rom[29873] = 25'b1111101100110110011110000;
    rom[29874] = 25'b1111101100111101111001001;
    rom[29875] = 25'b1111101101000101010100111;
    rom[29876] = 25'b1111101101001100110000111;
    rom[29877] = 25'b1111101101010100001101100;
    rom[29878] = 25'b1111101101011011101010101;
    rom[29879] = 25'b1111101101100011001000001;
    rom[29880] = 25'b1111101101101010100110001;
    rom[29881] = 25'b1111101101110010000100100;
    rom[29882] = 25'b1111101101111001100011011;
    rom[29883] = 25'b1111101110000001000010111;
    rom[29884] = 25'b1111101110001000100010110;
    rom[29885] = 25'b1111101110010000000011001;
    rom[29886] = 25'b1111101110010111100011111;
    rom[29887] = 25'b1111101110011111000101001;
    rom[29888] = 25'b1111101110100110100110111;
    rom[29889] = 25'b1111101110101110001001001;
    rom[29890] = 25'b1111101110110101101011110;
    rom[29891] = 25'b1111101110111101001110111;
    rom[29892] = 25'b1111101111000100110010100;
    rom[29893] = 25'b1111101111001100010110100;
    rom[29894] = 25'b1111101111010011111011001;
    rom[29895] = 25'b1111101111011011100000000;
    rom[29896] = 25'b1111101111100011000101100;
    rom[29897] = 25'b1111101111101010101011100;
    rom[29898] = 25'b1111101111110010010001110;
    rom[29899] = 25'b1111101111111001111000110;
    rom[29900] = 25'b1111110000000001100000000;
    rom[29901] = 25'b1111110000001001000111110;
    rom[29902] = 25'b1111110000010000110000001;
    rom[29903] = 25'b1111110000011000011000110;
    rom[29904] = 25'b1111110000100000000010000;
    rom[29905] = 25'b1111110000100111101011101;
    rom[29906] = 25'b1111110000101111010101101;
    rom[29907] = 25'b1111110000110111000000010;
    rom[29908] = 25'b1111110000111110101011010;
    rom[29909] = 25'b1111110001000110010110110;
    rom[29910] = 25'b1111110001001110000010110;
    rom[29911] = 25'b1111110001010101101111001;
    rom[29912] = 25'b1111110001011101011100000;
    rom[29913] = 25'b1111110001100101001001011;
    rom[29914] = 25'b1111110001101100110111001;
    rom[29915] = 25'b1111110001110100100101100;
    rom[29916] = 25'b1111110001111100010100010;
    rom[29917] = 25'b1111110010000100000011011;
    rom[29918] = 25'b1111110010001011110011000;
    rom[29919] = 25'b1111110010010011100011001;
    rom[29920] = 25'b1111110010011011010011110;
    rom[29921] = 25'b1111110010100011000100110;
    rom[29922] = 25'b1111110010101010110110010;
    rom[29923] = 25'b1111110010110010101000001;
    rom[29924] = 25'b1111110010111010011010101;
    rom[29925] = 25'b1111110011000010001101100;
    rom[29926] = 25'b1111110011001010000000110;
    rom[29927] = 25'b1111110011010001110100101;
    rom[29928] = 25'b1111110011011001101000111;
    rom[29929] = 25'b1111110011100001011101100;
    rom[29930] = 25'b1111110011101001010010110;
    rom[29931] = 25'b1111110011110001001000010;
    rom[29932] = 25'b1111110011111000111110100;
    rom[29933] = 25'b1111110100000000110101000;
    rom[29934] = 25'b1111110100001000101100000;
    rom[29935] = 25'b1111110100010000100011011;
    rom[29936] = 25'b1111110100011000011011011;
    rom[29937] = 25'b1111110100100000010011110;
    rom[29938] = 25'b1111110100101000001100100;
    rom[29939] = 25'b1111110100110000000101110;
    rom[29940] = 25'b1111110100110111111111100;
    rom[29941] = 25'b1111110100111111111001110;
    rom[29942] = 25'b1111110101000111110100011;
    rom[29943] = 25'b1111110101001111101111100;
    rom[29944] = 25'b1111110101010111101011001;
    rom[29945] = 25'b1111110101011111100111001;
    rom[29946] = 25'b1111110101100111100011101;
    rom[29947] = 25'b1111110101101111100000100;
    rom[29948] = 25'b1111110101110111011101111;
    rom[29949] = 25'b1111110101111111011011110;
    rom[29950] = 25'b1111110110000111011010000;
    rom[29951] = 25'b1111110110001111011000110;
    rom[29952] = 25'b1111110110010111011000000;
    rom[29953] = 25'b1111110110011111010111101;
    rom[29954] = 25'b1111110110100111010111110;
    rom[29955] = 25'b1111110110101111011000010;
    rom[29956] = 25'b1111110110110111011001010;
    rom[29957] = 25'b1111110110111111011010110;
    rom[29958] = 25'b1111110111000111011100110;
    rom[29959] = 25'b1111110111001111011111000;
    rom[29960] = 25'b1111110111010111100001111;
    rom[29961] = 25'b1111110111011111100101001;
    rom[29962] = 25'b1111110111100111101000111;
    rom[29963] = 25'b1111110111101111101101001;
    rom[29964] = 25'b1111110111110111110001110;
    rom[29965] = 25'b1111110111111111110110110;
    rom[29966] = 25'b1111111000000111111100010;
    rom[29967] = 25'b1111111000010000000010010;
    rom[29968] = 25'b1111111000011000001000101;
    rom[29969] = 25'b1111111000100000001111101;
    rom[29970] = 25'b1111111000101000010110111;
    rom[29971] = 25'b1111111000110000011110110;
    rom[29972] = 25'b1111111000111000100110111;
    rom[29973] = 25'b1111111001000000101111101;
    rom[29974] = 25'b1111111001001000111000110;
    rom[29975] = 25'b1111111001010001000010010;
    rom[29976] = 25'b1111111001011001001100010;
    rom[29977] = 25'b1111111001100001010110110;
    rom[29978] = 25'b1111111001101001100001101;
    rom[29979] = 25'b1111111001110001101101000;
    rom[29980] = 25'b1111111001111001111000111;
    rom[29981] = 25'b1111111010000010000101001;
    rom[29982] = 25'b1111111010001010010001111;
    rom[29983] = 25'b1111111010010010011111000;
    rom[29984] = 25'b1111111010011010101100101;
    rom[29985] = 25'b1111111010100010111010101;
    rom[29986] = 25'b1111111010101011001001001;
    rom[29987] = 25'b1111111010110011011000001;
    rom[29988] = 25'b1111111010111011100111100;
    rom[29989] = 25'b1111111011000011110111010;
    rom[29990] = 25'b1111111011001100000111100;
    rom[29991] = 25'b1111111011010100011000011;
    rom[29992] = 25'b1111111011011100101001100;
    rom[29993] = 25'b1111111011100100111011000;
    rom[29994] = 25'b1111111011101101001101001;
    rom[29995] = 25'b1111111011110101011111101;
    rom[29996] = 25'b1111111011111101110010100;
    rom[29997] = 25'b1111111100000110000101111;
    rom[29998] = 25'b1111111100001110011001110;
    rom[29999] = 25'b1111111100010110101110000;
    rom[30000] = 25'b1111111100011111000010110;
    rom[30001] = 25'b1111111100100111010111111;
    rom[30002] = 25'b1111111100101111101101100;
    rom[30003] = 25'b1111111100111000000011101;
    rom[30004] = 25'b1111111101000000011010000;
    rom[30005] = 25'b1111111101001000110001000;
    rom[30006] = 25'b1111111101010001001000011;
    rom[30007] = 25'b1111111101011001100000001;
    rom[30008] = 25'b1111111101100001111000011;
    rom[30009] = 25'b1111111101101010010001000;
    rom[30010] = 25'b1111111101110010101010010;
    rom[30011] = 25'b1111111101111011000011110;
    rom[30012] = 25'b1111111110000011011101110;
    rom[30013] = 25'b1111111110001011111000010;
    rom[30014] = 25'b1111111110010100010011000;
    rom[30015] = 25'b1111111110011100101110011;
    rom[30016] = 25'b1111111110100101001010001;
    rom[30017] = 25'b1111111110101101100110011;
    rom[30018] = 25'b1111111110110110000011000;
    rom[30019] = 25'b1111111110111110100000001;
    rom[30020] = 25'b1111111111000110111101101;
    rom[30021] = 25'b1111111111001111011011100;
    rom[30022] = 25'b1111111111010111111010000;
    rom[30023] = 25'b1111111111100000011000110;
    rom[30024] = 25'b1111111111101000111000000;
    rom[30025] = 25'b1111111111110001010111110;
    rom[30026] = 25'b1111111111111001110111110;
    rom[30027] = 25'b0000000000000010011000011;
    rom[30028] = 25'b0000000000001010111001011;
    rom[30029] = 25'b0000000000010011011010110;
    rom[30030] = 25'b0000000000011011111100101;
    rom[30031] = 25'b0000000000100100011111000;
    rom[30032] = 25'b0000000000101101000001101;
    rom[30033] = 25'b0000000000110101100100111;
    rom[30034] = 25'b0000000000111110001000100;
    rom[30035] = 25'b0000000001000110101100100;
    rom[30036] = 25'b0000000001001111010001000;
    rom[30037] = 25'b0000000001010111110101111;
    rom[30038] = 25'b0000000001100000011011010;
    rom[30039] = 25'b0000000001101001000001001;
    rom[30040] = 25'b0000000001110001100111010;
    rom[30041] = 25'b0000000001111010001110000;
    rom[30042] = 25'b0000000010000010110101000;
    rom[30043] = 25'b0000000010001011011100100;
    rom[30044] = 25'b0000000010010100000100011;
    rom[30045] = 25'b0000000010011100101100110;
    rom[30046] = 25'b0000000010100101010101101;
    rom[30047] = 25'b0000000010101101111110111;
    rom[30048] = 25'b0000000010110110101000100;
    rom[30049] = 25'b0000000010111111010010101;
    rom[30050] = 25'b0000000011000111111101001;
    rom[30051] = 25'b0000000011010000101000000;
    rom[30052] = 25'b0000000011011001010011011;
    rom[30053] = 25'b0000000011100001111111010;
    rom[30054] = 25'b0000000011101010101011100;
    rom[30055] = 25'b0000000011110011011000001;
    rom[30056] = 25'b0000000011111100000101010;
    rom[30057] = 25'b0000000100000100110010111;
    rom[30058] = 25'b0000000100001101100000110;
    rom[30059] = 25'b0000000100010110001111001;
    rom[30060] = 25'b0000000100011110111101111;
    rom[30061] = 25'b0000000100100111101101001;
    rom[30062] = 25'b0000000100110000011100110;
    rom[30063] = 25'b0000000100111001001100111;
    rom[30064] = 25'b0000000101000001111101011;
    rom[30065] = 25'b0000000101001010101110010;
    rom[30066] = 25'b0000000101010011011111110;
    rom[30067] = 25'b0000000101011100010001100;
    rom[30068] = 25'b0000000101100101000011110;
    rom[30069] = 25'b0000000101101101110110010;
    rom[30070] = 25'b0000000101110110101001011;
    rom[30071] = 25'b0000000101111111011100111;
    rom[30072] = 25'b0000000110001000010000110;
    rom[30073] = 25'b0000000110010001000101001;
    rom[30074] = 25'b0000000110011001111001111;
    rom[30075] = 25'b0000000110100010101111000;
    rom[30076] = 25'b0000000110101011100100101;
    rom[30077] = 25'b0000000110110100011010101;
    rom[30078] = 25'b0000000110111101010001001;
    rom[30079] = 25'b0000000111000110001000000;
    rom[30080] = 25'b0000000111001110111111010;
    rom[30081] = 25'b0000000111010111110111000;
    rom[30082] = 25'b0000000111100000101111001;
    rom[30083] = 25'b0000000111101001100111101;
    rom[30084] = 25'b0000000111110010100000101;
    rom[30085] = 25'b0000000111111011011010000;
    rom[30086] = 25'b0000001000000100010011111;
    rom[30087] = 25'b0000001000001101001110001;
    rom[30088] = 25'b0000001000010110001000110;
    rom[30089] = 25'b0000001000011111000011110;
    rom[30090] = 25'b0000001000100111111111011;
    rom[30091] = 25'b0000001000110000111011010;
    rom[30092] = 25'b0000001000111001110111101;
    rom[30093] = 25'b0000001001000010110100011;
    rom[30094] = 25'b0000001001001011110001100;
    rom[30095] = 25'b0000001001010100101111000;
    rom[30096] = 25'b0000001001011101101101000;
    rom[30097] = 25'b0000001001100110101011011;
    rom[30098] = 25'b0000001001101111101010010;
    rom[30099] = 25'b0000001001111000101001100;
    rom[30100] = 25'b0000001010000001101001010;
    rom[30101] = 25'b0000001010001010101001010;
    rom[30102] = 25'b0000001010010011101001110;
    rom[30103] = 25'b0000001010011100101010101;
    rom[30104] = 25'b0000001010100101101100000;
    rom[30105] = 25'b0000001010101110101101110;
    rom[30106] = 25'b0000001010110111101111111;
    rom[30107] = 25'b0000001011000000110010011;
    rom[30108] = 25'b0000001011001001110101011;
    rom[30109] = 25'b0000001011010010111000110;
    rom[30110] = 25'b0000001011011011111100100;
    rom[30111] = 25'b0000001011100101000000110;
    rom[30112] = 25'b0000001011101110000101100;
    rom[30113] = 25'b0000001011110111001010100;
    rom[30114] = 25'b0000001100000000001111111;
    rom[30115] = 25'b0000001100001001010101111;
    rom[30116] = 25'b0000001100010010011100001;
    rom[30117] = 25'b0000001100011011100010110;
    rom[30118] = 25'b0000001100100100101001111;
    rom[30119] = 25'b0000001100101101110001011;
    rom[30120] = 25'b0000001100110110111001010;
    rom[30121] = 25'b0000001101000000000001101;
    rom[30122] = 25'b0000001101001001001010010;
    rom[30123] = 25'b0000001101010010010011100;
    rom[30124] = 25'b0000001101011011011101000;
    rom[30125] = 25'b0000001101100100100111000;
    rom[30126] = 25'b0000001101101101110001011;
    rom[30127] = 25'b0000001101110110111100001;
    rom[30128] = 25'b0000001110000000000111011;
    rom[30129] = 25'b0000001110001001010010111;
    rom[30130] = 25'b0000001110010010011110111;
    rom[30131] = 25'b0000001110011011101011011;
    rom[30132] = 25'b0000001110100100111000001;
    rom[30133] = 25'b0000001110101110000101010;
    rom[30134] = 25'b0000001110110111010011000;
    rom[30135] = 25'b0000001111000000100001000;
    rom[30136] = 25'b0000001111001001101111011;
    rom[30137] = 25'b0000001111010010111110010;
    rom[30138] = 25'b0000001111011100001101100;
    rom[30139] = 25'b0000001111100101011101001;
    rom[30140] = 25'b0000001111101110101101001;
    rom[30141] = 25'b0000001111110111111101101;
    rom[30142] = 25'b0000010000000001001110100;
    rom[30143] = 25'b0000010000001010011111110;
    rom[30144] = 25'b0000010000010011110001011;
    rom[30145] = 25'b0000010000011101000011100;
    rom[30146] = 25'b0000010000100110010101111;
    rom[30147] = 25'b0000010000101111101000110;
    rom[30148] = 25'b0000010000111000111100001;
    rom[30149] = 25'b0000010001000010001111110;
    rom[30150] = 25'b0000010001001011100011111;
    rom[30151] = 25'b0000010001010100111000010;
    rom[30152] = 25'b0000010001011110001101001;
    rom[30153] = 25'b0000010001100111100010011;
    rom[30154] = 25'b0000010001110000111000001;
    rom[30155] = 25'b0000010001111010001110001;
    rom[30156] = 25'b0000010010000011100100101;
    rom[30157] = 25'b0000010010001100111011100;
    rom[30158] = 25'b0000010010010110010010110;
    rom[30159] = 25'b0000010010011111101010011;
    rom[30160] = 25'b0000010010101001000010100;
    rom[30161] = 25'b0000010010110010011011000;
    rom[30162] = 25'b0000010010111011110011110;
    rom[30163] = 25'b0000010011000101001101000;
    rom[30164] = 25'b0000010011001110100110101;
    rom[30165] = 25'b0000010011011000000000110;
    rom[30166] = 25'b0000010011100001011011001;
    rom[30167] = 25'b0000010011101010110110000;
    rom[30168] = 25'b0000010011110100010001010;
    rom[30169] = 25'b0000010011111101101100110;
    rom[30170] = 25'b0000010100000111001000111;
    rom[30171] = 25'b0000010100010000100101010;
    rom[30172] = 25'b0000010100011010000010001;
    rom[30173] = 25'b0000010100100011011111010;
    rom[30174] = 25'b0000010100101100111100111;
    rom[30175] = 25'b0000010100110110011010111;
    rom[30176] = 25'b0000010100111111111001010;
    rom[30177] = 25'b0000010101001001010111111;
    rom[30178] = 25'b0000010101010010110111001;
    rom[30179] = 25'b0000010101011100010110110;
    rom[30180] = 25'b0000010101100101110110101;
    rom[30181] = 25'b0000010101101111010111000;
    rom[30182] = 25'b0000010101111000110111101;
    rom[30183] = 25'b0000010110000010011000110;
    rom[30184] = 25'b0000010110001011111010010;
    rom[30185] = 25'b0000010110010101011100010;
    rom[30186] = 25'b0000010110011110111110100;
    rom[30187] = 25'b0000010110101000100001001;
    rom[30188] = 25'b0000010110110010000100001;
    rom[30189] = 25'b0000010110111011100111101;
    rom[30190] = 25'b0000010111000101001011100;
    rom[30191] = 25'b0000010111001110101111110;
    rom[30192] = 25'b0000010111011000010100010;
    rom[30193] = 25'b0000010111100001111001010;
    rom[30194] = 25'b0000010111101011011110101;
    rom[30195] = 25'b0000010111110101000100011;
    rom[30196] = 25'b0000010111111110101010101;
    rom[30197] = 25'b0000011000001000010001001;
    rom[30198] = 25'b0000011000010001111000000;
    rom[30199] = 25'b0000011000011011011111011;
    rom[30200] = 25'b0000011000100101000111000;
    rom[30201] = 25'b0000011000101110101111000;
    rom[30202] = 25'b0000011000111000010111101;
    rom[30203] = 25'b0000011001000010000000011;
    rom[30204] = 25'b0000011001001011101001101;
    rom[30205] = 25'b0000011001010101010011010;
    rom[30206] = 25'b0000011001011110111101010;
    rom[30207] = 25'b0000011001101000100111101;
    rom[30208] = 25'b0000011001110010010010011;
    rom[30209] = 25'b0000011001111011111101100;
    rom[30210] = 25'b0000011010000101101001000;
    rom[30211] = 25'b0000011010001111010100111;
    rom[30212] = 25'b0000011010011001000001001;
    rom[30213] = 25'b0000011010100010101101111;
    rom[30214] = 25'b0000011010101100011010111;
    rom[30215] = 25'b0000011010110110001000010;
    rom[30216] = 25'b0000011010111111110110001;
    rom[30217] = 25'b0000011011001001100100010;
    rom[30218] = 25'b0000011011010011010010110;
    rom[30219] = 25'b0000011011011101000001110;
    rom[30220] = 25'b0000011011100110110001000;
    rom[30221] = 25'b0000011011110000100000110;
    rom[30222] = 25'b0000011011111010010000110;
    rom[30223] = 25'b0000011100000100000001010;
    rom[30224] = 25'b0000011100001101110010000;
    rom[30225] = 25'b0000011100010111100011010;
    rom[30226] = 25'b0000011100100001010100110;
    rom[30227] = 25'b0000011100101011000110110;
    rom[30228] = 25'b0000011100110100111001001;
    rom[30229] = 25'b0000011100111110101011110;
    rom[30230] = 25'b0000011101001000011110110;
    rom[30231] = 25'b0000011101010010010010010;
    rom[30232] = 25'b0000011101011100000110000;
    rom[30233] = 25'b0000011101100101111010010;
    rom[30234] = 25'b0000011101101111101110110;
    rom[30235] = 25'b0000011101111001100011101;
    rom[30236] = 25'b0000011110000011011001000;
    rom[30237] = 25'b0000011110001101001110110;
    rom[30238] = 25'b0000011110010111000100110;
    rom[30239] = 25'b0000011110100000111011001;
    rom[30240] = 25'b0000011110101010110001111;
    rom[30241] = 25'b0000011110110100101001001;
    rom[30242] = 25'b0000011110111110100000101;
    rom[30243] = 25'b0000011111001000011000100;
    rom[30244] = 25'b0000011111010010010000110;
    rom[30245] = 25'b0000011111011100001001011;
    rom[30246] = 25'b0000011111100110000010011;
    rom[30247] = 25'b0000011111101111111011110;
    rom[30248] = 25'b0000011111111001110101100;
    rom[30249] = 25'b0000100000000011101111101;
    rom[30250] = 25'b0000100000001101101010001;
    rom[30251] = 25'b0000100000010111100100111;
    rom[30252] = 25'b0000100000100001100000000;
    rom[30253] = 25'b0000100000101011011011101;
    rom[30254] = 25'b0000100000110101010111101;
    rom[30255] = 25'b0000100000111111010011111;
    rom[30256] = 25'b0000100001001001010000101;
    rom[30257] = 25'b0000100001010011001101100;
    rom[30258] = 25'b0000100001011101001010111;
    rom[30259] = 25'b0000100001100111001000110;
    rom[30260] = 25'b0000100001110001000110111;
    rom[30261] = 25'b0000100001111011000101011;
    rom[30262] = 25'b0000100010000101000100001;
    rom[30263] = 25'b0000100010001111000011011;
    rom[30264] = 25'b0000100010011001000011000;
    rom[30265] = 25'b0000100010100011000010111;
    rom[30266] = 25'b0000100010101101000011001;
    rom[30267] = 25'b0000100010110111000011111;
    rom[30268] = 25'b0000100011000001000100111;
    rom[30269] = 25'b0000100011001011000110001;
    rom[30270] = 25'b0000100011010101000111111;
    rom[30271] = 25'b0000100011011111001010000;
    rom[30272] = 25'b0000100011101001001100100;
    rom[30273] = 25'b0000100011110011001111010;
    rom[30274] = 25'b0000100011111101010010100;
    rom[30275] = 25'b0000100100000111010110000;
    rom[30276] = 25'b0000100100010001011001111;
    rom[30277] = 25'b0000100100011011011110001;
    rom[30278] = 25'b0000100100100101100010101;
    rom[30279] = 25'b0000100100101111100111101;
    rom[30280] = 25'b0000100100111001101101000;
    rom[30281] = 25'b0000100101000011110010100;
    rom[30282] = 25'b0000100101001101111000101;
    rom[30283] = 25'b0000100101010111111111000;
    rom[30284] = 25'b0000100101100010000101110;
    rom[30285] = 25'b0000100101101100001100111;
    rom[30286] = 25'b0000100101110110010100010;
    rom[30287] = 25'b0000100110000000011100000;
    rom[30288] = 25'b0000100110001010100100010;
    rom[30289] = 25'b0000100110010100101100101;
    rom[30290] = 25'b0000100110011110110101100;
    rom[30291] = 25'b0000100110101000111110101;
    rom[30292] = 25'b0000100110110011001000010;
    rom[30293] = 25'b0000100110111101010010001;
    rom[30294] = 25'b0000100111000111011100011;
    rom[30295] = 25'b0000100111010001100111000;
    rom[30296] = 25'b0000100111011011110010000;
    rom[30297] = 25'b0000100111100101111101010;
    rom[30298] = 25'b0000100111110000001000111;
    rom[30299] = 25'b0000100111111010010100111;
    rom[30300] = 25'b0000101000000100100001010;
    rom[30301] = 25'b0000101000001110101110000;
    rom[30302] = 25'b0000101000011000111011000;
    rom[30303] = 25'b0000101000100011001000011;
    rom[30304] = 25'b0000101000101101010110001;
    rom[30305] = 25'b0000101000110111100100001;
    rom[30306] = 25'b0000101001000001110010101;
    rom[30307] = 25'b0000101001001100000001011;
    rom[30308] = 25'b0000101001010110010000101;
    rom[30309] = 25'b0000101001100000100000000;
    rom[30310] = 25'b0000101001101010101111110;
    rom[30311] = 25'b0000101001110101000000000;
    rom[30312] = 25'b0000101001111111010000100;
    rom[30313] = 25'b0000101010001001100001011;
    rom[30314] = 25'b0000101010010011110010100;
    rom[30315] = 25'b0000101010011110000100000;
    rom[30316] = 25'b0000101010101000010101111;
    rom[30317] = 25'b0000101010110010101000000;
    rom[30318] = 25'b0000101010111100111010101;
    rom[30319] = 25'b0000101011000111001101100;
    rom[30320] = 25'b0000101011010001100000110;
    rom[30321] = 25'b0000101011011011110100011;
    rom[30322] = 25'b0000101011100110001000010;
    rom[30323] = 25'b0000101011110000011100100;
    rom[30324] = 25'b0000101011111010110001001;
    rom[30325] = 25'b0000101100000101000110000;
    rom[30326] = 25'b0000101100001111011011010;
    rom[30327] = 25'b0000101100011001110000111;
    rom[30328] = 25'b0000101100100100000110111;
    rom[30329] = 25'b0000101100101110011101001;
    rom[30330] = 25'b0000101100111000110011111;
    rom[30331] = 25'b0000101101000011001010110;
    rom[30332] = 25'b0000101101001101100010000;
    rom[30333] = 25'b0000101101010111111001101;
    rom[30334] = 25'b0000101101100010010001101;
    rom[30335] = 25'b0000101101101100101010000;
    rom[30336] = 25'b0000101101110111000010101;
    rom[30337] = 25'b0000101110000001011011100;
    rom[30338] = 25'b0000101110001011110100110;
    rom[30339] = 25'b0000101110010110001110100;
    rom[30340] = 25'b0000101110100000101000011;
    rom[30341] = 25'b0000101110101011000010110;
    rom[30342] = 25'b0000101110110101011101011;
    rom[30343] = 25'b0000101110111111111000010;
    rom[30344] = 25'b0000101111001010010011101;
    rom[30345] = 25'b0000101111010100101111010;
    rom[30346] = 25'b0000101111011111001011001;
    rom[30347] = 25'b0000101111101001100111100;
    rom[30348] = 25'b0000101111110100000100001;
    rom[30349] = 25'b0000101111111110100001000;
    rom[30350] = 25'b0000110000001000111110011;
    rom[30351] = 25'b0000110000010011011011111;
    rom[30352] = 25'b0000110000011101111001111;
    rom[30353] = 25'b0000110000101000011000001;
    rom[30354] = 25'b0000110000110010110110110;
    rom[30355] = 25'b0000110000111101010101101;
    rom[30356] = 25'b0000110001000111110100111;
    rom[30357] = 25'b0000110001010010010100011;
    rom[30358] = 25'b0000110001011100110100011;
    rom[30359] = 25'b0000110001100111010100100;
    rom[30360] = 25'b0000110001110001110101001;
    rom[30361] = 25'b0000110001111100010110000;
    rom[30362] = 25'b0000110010000110110111001;
    rom[30363] = 25'b0000110010010001011000101;
    rom[30364] = 25'b0000110010011011111010100;
    rom[30365] = 25'b0000110010100110011100101;
    rom[30366] = 25'b0000110010110000111111001;
    rom[30367] = 25'b0000110010111011100001111;
    rom[30368] = 25'b0000110011000110000101000;
    rom[30369] = 25'b0000110011010000101000100;
    rom[30370] = 25'b0000110011011011001100010;
    rom[30371] = 25'b0000110011100101110000011;
    rom[30372] = 25'b0000110011110000010100110;
    rom[30373] = 25'b0000110011111010111001100;
    rom[30374] = 25'b0000110100000101011110100;
    rom[30375] = 25'b0000110100010000000011111;
    rom[30376] = 25'b0000110100011010101001101;
    rom[30377] = 25'b0000110100100101001111101;
    rom[30378] = 25'b0000110100101111110101111;
    rom[30379] = 25'b0000110100111010011100100;
    rom[30380] = 25'b0000110101000101000011100;
    rom[30381] = 25'b0000110101001111101010110;
    rom[30382] = 25'b0000110101011010010010011;
    rom[30383] = 25'b0000110101100100111010010;
    rom[30384] = 25'b0000110101101111100010011;
    rom[30385] = 25'b0000110101111010001011000;
    rom[30386] = 25'b0000110110000100110011111;
    rom[30387] = 25'b0000110110001111011101000;
    rom[30388] = 25'b0000110110011010000110011;
    rom[30389] = 25'b0000110110100100110000010;
    rom[30390] = 25'b0000110110101111011010011;
    rom[30391] = 25'b0000110110111010000100110;
    rom[30392] = 25'b0000110111000100101111100;
    rom[30393] = 25'b0000110111001111011010100;
    rom[30394] = 25'b0000110111011010000101111;
    rom[30395] = 25'b0000110111100100110001100;
    rom[30396] = 25'b0000110111101111011101100;
    rom[30397] = 25'b0000110111111010001001110;
    rom[30398] = 25'b0000111000000100110110011;
    rom[30399] = 25'b0000111000001111100011010;
    rom[30400] = 25'b0000111000011010010000011;
    rom[30401] = 25'b0000111000100100111101111;
    rom[30402] = 25'b0000111000101111101011110;
    rom[30403] = 25'b0000111000111010011001111;
    rom[30404] = 25'b0000111001000101001000010;
    rom[30405] = 25'b0000111001001111110111000;
    rom[30406] = 25'b0000111001011010100110000;
    rom[30407] = 25'b0000111001100101010101011;
    rom[30408] = 25'b0000111001110000000101001;
    rom[30409] = 25'b0000111001111010110101000;
    rom[30410] = 25'b0000111010000101100101010;
    rom[30411] = 25'b0000111010010000010101110;
    rom[30412] = 25'b0000111010011011000110101;
    rom[30413] = 25'b0000111010100101110111111;
    rom[30414] = 25'b0000111010110000101001010;
    rom[30415] = 25'b0000111010111011011011001;
    rom[30416] = 25'b0000111011000110001101001;
    rom[30417] = 25'b0000111011010000111111100;
    rom[30418] = 25'b0000111011011011110010001;
    rom[30419] = 25'b0000111011100110100101010;
    rom[30420] = 25'b0000111011110001011000100;
    rom[30421] = 25'b0000111011111100001100000;
    rom[30422] = 25'b0000111100000110111111111;
    rom[30423] = 25'b0000111100010001110100001;
    rom[30424] = 25'b0000111100011100101000100;
    rom[30425] = 25'b0000111100100111011101010;
    rom[30426] = 25'b0000111100110010010010011;
    rom[30427] = 25'b0000111100111101000111110;
    rom[30428] = 25'b0000111101000111111101011;
    rom[30429] = 25'b0000111101010010110011011;
    rom[30430] = 25'b0000111101011101101001101;
    rom[30431] = 25'b0000111101101000100000001;
    rom[30432] = 25'b0000111101110011010111000;
    rom[30433] = 25'b0000111101111110001110001;
    rom[30434] = 25'b0000111110001001000101100;
    rom[30435] = 25'b0000111110010011111101010;
    rom[30436] = 25'b0000111110011110110101010;
    rom[30437] = 25'b0000111110101001101101101;
    rom[30438] = 25'b0000111110110100100110001;
    rom[30439] = 25'b0000111110111111011111001;
    rom[30440] = 25'b0000111111001010011000010;
    rom[30441] = 25'b0000111111010101010001110;
    rom[30442] = 25'b0000111111100000001011100;
    rom[30443] = 25'b0000111111101011000101100;
    rom[30444] = 25'b0000111111110101111111111;
    rom[30445] = 25'b0001000000000000111010100;
    rom[30446] = 25'b0001000000001011110101011;
    rom[30447] = 25'b0001000000010110110000101;
    rom[30448] = 25'b0001000000100001101100001;
    rom[30449] = 25'b0001000000101100100111111;
    rom[30450] = 25'b0001000000110111100100000;
    rom[30451] = 25'b0001000001000010100000011;
    rom[30452] = 25'b0001000001001101011101000;
    rom[30453] = 25'b0001000001011000011001111;
    rom[30454] = 25'b0001000001100011010111001;
    rom[30455] = 25'b0001000001101110010100101;
    rom[30456] = 25'b0001000001111001010010011;
    rom[30457] = 25'b0001000010000100010000011;
    rom[30458] = 25'b0001000010001111001110110;
    rom[30459] = 25'b0001000010011010001101100;
    rom[30460] = 25'b0001000010100101001100011;
    rom[30461] = 25'b0001000010110000001011101;
    rom[30462] = 25'b0001000010111011001011000;
    rom[30463] = 25'b0001000011000110001010111;
    rom[30464] = 25'b0001000011010001001010110;
    rom[30465] = 25'b0001000011011100001011001;
    rom[30466] = 25'b0001000011100111001011110;
    rom[30467] = 25'b0001000011110010001100101;
    rom[30468] = 25'b0001000011111101001101110;
    rom[30469] = 25'b0001000100001000001111010;
    rom[30470] = 25'b0001000100010011010000111;
    rom[30471] = 25'b0001000100011110010010111;
    rom[30472] = 25'b0001000100101001010101001;
    rom[30473] = 25'b0001000100110100010111110;
    rom[30474] = 25'b0001000100111111011010100;
    rom[30475] = 25'b0001000101001010011101101;
    rom[30476] = 25'b0001000101010101100001000;
    rom[30477] = 25'b0001000101100000100100101;
    rom[30478] = 25'b0001000101101011101000100;
    rom[30479] = 25'b0001000101110110101100110;
    rom[30480] = 25'b0001000110000001110001010;
    rom[30481] = 25'b0001000110001100110101111;
    rom[30482] = 25'b0001000110010111111010111;
    rom[30483] = 25'b0001000110100011000000010;
    rom[30484] = 25'b0001000110101110000101111;
    rom[30485] = 25'b0001000110111001001011101;
    rom[30486] = 25'b0001000111000100010001110;
    rom[30487] = 25'b0001000111001111011000001;
    rom[30488] = 25'b0001000111011010011110110;
    rom[30489] = 25'b0001000111100101100101101;
    rom[30490] = 25'b0001000111110000101100110;
    rom[30491] = 25'b0001000111111011110100010;
    rom[30492] = 25'b0001001000000110111100000;
    rom[30493] = 25'b0001001000010010000100000;
    rom[30494] = 25'b0001001000011101001100010;
    rom[30495] = 25'b0001001000101000010100110;
    rom[30496] = 25'b0001001000110011011101100;
    rom[30497] = 25'b0001001000111110100110100;
    rom[30498] = 25'b0001001001001001101111111;
    rom[30499] = 25'b0001001001010100111001011;
    rom[30500] = 25'b0001001001100000000011010;
    rom[30501] = 25'b0001001001101011001101011;
    rom[30502] = 25'b0001001001110110010111110;
    rom[30503] = 25'b0001001010000001100010011;
    rom[30504] = 25'b0001001010001100101101010;
    rom[30505] = 25'b0001001010010111111000011;
    rom[30506] = 25'b0001001010100011000011111;
    rom[30507] = 25'b0001001010101110001111100;
    rom[30508] = 25'b0001001010111001011011100;
    rom[30509] = 25'b0001001011000100100111101;
    rom[30510] = 25'b0001001011001111110100001;
    rom[30511] = 25'b0001001011011011000000111;
    rom[30512] = 25'b0001001011100110001101110;
    rom[30513] = 25'b0001001011110001011011000;
    rom[30514] = 25'b0001001011111100101000100;
    rom[30515] = 25'b0001001100000111110110010;
    rom[30516] = 25'b0001001100010011000100011;
    rom[30517] = 25'b0001001100011110010010101;
    rom[30518] = 25'b0001001100101001100001001;
    rom[30519] = 25'b0001001100110100101111111;
    rom[30520] = 25'b0001001100111111111110111;
    rom[30521] = 25'b0001001101001011001110001;
    rom[30522] = 25'b0001001101010110011101101;
    rom[30523] = 25'b0001001101100001101101100;
    rom[30524] = 25'b0001001101101100111101100;
    rom[30525] = 25'b0001001101111000001101111;
    rom[30526] = 25'b0001001110000011011110011;
    rom[30527] = 25'b0001001110001110101111001;
    rom[30528] = 25'b0001001110011010000000010;
    rom[30529] = 25'b0001001110100101010001100;
    rom[30530] = 25'b0001001110110000100011001;
    rom[30531] = 25'b0001001110111011110100111;
    rom[30532] = 25'b0001001111000111000111000;
    rom[30533] = 25'b0001001111010010011001010;
    rom[30534] = 25'b0001001111011101101011111;
    rom[30535] = 25'b0001001111101000111110101;
    rom[30536] = 25'b0001001111110100010001101;
    rom[30537] = 25'b0001001111111111100101000;
    rom[30538] = 25'b0001010000001010111000100;
    rom[30539] = 25'b0001010000010110001100010;
    rom[30540] = 25'b0001010000100001100000010;
    rom[30541] = 25'b0001010000101100110100101;
    rom[30542] = 25'b0001010000111000001001001;
    rom[30543] = 25'b0001010001000011011101111;
    rom[30544] = 25'b0001010001001110110011000;
    rom[30545] = 25'b0001010001011010001000001;
    rom[30546] = 25'b0001010001100101011101110;
    rom[30547] = 25'b0001010001110000110011011;
    rom[30548] = 25'b0001010001111100001001011;
    rom[30549] = 25'b0001010010000111011111101;
    rom[30550] = 25'b0001010010010010110110000;
    rom[30551] = 25'b0001010010011110001100110;
    rom[30552] = 25'b0001010010101001100011110;
    rom[30553] = 25'b0001010010110100111010111;
    rom[30554] = 25'b0001010011000000010010011;
    rom[30555] = 25'b0001010011001011101010000;
    rom[30556] = 25'b0001010011010111000001111;
    rom[30557] = 25'b0001010011100010011010001;
    rom[30558] = 25'b0001010011101101110010011;
    rom[30559] = 25'b0001010011111001001011001;
    rom[30560] = 25'b0001010100000100100011111;
    rom[30561] = 25'b0001010100001111111101000;
    rom[30562] = 25'b0001010100011011010110010;
    rom[30563] = 25'b0001010100100110101111111;
    rom[30564] = 25'b0001010100110010001001101;
    rom[30565] = 25'b0001010100111101100011101;
    rom[30566] = 25'b0001010101001000111110000;
    rom[30567] = 25'b0001010101010100011000011;
    rom[30568] = 25'b0001010101011111110011010;
    rom[30569] = 25'b0001010101101011001110001;
    rom[30570] = 25'b0001010101110110101001010;
    rom[30571] = 25'b0001010110000010000100110;
    rom[30572] = 25'b0001010110001101100000011;
    rom[30573] = 25'b0001010110011000111100010;
    rom[30574] = 25'b0001010110100100011000011;
    rom[30575] = 25'b0001010110101111110100110;
    rom[30576] = 25'b0001010110111011010001010;
    rom[30577] = 25'b0001010111000110101110000;
    rom[30578] = 25'b0001010111010010001011000;
    rom[30579] = 25'b0001010111011101101000011;
    rom[30580] = 25'b0001010111101001000101110;
    rom[30581] = 25'b0001010111110100100011011;
    rom[30582] = 25'b0001011000000000000001011;
    rom[30583] = 25'b0001011000001011011111101;
    rom[30584] = 25'b0001011000010110111110000;
    rom[30585] = 25'b0001011000100010011100100;
    rom[30586] = 25'b0001011000101101111011011;
    rom[30587] = 25'b0001011000111001011010011;
    rom[30588] = 25'b0001011001000100111001110;
    rom[30589] = 25'b0001011001010000011001010;
    rom[30590] = 25'b0001011001011011111000111;
    rom[30591] = 25'b0001011001100111011000110;
    rom[30592] = 25'b0001011001110010111001000;
    rom[30593] = 25'b0001011001111110011001011;
    rom[30594] = 25'b0001011010001001111010000;
    rom[30595] = 25'b0001011010010101011010110;
    rom[30596] = 25'b0001011010100000111011110;
    rom[30597] = 25'b0001011010101100011101000;
    rom[30598] = 25'b0001011010110111111110100;
    rom[30599] = 25'b0001011011000011100000010;
    rom[30600] = 25'b0001011011001111000010001;
    rom[30601] = 25'b0001011011011010100100010;
    rom[30602] = 25'b0001011011100110000110100;
    rom[30603] = 25'b0001011011110001101001001;
    rom[30604] = 25'b0001011011111101001011111;
    rom[30605] = 25'b0001011100001000101110111;
    rom[30606] = 25'b0001011100010100010010000;
    rom[30607] = 25'b0001011100011111110101100;
    rom[30608] = 25'b0001011100101011011001001;
    rom[30609] = 25'b0001011100110110111100111;
    rom[30610] = 25'b0001011101000010100001000;
    rom[30611] = 25'b0001011101001110000101010;
    rom[30612] = 25'b0001011101011001101001101;
    rom[30613] = 25'b0001011101100101001110011;
    rom[30614] = 25'b0001011101110000110011010;
    rom[30615] = 25'b0001011101111100011000011;
    rom[30616] = 25'b0001011110000111111101101;
    rom[30617] = 25'b0001011110010011100011001;
    rom[30618] = 25'b0001011110011111001001000;
    rom[30619] = 25'b0001011110101010101110110;
    rom[30620] = 25'b0001011110110110010101000;
    rom[30621] = 25'b0001011111000001111011010;
    rom[30622] = 25'b0001011111001101100001111;
    rom[30623] = 25'b0001011111011001001000101;
    rom[30624] = 25'b0001011111100100101111101;
    rom[30625] = 25'b0001011111110000010110110;
    rom[30626] = 25'b0001011111111011111110001;
    rom[30627] = 25'b0001100000000111100101101;
    rom[30628] = 25'b0001100000010011001101100;
    rom[30629] = 25'b0001100000011110110101011;
    rom[30630] = 25'b0001100000101010011101101;
    rom[30631] = 25'b0001100000110110000110000;
    rom[30632] = 25'b0001100001000001101110101;
    rom[30633] = 25'b0001100001001101010111011;
    rom[30634] = 25'b0001100001011001000000011;
    rom[30635] = 25'b0001100001100100101001100;
    rom[30636] = 25'b0001100001110000010011000;
    rom[30637] = 25'b0001100001111011111100100;
    rom[30638] = 25'b0001100010000111100110011;
    rom[30639] = 25'b0001100010010011010000010;
    rom[30640] = 25'b0001100010011110111010100;
    rom[30641] = 25'b0001100010101010100100111;
    rom[30642] = 25'b0001100010110110001111011;
    rom[30643] = 25'b0001100011000001111010001;
    rom[30644] = 25'b0001100011001101100101001;
    rom[30645] = 25'b0001100011011001010000010;
    rom[30646] = 25'b0001100011100100111011101;
    rom[30647] = 25'b0001100011110000100111001;
    rom[30648] = 25'b0001100011111100010010111;
    rom[30649] = 25'b0001100100000111111110110;
    rom[30650] = 25'b0001100100010011101010111;
    rom[30651] = 25'b0001100100011111010111010;
    rom[30652] = 25'b0001100100101011000011110;
    rom[30653] = 25'b0001100100110110110000011;
    rom[30654] = 25'b0001100101000010011101010;
    rom[30655] = 25'b0001100101001110001010011;
    rom[30656] = 25'b0001100101011001110111101;
    rom[30657] = 25'b0001100101100101100101000;
    rom[30658] = 25'b0001100101110001010010110;
    rom[30659] = 25'b0001100101111101000000100;
    rom[30660] = 25'b0001100110001000101110100;
    rom[30661] = 25'b0001100110010100011100110;
    rom[30662] = 25'b0001100110100000001011001;
    rom[30663] = 25'b0001100110101011111001101;
    rom[30664] = 25'b0001100110110111101000100;
    rom[30665] = 25'b0001100111000011010111011;
    rom[30666] = 25'b0001100111001111000110100;
    rom[30667] = 25'b0001100111011010110101110;
    rom[30668] = 25'b0001100111100110100101010;
    rom[30669] = 25'b0001100111110010010101000;
    rom[30670] = 25'b0001100111111110000100110;
    rom[30671] = 25'b0001101000001001110100110;
    rom[30672] = 25'b0001101000010101100101000;
    rom[30673] = 25'b0001101000100001010101011;
    rom[30674] = 25'b0001101000101101000101111;
    rom[30675] = 25'b0001101000111000110110110;
    rom[30676] = 25'b0001101001000100100111101;
    rom[30677] = 25'b0001101001010000011000110;
    rom[30678] = 25'b0001101001011100001010000;
    rom[30679] = 25'b0001101001100111111011100;
    rom[30680] = 25'b0001101001110011101101001;
    rom[30681] = 25'b0001101001111111011110111;
    rom[30682] = 25'b0001101010001011010000111;
    rom[30683] = 25'b0001101010010111000011001;
    rom[30684] = 25'b0001101010100010110101011;
    rom[30685] = 25'b0001101010101110101000000;
    rom[30686] = 25'b0001101010111010011010101;
    rom[30687] = 25'b0001101011000110001101100;
    rom[30688] = 25'b0001101011010010000000100;
    rom[30689] = 25'b0001101011011101110011110;
    rom[30690] = 25'b0001101011101001100111000;
    rom[30691] = 25'b0001101011110101011010101;
    rom[30692] = 25'b0001101100000001001110011;
    rom[30693] = 25'b0001101100001101000010010;
    rom[30694] = 25'b0001101100011000110110010;
    rom[30695] = 25'b0001101100100100101010100;
    rom[30696] = 25'b0001101100110000011111000;
    rom[30697] = 25'b0001101100111100010011100;
    rom[30698] = 25'b0001101101001000001000010;
    rom[30699] = 25'b0001101101010011111101001;
    rom[30700] = 25'b0001101101011111110010010;
    rom[30701] = 25'b0001101101101011100111011;
    rom[30702] = 25'b0001101101110111011100111;
    rom[30703] = 25'b0001101110000011010010011;
    rom[30704] = 25'b0001101110001111001000000;
    rom[30705] = 25'b0001101110011010111110000;
    rom[30706] = 25'b0001101110100110110100000;
    rom[30707] = 25'b0001101110110010101010010;
    rom[30708] = 25'b0001101110111110100000101;
    rom[30709] = 25'b0001101111001010010111001;
    rom[30710] = 25'b0001101111010110001101111;
    rom[30711] = 25'b0001101111100010000100110;
    rom[30712] = 25'b0001101111101101111011101;
    rom[30713] = 25'b0001101111111001110010111;
    rom[30714] = 25'b0001110000000101101010010;
    rom[30715] = 25'b0001110000010001100001110;
    rom[30716] = 25'b0001110000011101011001011;
    rom[30717] = 25'b0001110000101001010001001;
    rom[30718] = 25'b0001110000110101001001001;
    rom[30719] = 25'b0001110001000001000001010;
    rom[30720] = 25'b0001110001001100111001101;
    rom[30721] = 25'b0001110001011000110010000;
    rom[30722] = 25'b0001110001100100101010101;
    rom[30723] = 25'b0001110001110000100011010;
    rom[30724] = 25'b0001110001111100011100010;
    rom[30725] = 25'b0001110010001000010101010;
    rom[30726] = 25'b0001110010010100001110011;
    rom[30727] = 25'b0001110010100000000111111;
    rom[30728] = 25'b0001110010101100000001010;
    rom[30729] = 25'b0001110010110111111011000;
    rom[30730] = 25'b0001110011000011110100110;
    rom[30731] = 25'b0001110011001111101110110;
    rom[30732] = 25'b0001110011011011101000111;
    rom[30733] = 25'b0001110011100111100011001;
    rom[30734] = 25'b0001110011110011011101100;
    rom[30735] = 25'b0001110011111111011000000;
    rom[30736] = 25'b0001110100001011010010110;
    rom[30737] = 25'b0001110100010111001101101;
    rom[30738] = 25'b0001110100100011001000101;
    rom[30739] = 25'b0001110100101111000011110;
    rom[30740] = 25'b0001110100111010111111001;
    rom[30741] = 25'b0001110101000110111010011;
    rom[30742] = 25'b0001110101010010110110000;
    rom[30743] = 25'b0001110101011110110001110;
    rom[30744] = 25'b0001110101101010101101101;
    rom[30745] = 25'b0001110101110110101001101;
    rom[30746] = 25'b0001110110000010100101110;
    rom[30747] = 25'b0001110110001110100010000;
    rom[30748] = 25'b0001110110011010011110100;
    rom[30749] = 25'b0001110110100110011011001;
    rom[30750] = 25'b0001110110110010010111110;
    rom[30751] = 25'b0001110110111110010100100;
    rom[30752] = 25'b0001110111001010010001101;
    rom[30753] = 25'b0001110111010110001110110;
    rom[30754] = 25'b0001110111100010001100000;
    rom[30755] = 25'b0001110111101110001001011;
    rom[30756] = 25'b0001110111111010000110111;
    rom[30757] = 25'b0001111000000110000100101;
    rom[30758] = 25'b0001111000010010000010011;
    rom[30759] = 25'b0001111000011110000000011;
    rom[30760] = 25'b0001111000101001111110100;
    rom[30761] = 25'b0001111000110101111100101;
    rom[30762] = 25'b0001111001000001111011000;
    rom[30763] = 25'b0001111001001101111001100;
    rom[30764] = 25'b0001111001011001111000001;
    rom[30765] = 25'b0001111001100101110110110;
    rom[30766] = 25'b0001111001110001110101101;
    rom[30767] = 25'b0001111001111101110100101;
    rom[30768] = 25'b0001111010001001110011111;
    rom[30769] = 25'b0001111010010101110011001;
    rom[30770] = 25'b0001111010100001110010100;
    rom[30771] = 25'b0001111010101101110010000;
    rom[30772] = 25'b0001111010111001110001101;
    rom[30773] = 25'b0001111011000101110001100;
    rom[30774] = 25'b0001111011010001110001011;
    rom[30775] = 25'b0001111011011101110001011;
    rom[30776] = 25'b0001111011101001110001100;
    rom[30777] = 25'b0001111011110101110001111;
    rom[30778] = 25'b0001111100000001110010011;
    rom[30779] = 25'b0001111100001101110010110;
    rom[30780] = 25'b0001111100011001110011100;
    rom[30781] = 25'b0001111100100101110100010;
    rom[30782] = 25'b0001111100110001110101001;
    rom[30783] = 25'b0001111100111101110110010;
    rom[30784] = 25'b0001111101001001110111011;
    rom[30785] = 25'b0001111101010101111000101;
    rom[30786] = 25'b0001111101100001111010000;
    rom[30787] = 25'b0001111101101101111011100;
    rom[30788] = 25'b0001111101111001111101001;
    rom[30789] = 25'b0001111110000101111110111;
    rom[30790] = 25'b0001111110010010000000110;
    rom[30791] = 25'b0001111110011110000010110;
    rom[30792] = 25'b0001111110101010000100111;
    rom[30793] = 25'b0001111110110110000111001;
    rom[30794] = 25'b0001111111000010001001011;
    rom[30795] = 25'b0001111111001110001011111;
    rom[30796] = 25'b0001111111011010001110011;
    rom[30797] = 25'b0001111111100110010001001;
    rom[30798] = 25'b0001111111110010010100000;
    rom[30799] = 25'b0001111111111110010110111;
    rom[30800] = 25'b0010000000001010011001111;
    rom[30801] = 25'b0010000000010110011101000;
    rom[30802] = 25'b0010000000100010100000010;
    rom[30803] = 25'b0010000000101110100011101;
    rom[30804] = 25'b0010000000111010100111001;
    rom[30805] = 25'b0010000001000110101010101;
    rom[30806] = 25'b0010000001010010101110011;
    rom[30807] = 25'b0010000001011110110010001;
    rom[30808] = 25'b0010000001101010110110001;
    rom[30809] = 25'b0010000001110110111010001;
    rom[30810] = 25'b0010000010000010111110010;
    rom[30811] = 25'b0010000010001111000010100;
    rom[30812] = 25'b0010000010011011000110110;
    rom[30813] = 25'b0010000010100111001011010;
    rom[30814] = 25'b0010000010110011001111110;
    rom[30815] = 25'b0010000010111111010100100;
    rom[30816] = 25'b0010000011001011011001010;
    rom[30817] = 25'b0010000011010111011110001;
    rom[30818] = 25'b0010000011100011100011001;
    rom[30819] = 25'b0010000011101111101000001;
    rom[30820] = 25'b0010000011111011101101010;
    rom[30821] = 25'b0010000100000111110010100;
    rom[30822] = 25'b0010000100010011111000000;
    rom[30823] = 25'b0010000100011111111101011;
    rom[30824] = 25'b0010000100101100000011000;
    rom[30825] = 25'b0010000100111000001000101;
    rom[30826] = 25'b0010000101000100001110011;
    rom[30827] = 25'b0010000101010000010100011;
    rom[30828] = 25'b0010000101011100011010010;
    rom[30829] = 25'b0010000101101000100000010;
    rom[30830] = 25'b0010000101110100100110100;
    rom[30831] = 25'b0010000110000000101100110;
    rom[30832] = 25'b0010000110001100110011001;
    rom[30833] = 25'b0010000110011000111001101;
    rom[30834] = 25'b0010000110100101000000001;
    rom[30835] = 25'b0010000110110001000110110;
    rom[30836] = 25'b0010000110111101001101100;
    rom[30837] = 25'b0010000111001001010100010;
    rom[30838] = 25'b0010000111010101011011001;
    rom[30839] = 25'b0010000111100001100010010;
    rom[30840] = 25'b0010000111101101101001010;
    rom[30841] = 25'b0010000111111001110000100;
    rom[30842] = 25'b0010001000000101110111111;
    rom[30843] = 25'b0010001000010001111111001;
    rom[30844] = 25'b0010001000011110000110101;
    rom[30845] = 25'b0010001000101010001110001;
    rom[30846] = 25'b0010001000110110010101110;
    rom[30847] = 25'b0010001001000010011101100;
    rom[30848] = 25'b0010001001001110100101010;
    rom[30849] = 25'b0010001001011010101101010;
    rom[30850] = 25'b0010001001100110110101010;
    rom[30851] = 25'b0010001001110010111101010;
    rom[30852] = 25'b0010001001111111000101011;
    rom[30853] = 25'b0010001010001011001101101;
    rom[30854] = 25'b0010001010010111010110000;
    rom[30855] = 25'b0010001010100011011110011;
    rom[30856] = 25'b0010001010101111100110111;
    rom[30857] = 25'b0010001010111011101111011;
    rom[30858] = 25'b0010001011000111111000001;
    rom[30859] = 25'b0010001011010100000000110;
    rom[30860] = 25'b0010001011100000001001101;
    rom[30861] = 25'b0010001011101100010010100;
    rom[30862] = 25'b0010001011111000011011100;
    rom[30863] = 25'b0010001100000100100100100;
    rom[30864] = 25'b0010001100010000101101101;
    rom[30865] = 25'b0010001100011100110110111;
    rom[30866] = 25'b0010001100101001000000001;
    rom[30867] = 25'b0010001100110101001001100;
    rom[30868] = 25'b0010001101000001010010111;
    rom[30869] = 25'b0010001101001101011100011;
    rom[30870] = 25'b0010001101011001100110000;
    rom[30871] = 25'b0010001101100101101111101;
    rom[30872] = 25'b0010001101110001111001011;
    rom[30873] = 25'b0010001101111110000011001;
    rom[30874] = 25'b0010001110001010001101000;
    rom[30875] = 25'b0010001110010110010110111;
    rom[30876] = 25'b0010001110100010100000111;
    rom[30877] = 25'b0010001110101110101011000;
    rom[30878] = 25'b0010001110111010110101010;
    rom[30879] = 25'b0010001111000110111111011;
    rom[30880] = 25'b0010001111010011001001110;
    rom[30881] = 25'b0010001111011111010100001;
    rom[30882] = 25'b0010001111101011011110100;
    rom[30883] = 25'b0010001111110111101001000;
    rom[30884] = 25'b0010010000000011110011101;
    rom[30885] = 25'b0010010000001111111110001;
    rom[30886] = 25'b0010010000011100001000111;
    rom[30887] = 25'b0010010000101000010011101;
    rom[30888] = 25'b0010010000110100011110011;
    rom[30889] = 25'b0010010001000000101001011;
    rom[30890] = 25'b0010010001001100110100010;
    rom[30891] = 25'b0010010001011000111111011;
    rom[30892] = 25'b0010010001100101001010011;
    rom[30893] = 25'b0010010001110001010101100;
    rom[30894] = 25'b0010010001111101100000110;
    rom[30895] = 25'b0010010010001001101100000;
    rom[30896] = 25'b0010010010010101110111010;
    rom[30897] = 25'b0010010010100010000010101;
    rom[30898] = 25'b0010010010101110001110001;
    rom[30899] = 25'b0010010010111010011001101;
    rom[30900] = 25'b0010010011000110100101001;
    rom[30901] = 25'b0010010011010010110000110;
    rom[30902] = 25'b0010010011011110111100100;
    rom[30903] = 25'b0010010011101011001000001;
    rom[30904] = 25'b0010010011110111010011111;
    rom[30905] = 25'b0010010100000011011111110;
    rom[30906] = 25'b0010010100001111101011101;
    rom[30907] = 25'b0010010100011011110111100;
    rom[30908] = 25'b0010010100101000000011101;
    rom[30909] = 25'b0010010100110100001111101;
    rom[30910] = 25'b0010010101000000011011110;
    rom[30911] = 25'b0010010101001100100111111;
    rom[30912] = 25'b0010010101011000110100000;
    rom[30913] = 25'b0010010101100101000000010;
    rom[30914] = 25'b0010010101110001001100101;
    rom[30915] = 25'b0010010101111101011001000;
    rom[30916] = 25'b0010010110001001100101011;
    rom[30917] = 25'b0010010110010101110001111;
    rom[30918] = 25'b0010010110100001111110010;
    rom[30919] = 25'b0010010110101110001010110;
    rom[30920] = 25'b0010010110111010010111011;
    rom[30921] = 25'b0010010111000110100100000;
    rom[30922] = 25'b0010010111010010110000110;
    rom[30923] = 25'b0010010111011110111101100;
    rom[30924] = 25'b0010010111101011001010010;
    rom[30925] = 25'b0010010111110111010111000;
    rom[30926] = 25'b0010011000000011100011111;
    rom[30927] = 25'b0010011000001111110000111;
    rom[30928] = 25'b0010011000011011111101110;
    rom[30929] = 25'b0010011000101000001010110;
    rom[30930] = 25'b0010011000110100010111110;
    rom[30931] = 25'b0010011001000000100100110;
    rom[30932] = 25'b0010011001001100110001111;
    rom[30933] = 25'b0010011001011000111111001;
    rom[30934] = 25'b0010011001100101001100001;
    rom[30935] = 25'b0010011001110001011001011;
    rom[30936] = 25'b0010011001111101100110110;
    rom[30937] = 25'b0010011010001001110100000;
    rom[30938] = 25'b0010011010010110000001010;
    rom[30939] = 25'b0010011010100010001110101;
    rom[30940] = 25'b0010011010101110011100000;
    rom[30941] = 25'b0010011010111010101001100;
    rom[30942] = 25'b0010011011000110110110111;
    rom[30943] = 25'b0010011011010011000100100;
    rom[30944] = 25'b0010011011011111010010000;
    rom[30945] = 25'b0010011011101011011111100;
    rom[30946] = 25'b0010011011110111101101001;
    rom[30947] = 25'b0010011100000011111010110;
    rom[30948] = 25'b0010011100010000001000100;
    rom[30949] = 25'b0010011100011100010110001;
    rom[30950] = 25'b0010011100101000100011111;
    rom[30951] = 25'b0010011100110100110001101;
    rom[30952] = 25'b0010011101000000111111011;
    rom[30953] = 25'b0010011101001101001101001;
    rom[30954] = 25'b0010011101011001011010111;
    rom[30955] = 25'b0010011101100101101000111;
    rom[30956] = 25'b0010011101110001110110101;
    rom[30957] = 25'b0010011101111110000100101;
    rom[30958] = 25'b0010011110001010010010100;
    rom[30959] = 25'b0010011110010110100000100;
    rom[30960] = 25'b0010011110100010101110100;
    rom[30961] = 25'b0010011110101110111100011;
    rom[30962] = 25'b0010011110111011001010011;
    rom[30963] = 25'b0010011111000111011000100;
    rom[30964] = 25'b0010011111010011100110101;
    rom[30965] = 25'b0010011111011111110100110;
    rom[30966] = 25'b0010011111101100000010110;
    rom[30967] = 25'b0010011111111000010000111;
    rom[30968] = 25'b0010100000000100011111000;
    rom[30969] = 25'b0010100000010000101101010;
    rom[30970] = 25'b0010100000011100111011011;
    rom[30971] = 25'b0010100000101001001001101;
    rom[30972] = 25'b0010100000110101010111110;
    rom[30973] = 25'b0010100001000001100110001;
    rom[30974] = 25'b0010100001001101110100010;
    rom[30975] = 25'b0010100001011010000010101;
    rom[30976] = 25'b0010100001100110010000110;
    rom[30977] = 25'b0010100001110010011111001;
    rom[30978] = 25'b0010100001111110101101011;
    rom[30979] = 25'b0010100010001010111011110;
    rom[30980] = 25'b0010100010010111001010001;
    rom[30981] = 25'b0010100010100011011000011;
    rom[30982] = 25'b0010100010101111100110110;
    rom[30983] = 25'b0010100010111011110101001;
    rom[30984] = 25'b0010100011001000000011100;
    rom[30985] = 25'b0010100011010100010001111;
    rom[30986] = 25'b0010100011100000100000010;
    rom[30987] = 25'b0010100011101100101110110;
    rom[30988] = 25'b0010100011111000111101001;
    rom[30989] = 25'b0010100100000101001011100;
    rom[30990] = 25'b0010100100010001011001111;
    rom[30991] = 25'b0010100100011101101000011;
    rom[30992] = 25'b0010100100101001110110110;
    rom[30993] = 25'b0010100100110110000101001;
    rom[30994] = 25'b0010100101000010010011101;
    rom[30995] = 25'b0010100101001110100010000;
    rom[30996] = 25'b0010100101011010110000100;
    rom[30997] = 25'b0010100101100110111111000;
    rom[30998] = 25'b0010100101110011001101011;
    rom[30999] = 25'b0010100101111111011011111;
    rom[31000] = 25'b0010100110001011101010011;
    rom[31001] = 25'b0010100110010111111000110;
    rom[31002] = 25'b0010100110100100000111010;
    rom[31003] = 25'b0010100110110000010101110;
    rom[31004] = 25'b0010100110111100100100001;
    rom[31005] = 25'b0010100111001000110010101;
    rom[31006] = 25'b0010100111010101000001001;
    rom[31007] = 25'b0010100111100001001111100;
    rom[31008] = 25'b0010100111101101011101111;
    rom[31009] = 25'b0010100111111001101100011;
    rom[31010] = 25'b0010101000000101111010110;
    rom[31011] = 25'b0010101000010010001001001;
    rom[31012] = 25'b0010101000011110010111101;
    rom[31013] = 25'b0010101000101010100110000;
    rom[31014] = 25'b0010101000110110110100011;
    rom[31015] = 25'b0010101001000011000010111;
    rom[31016] = 25'b0010101001001111010001010;
    rom[31017] = 25'b0010101001011011011111100;
    rom[31018] = 25'b0010101001100111101101111;
    rom[31019] = 25'b0010101001110011111100011;
    rom[31020] = 25'b0010101010000000001010101;
    rom[31021] = 25'b0010101010001100011000111;
    rom[31022] = 25'b0010101010011000100111010;
    rom[31023] = 25'b0010101010100100110101101;
    rom[31024] = 25'b0010101010110001000011111;
    rom[31025] = 25'b0010101010111101010010001;
    rom[31026] = 25'b0010101011001001100000100;
    rom[31027] = 25'b0010101011010101101110101;
    rom[31028] = 25'b0010101011100001111101000;
    rom[31029] = 25'b0010101011101110001011001;
    rom[31030] = 25'b0010101011111010011001011;
    rom[31031] = 25'b0010101100000110100111100;
    rom[31032] = 25'b0010101100010010110101110;
    rom[31033] = 25'b0010101100011111000011111;
    rom[31034] = 25'b0010101100101011010001111;
    rom[31035] = 25'b0010101100110111100000000;
    rom[31036] = 25'b0010101101000011101110001;
    rom[31037] = 25'b0010101101001111111100010;
    rom[31038] = 25'b0010101101011100001010010;
    rom[31039] = 25'b0010101101101000011000011;
    rom[31040] = 25'b0010101101110100100110011;
    rom[31041] = 25'b0010101110000000110100010;
    rom[31042] = 25'b0010101110001101000010010;
    rom[31043] = 25'b0010101110011001010000001;
    rom[31044] = 25'b0010101110100101011110001;
    rom[31045] = 25'b0010101110110001101100000;
    rom[31046] = 25'b0010101110111101111001111;
    rom[31047] = 25'b0010101111001010000111101;
    rom[31048] = 25'b0010101111010110010101100;
    rom[31049] = 25'b0010101111100010100011010;
    rom[31050] = 25'b0010101111101110110001000;
    rom[31051] = 25'b0010101111111010111110110;
    rom[31052] = 25'b0010110000000111001100011;
    rom[31053] = 25'b0010110000010011011010000;
    rom[31054] = 25'b0010110000011111100111101;
    rom[31055] = 25'b0010110000101011110101010;
    rom[31056] = 25'b0010110000111000000010110;
    rom[31057] = 25'b0010110001000100010000011;
    rom[31058] = 25'b0010110001010000011101111;
    rom[31059] = 25'b0010110001011100101011011;
    rom[31060] = 25'b0010110001101000111000110;
    rom[31061] = 25'b0010110001110101000110010;
    rom[31062] = 25'b0010110010000001010011100;
    rom[31063] = 25'b0010110010001101100000111;
    rom[31064] = 25'b0010110010011001101110001;
    rom[31065] = 25'b0010110010100101111011011;
    rom[31066] = 25'b0010110010110010001000101;
    rom[31067] = 25'b0010110010111110010101110;
    rom[31068] = 25'b0010110011001010100011000;
    rom[31069] = 25'b0010110011010110110000000;
    rom[31070] = 25'b0010110011100010111101000;
    rom[31071] = 25'b0010110011101111001010001;
    rom[31072] = 25'b0010110011111011010111000;
    rom[31073] = 25'b0010110100000111100100000;
    rom[31074] = 25'b0010110100010011110000111;
    rom[31075] = 25'b0010110100011111111101110;
    rom[31076] = 25'b0010110100101100001010100;
    rom[31077] = 25'b0010110100111000010111010;
    rom[31078] = 25'b0010110101000100100100000;
    rom[31079] = 25'b0010110101010000110000101;
    rom[31080] = 25'b0010110101011100111101010;
    rom[31081] = 25'b0010110101101001001001111;
    rom[31082] = 25'b0010110101110101010110100;
    rom[31083] = 25'b0010110110000001100010111;
    rom[31084] = 25'b0010110110001101101111011;
    rom[31085] = 25'b0010110110011001111011110;
    rom[31086] = 25'b0010110110100110001000001;
    rom[31087] = 25'b0010110110110010010100011;
    rom[31088] = 25'b0010110110111110100000101;
    rom[31089] = 25'b0010110111001010101100110;
    rom[31090] = 25'b0010110111010110111000111;
    rom[31091] = 25'b0010110111100011000101000;
    rom[31092] = 25'b0010110111101111010001000;
    rom[31093] = 25'b0010110111111011011101000;
    rom[31094] = 25'b0010111000000111101001000;
    rom[31095] = 25'b0010111000010011110100110;
    rom[31096] = 25'b0010111000100000000000101;
    rom[31097] = 25'b0010111000101100001100011;
    rom[31098] = 25'b0010111000111000011000001;
    rom[31099] = 25'b0010111001000100100011110;
    rom[31100] = 25'b0010111001010000101111010;
    rom[31101] = 25'b0010111001011100111010110;
    rom[31102] = 25'b0010111001101001000110010;
    rom[31103] = 25'b0010111001110101010001110;
    rom[31104] = 25'b0010111010000001011101000;
    rom[31105] = 25'b0010111010001101101000011;
    rom[31106] = 25'b0010111010011001110011100;
    rom[31107] = 25'b0010111010100101111110110;
    rom[31108] = 25'b0010111010110010001001110;
    rom[31109] = 25'b0010111010111110010100111;
    rom[31110] = 25'b0010111011001010011111111;
    rom[31111] = 25'b0010111011010110101010111;
    rom[31112] = 25'b0010111011100010110101101;
    rom[31113] = 25'b0010111011101111000000011;
    rom[31114] = 25'b0010111011111011001011001;
    rom[31115] = 25'b0010111100000111010101111;
    rom[31116] = 25'b0010111100010011100000011;
    rom[31117] = 25'b0010111100011111101010111;
    rom[31118] = 25'b0010111100101011110101011;
    rom[31119] = 25'b0010111100110111111111110;
    rom[31120] = 25'b0010111101000100001010000;
    rom[31121] = 25'b0010111101010000010100010;
    rom[31122] = 25'b0010111101011100011110100;
    rom[31123] = 25'b0010111101101000101000101;
    rom[31124] = 25'b0010111101110100110010101;
    rom[31125] = 25'b0010111110000000111100100;
    rom[31126] = 25'b0010111110001101000110011;
    rom[31127] = 25'b0010111110011001010000010;
    rom[31128] = 25'b0010111110100101011010000;
    rom[31129] = 25'b0010111110110001100011101;
    rom[31130] = 25'b0010111110111101101101010;
    rom[31131] = 25'b0010111111001001110110110;
    rom[31132] = 25'b0010111111010110000000001;
    rom[31133] = 25'b0010111111100010001001100;
    rom[31134] = 25'b0010111111101110010010111;
    rom[31135] = 25'b0010111111111010011100000;
    rom[31136] = 25'b0011000000000110100101001;
    rom[31137] = 25'b0011000000010010101110001;
    rom[31138] = 25'b0011000000011110110111001;
    rom[31139] = 25'b0011000000101011000000000;
    rom[31140] = 25'b0011000000110111001000111;
    rom[31141] = 25'b0011000001000011010001100;
    rom[31142] = 25'b0011000001001111011010010;
    rom[31143] = 25'b0011000001011011100010110;
    rom[31144] = 25'b0011000001100111101011010;
    rom[31145] = 25'b0011000001110011110011101;
    rom[31146] = 25'b0011000001111111111011111;
    rom[31147] = 25'b0011000010001100000100001;
    rom[31148] = 25'b0011000010011000001100010;
    rom[31149] = 25'b0011000010100100010100011;
    rom[31150] = 25'b0011000010110000011100010;
    rom[31151] = 25'b0011000010111100100100010;
    rom[31152] = 25'b0011000011001000101100000;
    rom[31153] = 25'b0011000011010100110011101;
    rom[31154] = 25'b0011000011100000111011010;
    rom[31155] = 25'b0011000011101101000010111;
    rom[31156] = 25'b0011000011111001001010010;
    rom[31157] = 25'b0011000100000101010001100;
    rom[31158] = 25'b0011000100010001011000111;
    rom[31159] = 25'b0011000100011101011111111;
    rom[31160] = 25'b0011000100101001100111000;
    rom[31161] = 25'b0011000100110101101110000;
    rom[31162] = 25'b0011000101000001110100111;
    rom[31163] = 25'b0011000101001101111011101;
    rom[31164] = 25'b0011000101011010000010011;
    rom[31165] = 25'b0011000101100110001000111;
    rom[31166] = 25'b0011000101110010001111011;
    rom[31167] = 25'b0011000101111110010101111;
    rom[31168] = 25'b0011000110001010011100001;
    rom[31169] = 25'b0011000110010110100010010;
    rom[31170] = 25'b0011000110100010101000011;
    rom[31171] = 25'b0011000110101110101110011;
    rom[31172] = 25'b0011000110111010110100011;
    rom[31173] = 25'b0011000111000110111010001;
    rom[31174] = 25'b0011000111010010111111110;
    rom[31175] = 25'b0011000111011111000101011;
    rom[31176] = 25'b0011000111101011001010111;
    rom[31177] = 25'b0011000111110111010000011;
    rom[31178] = 25'b0011001000000011010101101;
    rom[31179] = 25'b0011001000001111011010110;
    rom[31180] = 25'b0011001000011011011111111;
    rom[31181] = 25'b0011001000100111100100111;
    rom[31182] = 25'b0011001000110011101001110;
    rom[31183] = 25'b0011001000111111101110100;
    rom[31184] = 25'b0011001001001011110011001;
    rom[31185] = 25'b0011001001010111110111110;
    rom[31186] = 25'b0011001001100011111100001;
    rom[31187] = 25'b0011001001110000000000100;
    rom[31188] = 25'b0011001001111100000100110;
    rom[31189] = 25'b0011001010001000001000111;
    rom[31190] = 25'b0011001010010100001100110;
    rom[31191] = 25'b0011001010100000010000110;
    rom[31192] = 25'b0011001010101100010100100;
    rom[31193] = 25'b0011001010111000011000010;
    rom[31194] = 25'b0011001011000100011011101;
    rom[31195] = 25'b0011001011010000011111001;
    rom[31196] = 25'b0011001011011100100010100;
    rom[31197] = 25'b0011001011101000100101110;
    rom[31198] = 25'b0011001011110100101000111;
    rom[31199] = 25'b0011001100000000101011111;
    rom[31200] = 25'b0011001100001100101110101;
    rom[31201] = 25'b0011001100011000110001100;
    rom[31202] = 25'b0011001100100100110100001;
    rom[31203] = 25'b0011001100110000110110101;
    rom[31204] = 25'b0011001100111100111001000;
    rom[31205] = 25'b0011001101001000111011010;
    rom[31206] = 25'b0011001101010100111101011;
    rom[31207] = 25'b0011001101100000111111100;
    rom[31208] = 25'b0011001101101101000001011;
    rom[31209] = 25'b0011001101111001000011010;
    rom[31210] = 25'b0011001110000101000100111;
    rom[31211] = 25'b0011001110010001000110011;
    rom[31212] = 25'b0011001110011101000111111;
    rom[31213] = 25'b0011001110101001001001001;
    rom[31214] = 25'b0011001110110101001010010;
    rom[31215] = 25'b0011001111000001001011011;
    rom[31216] = 25'b0011001111001101001100010;
    rom[31217] = 25'b0011001111011001001101001;
    rom[31218] = 25'b0011001111100101001101111;
    rom[31219] = 25'b0011001111110001001110010;
    rom[31220] = 25'b0011001111111101001110110;
    rom[31221] = 25'b0011010000001001001111001;
    rom[31222] = 25'b0011010000010101001111001;
    rom[31223] = 25'b0011010000100001001111010;
    rom[31224] = 25'b0011010000101101001111001;
    rom[31225] = 25'b0011010000111001001111000;
    rom[31226] = 25'b0011010001000101001110101;
    rom[31227] = 25'b0011010001010001001110000;
    rom[31228] = 25'b0011010001011101001101011;
    rom[31229] = 25'b0011010001101001001100101;
    rom[31230] = 25'b0011010001110101001011110;
    rom[31231] = 25'b0011010010000001001010110;
    rom[31232] = 25'b0011010010001101001001101;
    rom[31233] = 25'b0011010010011001001000011;
    rom[31234] = 25'b0011010010100101000110111;
    rom[31235] = 25'b0011010010110001000101010;
    rom[31236] = 25'b0011010010111101000011101;
    rom[31237] = 25'b0011010011001001000001110;
    rom[31238] = 25'b0011010011010100111111110;
    rom[31239] = 25'b0011010011100000111101101;
    rom[31240] = 25'b0011010011101100111011011;
    rom[31241] = 25'b0011010011111000111001000;
    rom[31242] = 25'b0011010100000100110110100;
    rom[31243] = 25'b0011010100010000110011110;
    rom[31244] = 25'b0011010100011100110000111;
    rom[31245] = 25'b0011010100101000101101111;
    rom[31246] = 25'b0011010100110100101010111;
    rom[31247] = 25'b0011010101000000100111101;
    rom[31248] = 25'b0011010101001100100100001;
    rom[31249] = 25'b0011010101011000100000101;
    rom[31250] = 25'b0011010101100100011100111;
    rom[31251] = 25'b0011010101110000011001001;
    rom[31252] = 25'b0011010101111100010101001;
    rom[31253] = 25'b0011010110001000010001000;
    rom[31254] = 25'b0011010110010100001100110;
    rom[31255] = 25'b0011010110100000001000010;
    rom[31256] = 25'b0011010110101100000011101;
    rom[31257] = 25'b0011010110110111111110111;
    rom[31258] = 25'b0011010111000011111010001;
    rom[31259] = 25'b0011010111001111110101000;
    rom[31260] = 25'b0011010111011011101111111;
    rom[31261] = 25'b0011010111100111101010100;
    rom[31262] = 25'b0011010111110011100101000;
    rom[31263] = 25'b0011010111111111011111011;
    rom[31264] = 25'b0011011000001011011001101;
    rom[31265] = 25'b0011011000010111010011101;
    rom[31266] = 25'b0011011000100011001101100;
    rom[31267] = 25'b0011011000101111000111010;
    rom[31268] = 25'b0011011000111011000000111;
    rom[31269] = 25'b0011011001000110111010010;
    rom[31270] = 25'b0011011001010010110011101;
    rom[31271] = 25'b0011011001011110101100101;
    rom[31272] = 25'b0011011001101010100101101;
    rom[31273] = 25'b0011011001110110011110011;
    rom[31274] = 25'b0011011010000010010111000;
    rom[31275] = 25'b0011011010001110001111100;
    rom[31276] = 25'b0011011010011010000111111;
    rom[31277] = 25'b0011011010100101111111111;
    rom[31278] = 25'b0011011010110001110111111;
    rom[31279] = 25'b0011011010111101101111110;
    rom[31280] = 25'b0011011011001001100111011;
    rom[31281] = 25'b0011011011010101011110111;
    rom[31282] = 25'b0011011011100001010110010;
    rom[31283] = 25'b0011011011101101001101011;
    rom[31284] = 25'b0011011011111001000100100;
    rom[31285] = 25'b0011011100000100111011011;
    rom[31286] = 25'b0011011100010000110010000;
    rom[31287] = 25'b0011011100011100101000100;
    rom[31288] = 25'b0011011100101000011110110;
    rom[31289] = 25'b0011011100110100010101000;
    rom[31290] = 25'b0011011101000000001010111;
    rom[31291] = 25'b0011011101001100000000110;
    rom[31292] = 25'b0011011101010111110110011;
    rom[31293] = 25'b0011011101100011101100000;
    rom[31294] = 25'b0011011101101111100001010;
    rom[31295] = 25'b0011011101111011010110011;
    rom[31296] = 25'b0011011110000111001011011;
    rom[31297] = 25'b0011011110010011000000001;
    rom[31298] = 25'b0011011110011110110100110;
    rom[31299] = 25'b0011011110101010101001010;
    rom[31300] = 25'b0011011110110110011101100;
    rom[31301] = 25'b0011011111000010010001101;
    rom[31302] = 25'b0011011111001110000101100;
    rom[31303] = 25'b0011011111011001111001010;
    rom[31304] = 25'b0011011111100101101100111;
    rom[31305] = 25'b0011011111110001100000010;
    rom[31306] = 25'b0011011111111101010011100;
    rom[31307] = 25'b0011100000001001000110100;
    rom[31308] = 25'b0011100000010100111001011;
    rom[31309] = 25'b0011100000100000101100000;
    rom[31310] = 25'b0011100000101100011110100;
    rom[31311] = 25'b0011100000111000010000110;
    rom[31312] = 25'b0011100001000100000011000;
    rom[31313] = 25'b0011100001001111110100111;
    rom[31314] = 25'b0011100001011011100110101;
    rom[31315] = 25'b0011100001100111011000010;
    rom[31316] = 25'b0011100001110011001001101;
    rom[31317] = 25'b0011100001111110111010111;
    rom[31318] = 25'b0011100010001010101011111;
    rom[31319] = 25'b0011100010010110011100110;
    rom[31320] = 25'b0011100010100010001101011;
    rom[31321] = 25'b0011100010101101111101111;
    rom[31322] = 25'b0011100010111001101110001;
    rom[31323] = 25'b0011100011000101011110001;
    rom[31324] = 25'b0011100011010001001110001;
    rom[31325] = 25'b0011100011011100111101110;
    rom[31326] = 25'b0011100011101000101101011;
    rom[31327] = 25'b0011100011110100011100101;
    rom[31328] = 25'b0011100100000000001011110;
    rom[31329] = 25'b0011100100001011111010101;
    rom[31330] = 25'b0011100100010111101001100;
    rom[31331] = 25'b0011100100100011011000000;
    rom[31332] = 25'b0011100100101111000110011;
    rom[31333] = 25'b0011100100111010110100101;
    rom[31334] = 25'b0011100101000110100010100;
    rom[31335] = 25'b0011100101010010010000010;
    rom[31336] = 25'b0011100101011101111101111;
    rom[31337] = 25'b0011100101101001101011010;
    rom[31338] = 25'b0011100101110101011000100;
    rom[31339] = 25'b0011100110000001000101100;
    rom[31340] = 25'b0011100110001100110010010;
    rom[31341] = 25'b0011100110011000011110110;
    rom[31342] = 25'b0011100110100100001011010;
    rom[31343] = 25'b0011100110101111110111011;
    rom[31344] = 25'b0011100110111011100011100;
    rom[31345] = 25'b0011100111000111001111010;
    rom[31346] = 25'b0011100111010010111010110;
    rom[31347] = 25'b0011100111011110100110001;
    rom[31348] = 25'b0011100111101010010001011;
    rom[31349] = 25'b0011100111110101111100011;
    rom[31350] = 25'b0011101000000001100111001;
    rom[31351] = 25'b0011101000001101010001110;
    rom[31352] = 25'b0011101000011000111100000;
    rom[31353] = 25'b0011101000100100100110010;
    rom[31354] = 25'b0011101000110000010000001;
    rom[31355] = 25'b0011101000111011111010000;
    rom[31356] = 25'b0011101001000111100011100;
    rom[31357] = 25'b0011101001010011001100110;
    rom[31358] = 25'b0011101001011110110101111;
    rom[31359] = 25'b0011101001101010011110111;
    rom[31360] = 25'b0011101001110110000111100;
    rom[31361] = 25'b0011101010000001110000000;
    rom[31362] = 25'b0011101010001101011000011;
    rom[31363] = 25'b0011101010011001000000011;
    rom[31364] = 25'b0011101010100100101000010;
    rom[31365] = 25'b0011101010110000001111111;
    rom[31366] = 25'b0011101010111011110111011;
    rom[31367] = 25'b0011101011000111011110100;
    rom[31368] = 25'b0011101011010011000101100;
    rom[31369] = 25'b0011101011011110101100011;
    rom[31370] = 25'b0011101011101010010010111;
    rom[31371] = 25'b0011101011110101111001010;
    rom[31372] = 25'b0011101100000001011111011;
    rom[31373] = 25'b0011101100001101000101011;
    rom[31374] = 25'b0011101100011000101011000;
    rom[31375] = 25'b0011101100100100010000100;
    rom[31376] = 25'b0011101100101111110101110;
    rom[31377] = 25'b0011101100111011011010110;
    rom[31378] = 25'b0011101101000110111111101;
    rom[31379] = 25'b0011101101010010100100010;
    rom[31380] = 25'b0011101101011110001000101;
    rom[31381] = 25'b0011101101101001101100111;
    rom[31382] = 25'b0011101101110101010000110;
    rom[31383] = 25'b0011101110000000110100100;
    rom[31384] = 25'b0011101110001100010111111;
    rom[31385] = 25'b0011101110010111111011010;
    rom[31386] = 25'b0011101110100011011110010;
    rom[31387] = 25'b0011101110101111000001001;
    rom[31388] = 25'b0011101110111010100011101;
    rom[31389] = 25'b0011101111000110000110000;
    rom[31390] = 25'b0011101111010001101000001;
    rom[31391] = 25'b0011101111011101001010000;
    rom[31392] = 25'b0011101111101000101011110;
    rom[31393] = 25'b0011101111110100001101001;
    rom[31394] = 25'b0011101111111111101110011;
    rom[31395] = 25'b0011110000001011001111011;
    rom[31396] = 25'b0011110000010110110000001;
    rom[31397] = 25'b0011110000100010010000101;
    rom[31398] = 25'b0011110000101101110001000;
    rom[31399] = 25'b0011110000111001010001000;
    rom[31400] = 25'b0011110001000100110000111;
    rom[31401] = 25'b0011110001010000010000100;
    rom[31402] = 25'b0011110001011011101111110;
    rom[31403] = 25'b0011110001100111001110111;
    rom[31404] = 25'b0011110001110010101101110;
    rom[31405] = 25'b0011110001111110001100100;
    rom[31406] = 25'b0011110010001001101010111;
    rom[31407] = 25'b0011110010010101001001001;
    rom[31408] = 25'b0011110010100000100111000;
    rom[31409] = 25'b0011110010101100000100101;
    rom[31410] = 25'b0011110010110111100010001;
    rom[31411] = 25'b0011110011000010111111011;
    rom[31412] = 25'b0011110011001110011100011;
    rom[31413] = 25'b0011110011011001111001001;
    rom[31414] = 25'b0011110011100101010101101;
    rom[31415] = 25'b0011110011110000110001111;
    rom[31416] = 25'b0011110011111100001101111;
    rom[31417] = 25'b0011110100000111101001101;
    rom[31418] = 25'b0011110100010011000101010;
    rom[31419] = 25'b0011110100011110100000100;
    rom[31420] = 25'b0011110100101001111011100;
    rom[31421] = 25'b0011110100110101010110010;
    rom[31422] = 25'b0011110101000000110000111;
    rom[31423] = 25'b0011110101001100001011001;
    rom[31424] = 25'b0011110101010111100101010;
    rom[31425] = 25'b0011110101100010111111001;
    rom[31426] = 25'b0011110101101110011000101;
    rom[31427] = 25'b0011110101111001110001111;
    rom[31428] = 25'b0011110110000101001011000;
    rom[31429] = 25'b0011110110010000100011111;
    rom[31430] = 25'b0011110110011011111100011;
    rom[31431] = 25'b0011110110100111010100101;
    rom[31432] = 25'b0011110110110010101100110;
    rom[31433] = 25'b0011110110111110000100101;
    rom[31434] = 25'b0011110111001001011100000;
    rom[31435] = 25'b0011110111010100110011011;
    rom[31436] = 25'b0011110111100000001010100;
    rom[31437] = 25'b0011110111101011100001010;
    rom[31438] = 25'b0011110111110110110111110;
    rom[31439] = 25'b0011111000000010001110000;
    rom[31440] = 25'b0011111000001101100100001;
    rom[31441] = 25'b0011111000011000111001111;
    rom[31442] = 25'b0011111000100100001111011;
    rom[31443] = 25'b0011111000101111100100101;
    rom[31444] = 25'b0011111000111010111001101;
    rom[31445] = 25'b0011111001000110001110011;
    rom[31446] = 25'b0011111001010001100010111;
    rom[31447] = 25'b0011111001011100110111000;
    rom[31448] = 25'b0011111001101000001011000;
    rom[31449] = 25'b0011111001110011011110110;
    rom[31450] = 25'b0011111001111110110010001;
    rom[31451] = 25'b0011111010001010000101010;
    rom[31452] = 25'b0011111010010101011000010;
    rom[31453] = 25'b0011111010100000101010111;
    rom[31454] = 25'b0011111010101011111101010;
    rom[31455] = 25'b0011111010110111001111011;
    rom[31456] = 25'b0011111011000010100001010;
    rom[31457] = 25'b0011111011001101110010111;
    rom[31458] = 25'b0011111011011001000100001;
    rom[31459] = 25'b0011111011100100010101010;
    rom[31460] = 25'b0011111011101111100110000;
    rom[31461] = 25'b0011111011111010110110100;
    rom[31462] = 25'b0011111100000110000110110;
    rom[31463] = 25'b0011111100010001010110110;
    rom[31464] = 25'b0011111100011100100110011;
    rom[31465] = 25'b0011111100100111110101111;
    rom[31466] = 25'b0011111100110011000101000;
    rom[31467] = 25'b0011111100111110010011111;
    rom[31468] = 25'b0011111101001001100010100;
    rom[31469] = 25'b0011111101010100110000111;
    rom[31470] = 25'b0011111101011111111111000;
    rom[31471] = 25'b0011111101101011001100110;
    rom[31472] = 25'b0011111101110110011010010;
    rom[31473] = 25'b0011111110000001100111101;
    rom[31474] = 25'b0011111110001100110100100;
    rom[31475] = 25'b0011111110011000000001010;
    rom[31476] = 25'b0011111110100011001101101;
    rom[31477] = 25'b0011111110101110011001110;
    rom[31478] = 25'b0011111110111001100101110;
    rom[31479] = 25'b0011111111000100110001010;
    rom[31480] = 25'b0011111111001111111100101;
    rom[31481] = 25'b0011111111011011000111101;
    rom[31482] = 25'b0011111111100110010010011;
    rom[31483] = 25'b0011111111110001011100111;
    rom[31484] = 25'b0011111111111100100111000;
    rom[31485] = 25'b0100000000000111110000111;
    rom[31486] = 25'b0100000000010010111010101;
    rom[31487] = 25'b0100000000011110000100000;
    rom[31488] = 25'b0100000000101001001101000;
    rom[31489] = 25'b0100000000110100010101110;
    rom[31490] = 25'b0100000000111111011110010;
    rom[31491] = 25'b0100000001001010100110011;
    rom[31492] = 25'b0100000001010101101110011;
    rom[31493] = 25'b0100000001100000110110000;
    rom[31494] = 25'b0100000001101011111101011;
    rom[31495] = 25'b0100000001110111000100011;
    rom[31496] = 25'b0100000010000010001011001;
    rom[31497] = 25'b0100000010001101010001101;
    rom[31498] = 25'b0100000010011000010111111;
    rom[31499] = 25'b0100000010100011011101110;
    rom[31500] = 25'b0100000010101110100011011;
    rom[31501] = 25'b0100000010111001101000110;
    rom[31502] = 25'b0100000011000100101101110;
    rom[31503] = 25'b0100000011001111110010100;
    rom[31504] = 25'b0100000011011010110110111;
    rom[31505] = 25'b0100000011100101111011001;
    rom[31506] = 25'b0100000011110000111111000;
    rom[31507] = 25'b0100000011111100000010100;
    rom[31508] = 25'b0100000100000111000101110;
    rom[31509] = 25'b0100000100010010001000110;
    rom[31510] = 25'b0100000100011101001011100;
    rom[31511] = 25'b0100000100101000001101111;
    rom[31512] = 25'b0100000100110011010000000;
    rom[31513] = 25'b0100000100111110010001110;
    rom[31514] = 25'b0100000101001001010011010;
    rom[31515] = 25'b0100000101010100010100011;
    rom[31516] = 25'b0100000101011111010101011;
    rom[31517] = 25'b0100000101101010010101111;
    rom[31518] = 25'b0100000101110101010110010;
    rom[31519] = 25'b0100000110000000010110010;
    rom[31520] = 25'b0100000110001011010101111;
    rom[31521] = 25'b0100000110010110010101010;
    rom[31522] = 25'b0100000110100001010100011;
    rom[31523] = 25'b0100000110101100010011001;
    rom[31524] = 25'b0100000110110111010001101;
    rom[31525] = 25'b0100000111000010001111110;
    rom[31526] = 25'b0100000111001101001101101;
    rom[31527] = 25'b0100000111011000001011010;
    rom[31528] = 25'b0100000111100011001000100;
    rom[31529] = 25'b0100000111101110000101100;
    rom[31530] = 25'b0100000111111001000010001;
    rom[31531] = 25'b0100001000000011111110100;
    rom[31532] = 25'b0100001000001110111010100;
    rom[31533] = 25'b0100001000011001110110001;
    rom[31534] = 25'b0100001000100100110001101;
    rom[31535] = 25'b0100001000101111101100110;
    rom[31536] = 25'b0100001000111010100111100;
    rom[31537] = 25'b0100001001000101100010000;
    rom[31538] = 25'b0100001001010000011100001;
    rom[31539] = 25'b0100001001011011010110000;
    rom[31540] = 25'b0100001001100110001111100;
    rom[31541] = 25'b0100001001110001001000110;
    rom[31542] = 25'b0100001001111100000001110;
    rom[31543] = 25'b0100001010000110111010011;
    rom[31544] = 25'b0100001010010001110010101;
    rom[31545] = 25'b0100001010011100101010101;
    rom[31546] = 25'b0100001010100111100010010;
    rom[31547] = 25'b0100001010110010011001101;
    rom[31548] = 25'b0100001010111101010000101;
    rom[31549] = 25'b0100001011001000000111011;
    rom[31550] = 25'b0100001011010010111101110;
    rom[31551] = 25'b0100001011011101110011110;
    rom[31552] = 25'b0100001011101000101001100;
    rom[31553] = 25'b0100001011110011011111000;
    rom[31554] = 25'b0100001011111110010100000;
    rom[31555] = 25'b0100001100001001001000111;
    rom[31556] = 25'b0100001100010011111101011;
    rom[31557] = 25'b0100001100011110110001100;
    rom[31558] = 25'b0100001100101001100101011;
    rom[31559] = 25'b0100001100110100011000110;
    rom[31560] = 25'b0100001100111111001100000;
    rom[31561] = 25'b0100001101001001111110111;
    rom[31562] = 25'b0100001101010100110001011;
    rom[31563] = 25'b0100001101011111100011100;
    rom[31564] = 25'b0100001101101010010101100;
    rom[31565] = 25'b0100001101110101000111001;
    rom[31566] = 25'b0100001101111111111000010;
    rom[31567] = 25'b0100001110001010101001001;
    rom[31568] = 25'b0100001110010101011001110;
    rom[31569] = 25'b0100001110100000001010000;
    rom[31570] = 25'b0100001110101010111001111;
    rom[31571] = 25'b0100001110110101101001100;
    rom[31572] = 25'b0100001111000000011000110;
    rom[31573] = 25'b0100001111001011000111101;
    rom[31574] = 25'b0100001111010101110110010;
    rom[31575] = 25'b0100001111100000100100100;
    rom[31576] = 25'b0100001111101011010010011;
    rom[31577] = 25'b0100001111110110000000000;
    rom[31578] = 25'b0100010000000000101101010;
    rom[31579] = 25'b0100010000001011011010010;
    rom[31580] = 25'b0100010000010110000110110;
    rom[31581] = 25'b0100010000100000110011000;
    rom[31582] = 25'b0100010000101011011111000;
    rom[31583] = 25'b0100010000110110001010100;
    rom[31584] = 25'b0100010001000000110101110;
    rom[31585] = 25'b0100010001001011100000110;
    rom[31586] = 25'b0100010001010110001011010;
    rom[31587] = 25'b0100010001100000110101100;
    rom[31588] = 25'b0100010001101011011111011;
    rom[31589] = 25'b0100010001110110001000111;
    rom[31590] = 25'b0100010010000000110010001;
    rom[31591] = 25'b0100010010001011011011000;
    rom[31592] = 25'b0100010010010110000011101;
    rom[31593] = 25'b0100010010100000101011110;
    rom[31594] = 25'b0100010010101011010011101;
    rom[31595] = 25'b0100010010110101111011000;
    rom[31596] = 25'b0100010011000000100010010;
    rom[31597] = 25'b0100010011001011001001001;
    rom[31598] = 25'b0100010011010101101111100;
    rom[31599] = 25'b0100010011100000010101101;
    rom[31600] = 25'b0100010011101010111011011;
    rom[31601] = 25'b0100010011110101100000111;
    rom[31602] = 25'b0100010100000000000101111;
    rom[31603] = 25'b0100010100001010101010101;
    rom[31604] = 25'b0100010100010101001111001;
    rom[31605] = 25'b0100010100011111110011001;
    rom[31606] = 25'b0100010100101010010110111;
    rom[31607] = 25'b0100010100110100111010001;
    rom[31608] = 25'b0100010100111111011101001;
    rom[31609] = 25'b0100010101001001111111110;
    rom[31610] = 25'b0100010101010100100010001;
    rom[31611] = 25'b0100010101011111000100000;
    rom[31612] = 25'b0100010101101001100101101;
    rom[31613] = 25'b0100010101110100000110111;
    rom[31614] = 25'b0100010101111110100111110;
    rom[31615] = 25'b0100010110001001001000010;
    rom[31616] = 25'b0100010110010011101000100;
    rom[31617] = 25'b0100010110011110001000010;
    rom[31618] = 25'b0100010110101000100111110;
    rom[31619] = 25'b0100010110110011000110111;
    rom[31620] = 25'b0100010110111101100101101;
    rom[31621] = 25'b0100010111001000000100000;
    rom[31622] = 25'b0100010111010010100010001;
    rom[31623] = 25'b0100010111011100111111110;
    rom[31624] = 25'b0100010111100111011101001;
    rom[31625] = 25'b0100010111110001111010001;
    rom[31626] = 25'b0100010111111100010110101;
    rom[31627] = 25'b0100011000000110110010111;
    rom[31628] = 25'b0100011000010001001110111;
    rom[31629] = 25'b0100011000011011101010010;
    rom[31630] = 25'b0100011000100110000101100;
    rom[31631] = 25'b0100011000110000100000010;
    rom[31632] = 25'b0100011000111010111010110;
    rom[31633] = 25'b0100011001000101010100110;
    rom[31634] = 25'b0100011001001111101110100;
    rom[31635] = 25'b0100011001011010000111111;
    rom[31636] = 25'b0100011001100100100000110;
    rom[31637] = 25'b0100011001101110111001100;
    rom[31638] = 25'b0100011001111001010001110;
    rom[31639] = 25'b0100011010000011101001101;
    rom[31640] = 25'b0100011010001110000001001;
    rom[31641] = 25'b0100011010011000011000010;
    rom[31642] = 25'b0100011010100010101111000;
    rom[31643] = 25'b0100011010101101000101011;
    rom[31644] = 25'b0100011010110111011011011;
    rom[31645] = 25'b0100011011000001110001001;
    rom[31646] = 25'b0100011011001100000110100;
    rom[31647] = 25'b0100011011010110011011011;
    rom[31648] = 25'b0100011011100000110000000;
    rom[31649] = 25'b0100011011101011000100001;
    rom[31650] = 25'b0100011011110101010111111;
    rom[31651] = 25'b0100011011111111101011011;
    rom[31652] = 25'b0100011100001001111110011;
    rom[31653] = 25'b0100011100010100010001001;
    rom[31654] = 25'b0100011100011110100011100;
    rom[31655] = 25'b0100011100101000110101011;
    rom[31656] = 25'b0100011100110011000111000;
    rom[31657] = 25'b0100011100111101011000001;
    rom[31658] = 25'b0100011101000111101001000;
    rom[31659] = 25'b0100011101010001111001100;
    rom[31660] = 25'b0100011101011100001001100;
    rom[31661] = 25'b0100011101100110011001010;
    rom[31662] = 25'b0100011101110000101000100;
    rom[31663] = 25'b0100011101111010110111011;
    rom[31664] = 25'b0100011110000101000110000;
    rom[31665] = 25'b0100011110001111010100001;
    rom[31666] = 25'b0100011110011001100010000;
    rom[31667] = 25'b0100011110100011101111010;
    rom[31668] = 25'b0100011110101101111100011;
    rom[31669] = 25'b0100011110111000001001000;
    rom[31670] = 25'b0100011111000010010101010;
    rom[31671] = 25'b0100011111001100100001001;
    rom[31672] = 25'b0100011111010110101100101;
    rom[31673] = 25'b0100011111100000110111110;
    rom[31674] = 25'b0100011111101011000010100;
    rom[31675] = 25'b0100011111110101001100110;
    rom[31676] = 25'b0100011111111111010110101;
    rom[31677] = 25'b0100100000001001100000010;
    rom[31678] = 25'b0100100000010011101001011;
    rom[31679] = 25'b0100100000011101110010001;
    rom[31680] = 25'b0100100000100111111010101;
    rom[31681] = 25'b0100100000110010000010101;
    rom[31682] = 25'b0100100000111100001010010;
    rom[31683] = 25'b0100100001000110010001100;
    rom[31684] = 25'b0100100001010000011000010;
    rom[31685] = 25'b0100100001011010011110110;
    rom[31686] = 25'b0100100001100100100100111;
    rom[31687] = 25'b0100100001101110101010100;
    rom[31688] = 25'b0100100001111000101111110;
    rom[31689] = 25'b0100100010000010110100101;
    rom[31690] = 25'b0100100010001100111001001;
    rom[31691] = 25'b0100100010010110111101010;
    rom[31692] = 25'b0100100010100001000000111;
    rom[31693] = 25'b0100100010101011000100001;
    rom[31694] = 25'b0100100010110101000111001;
    rom[31695] = 25'b0100100010111111001001101;
    rom[31696] = 25'b0100100011001001001011101;
    rom[31697] = 25'b0100100011010011001101100;
    rom[31698] = 25'b0100100011011101001110110;
    rom[31699] = 25'b0100100011100111001111101;
    rom[31700] = 25'b0100100011110001010000001;
    rom[31701] = 25'b0100100011111011010000011;
    rom[31702] = 25'b0100100100000101010000000;
    rom[31703] = 25'b0100100100001111001111011;
    rom[31704] = 25'b0100100100011001001110011;
    rom[31705] = 25'b0100100100100011001100111;
    rom[31706] = 25'b0100100100101101001010111;
    rom[31707] = 25'b0100100100110111001000101;
    rom[31708] = 25'b0100100101000001000110000;
    rom[31709] = 25'b0100100101001011000010111;
    rom[31710] = 25'b0100100101010100111111011;
    rom[31711] = 25'b0100100101011110111011100;
    rom[31712] = 25'b0100100101101000110111010;
    rom[31713] = 25'b0100100101110010110010100;
    rom[31714] = 25'b0100100101111100101101011;
    rom[31715] = 25'b0100100110000110100111111;
    rom[31716] = 25'b0100100110010000100010000;
    rom[31717] = 25'b0100100110011010011011101;
    rom[31718] = 25'b0100100110100100010100111;
    rom[31719] = 25'b0100100110101110001101110;
    rom[31720] = 25'b0100100110111000000110001;
    rom[31721] = 25'b0100100111000001111110001;
    rom[31722] = 25'b0100100111001011110101111;
    rom[31723] = 25'b0100100111010101101101000;
    rom[31724] = 25'b0100100111011111100011110;
    rom[31725] = 25'b0100100111101001011010010;
    rom[31726] = 25'b0100100111110011010000010;
    rom[31727] = 25'b0100100111111101000101110;
    rom[31728] = 25'b0100101000000110111010111;
    rom[31729] = 25'b0100101000010000101111101;
    rom[31730] = 25'b0100101000011010100100000;
    rom[31731] = 25'b0100101000100100010111111;
    rom[31732] = 25'b0100101000101110001011011;
    rom[31733] = 25'b0100101000110111111110100;
    rom[31734] = 25'b0100101001000001110001001;
    rom[31735] = 25'b0100101001001011100011011;
    rom[31736] = 25'b0100101001010101010101001;
    rom[31737] = 25'b0100101001011111000110100;
    rom[31738] = 25'b0100101001101000110111101;
    rom[31739] = 25'b0100101001110010101000001;
    rom[31740] = 25'b0100101001111100011000010;
    rom[31741] = 25'b0100101010000110001000001;
    rom[31742] = 25'b0100101010001111110111011;
    rom[31743] = 25'b0100101010011001100110010;
    rom[31744] = 25'b0100101010100011010100110;
    rom[31745] = 25'b0100101010101101000010111;
    rom[31746] = 25'b0100101010110110110000011;
    rom[31747] = 25'b0100101011000000011101101;
    rom[31748] = 25'b0100101011001010001010100;
    rom[31749] = 25'b0100101011010011110110110;
    rom[31750] = 25'b0100101011011101100010110;
    rom[31751] = 25'b0100101011100111001110010;
    rom[31752] = 25'b0100101011110000111001011;
    rom[31753] = 25'b0100101011111010100100000;
    rom[31754] = 25'b0100101100000100001110010;
    rom[31755] = 25'b0100101100001101111000000;
    rom[31756] = 25'b0100101100010111100001011;
    rom[31757] = 25'b0100101100100001001010011;
    rom[31758] = 25'b0100101100101010110010111;
    rom[31759] = 25'b0100101100110100011011000;
    rom[31760] = 25'b0100101100111110000010101;
    rom[31761] = 25'b0100101101000111101001111;
    rom[31762] = 25'b0100101101010001010000110;
    rom[31763] = 25'b0100101101011010110111001;
    rom[31764] = 25'b0100101101100100011101000;
    rom[31765] = 25'b0100101101101110000010100;
    rom[31766] = 25'b0100101101110111100111100;
    rom[31767] = 25'b0100101110000001001100010;
    rom[31768] = 25'b0100101110001010110000011;
    rom[31769] = 25'b0100101110010100010100010;
    rom[31770] = 25'b0100101110011101110111101;
    rom[31771] = 25'b0100101110100111011010100;
    rom[31772] = 25'b0100101110110000111101000;
    rom[31773] = 25'b0100101110111010011111000;
    rom[31774] = 25'b0100101111000100000000101;
    rom[31775] = 25'b0100101111001101100001110;
    rom[31776] = 25'b0100101111010111000010100;
    rom[31777] = 25'b0100101111100000100010111;
    rom[31778] = 25'b0100101111101010000010101;
    rom[31779] = 25'b0100101111110011100010001;
    rom[31780] = 25'b0100101111111101000001001;
    rom[31781] = 25'b0100110000000110011111101;
    rom[31782] = 25'b0100110000001111111101110;
    rom[31783] = 25'b0100110000011001011011011;
    rom[31784] = 25'b0100110000100010111000101;
    rom[31785] = 25'b0100110000101100010101011;
    rom[31786] = 25'b0100110000110101110001101;
    rom[31787] = 25'b0100110000111111001101101;
    rom[31788] = 25'b0100110001001000101001000;
    rom[31789] = 25'b0100110001010010000100000;
    rom[31790] = 25'b0100110001011011011110101;
    rom[31791] = 25'b0100110001100100111000110;
    rom[31792] = 25'b0100110001101110010010011;
    rom[31793] = 25'b0100110001110111101011101;
    rom[31794] = 25'b0100110010000001000100011;
    rom[31795] = 25'b0100110010001010011100110;
    rom[31796] = 25'b0100110010010011110100101;
    rom[31797] = 25'b0100110010011101001100001;
    rom[31798] = 25'b0100110010100110100011001;
    rom[31799] = 25'b0100110010101111111001101;
    rom[31800] = 25'b0100110010111001001111101;
    rom[31801] = 25'b0100110011000010100101011;
    rom[31802] = 25'b0100110011001011111010100;
    rom[31803] = 25'b0100110011010101001111010;
    rom[31804] = 25'b0100110011011110100011100;
    rom[31805] = 25'b0100110011100111110111011;
    rom[31806] = 25'b0100110011110001001010110;
    rom[31807] = 25'b0100110011111010011101110;
    rom[31808] = 25'b0100110100000011110000001;
    rom[31809] = 25'b0100110100001101000010010;
    rom[31810] = 25'b0100110100010110010011110;
    rom[31811] = 25'b0100110100011111100101000;
    rom[31812] = 25'b0100110100101000110101101;
    rom[31813] = 25'b0100110100110010000101110;
    rom[31814] = 25'b0100110100111011010101100;
    rom[31815] = 25'b0100110101000100100100111;
    rom[31816] = 25'b0100110101001101110011110;
    rom[31817] = 25'b0100110101010111000010001;
    rom[31818] = 25'b0100110101100000010000001;
    rom[31819] = 25'b0100110101101001011101100;
    rom[31820] = 25'b0100110101110010101010100;
    rom[31821] = 25'b0100110101111011110111000;
    rom[31822] = 25'b0100110110000101000011010;
    rom[31823] = 25'b0100110110001110001110110;
    rom[31824] = 25'b0100110110010111011010000;
    rom[31825] = 25'b0100110110100000100100101;
    rom[31826] = 25'b0100110110101001101111000;
    rom[31827] = 25'b0100110110110010111000110;
    rom[31828] = 25'b0100110110111100000010000;
    rom[31829] = 25'b0100110111000101001010111;
    rom[31830] = 25'b0100110111001110010011011;
    rom[31831] = 25'b0100110111010111011011010;
    rom[31832] = 25'b0100110111100000100010110;
    rom[31833] = 25'b0100110111101001101001110;
    rom[31834] = 25'b0100110111110010110000010;
    rom[31835] = 25'b0100110111111011110110010;
    rom[31836] = 25'b0100111000000100111011111;
    rom[31837] = 25'b0100111000001110000001000;
    rom[31838] = 25'b0100111000010111000101110;
    rom[31839] = 25'b0100111000100000001010000;
    rom[31840] = 25'b0100111000101001001101110;
    rom[31841] = 25'b0100111000110010010001000;
    rom[31842] = 25'b0100111000111011010011110;
    rom[31843] = 25'b0100111001000100010110001;
    rom[31844] = 25'b0100111001001101011000000;
    rom[31845] = 25'b0100111001010110011001011;
    rom[31846] = 25'b0100111001011111011010010;
    rom[31847] = 25'b0100111001101000011010110;
    rom[31848] = 25'b0100111001110001011010101;
    rom[31849] = 25'b0100111001111010011010010;
    rom[31850] = 25'b0100111010000011011001010;
    rom[31851] = 25'b0100111010001100010111110;
    rom[31852] = 25'b0100111010010101010101111;
    rom[31853] = 25'b0100111010011110010011100;
    rom[31854] = 25'b0100111010100111010000101;
    rom[31855] = 25'b0100111010110000001101010;
    rom[31856] = 25'b0100111010111001001001100;
    rom[31857] = 25'b0100111011000010000101010;
    rom[31858] = 25'b0100111011001011000000100;
    rom[31859] = 25'b0100111011010011111011010;
    rom[31860] = 25'b0100111011011100110101100;
    rom[31861] = 25'b0100111011100101101111010;
    rom[31862] = 25'b0100111011101110101000101;
    rom[31863] = 25'b0100111011110111100001011;
    rom[31864] = 25'b0100111100000000011001110;
    rom[31865] = 25'b0100111100001001010001101;
    rom[31866] = 25'b0100111100010010001001001;
    rom[31867] = 25'b0100111100011011000000000;
    rom[31868] = 25'b0100111100100011110110011;
    rom[31869] = 25'b0100111100101100101100011;
    rom[31870] = 25'b0100111100110101100001111;
    rom[31871] = 25'b0100111100111110010110111;
    rom[31872] = 25'b0100111101000111001011011;
    rom[31873] = 25'b0100111101001111111111011;
    rom[31874] = 25'b0100111101011000110011000;
    rom[31875] = 25'b0100111101100001100110000;
    rom[31876] = 25'b0100111101101010011000100;
    rom[31877] = 25'b0100111101110011001010101;
    rom[31878] = 25'b0100111101111011111100010;
    rom[31879] = 25'b0100111110000100101101011;
    rom[31880] = 25'b0100111110001101011110000;
    rom[31881] = 25'b0100111110010110001110001;
    rom[31882] = 25'b0100111110011110111101111;
    rom[31883] = 25'b0100111110100111101101000;
    rom[31884] = 25'b0100111110110000011011110;
    rom[31885] = 25'b0100111110111001001001111;
    rom[31886] = 25'b0100111111000001110111101;
    rom[31887] = 25'b0100111111001010100100110;
    rom[31888] = 25'b0100111111010011010001100;
    rom[31889] = 25'b0100111111011011111101110;
    rom[31890] = 25'b0100111111100100101001100;
    rom[31891] = 25'b0100111111101101010100101;
    rom[31892] = 25'b0100111111110101111111100;
    rom[31893] = 25'b0100111111111110101001110;
    rom[31894] = 25'b0101000000000111010011100;
    rom[31895] = 25'b0101000000001111111100110;
    rom[31896] = 25'b0101000000011000100101100;
    rom[31897] = 25'b0101000000100001001101110;
    rom[31898] = 25'b0101000000101001110101101;
    rom[31899] = 25'b0101000000110010011100111;
    rom[31900] = 25'b0101000000111011000011101;
    rom[31901] = 25'b0101000001000011101010000;
    rom[31902] = 25'b0101000001001100001111110;
    rom[31903] = 25'b0101000001010100110101000;
    rom[31904] = 25'b0101000001011101011001111;
    rom[31905] = 25'b0101000001100101111110001;
    rom[31906] = 25'b0101000001101110100010000;
    rom[31907] = 25'b0101000001110111000101010;
    rom[31908] = 25'b0101000001111111101000001;
    rom[31909] = 25'b0101000010001000001010100;
    rom[31910] = 25'b0101000010010000101100010;
    rom[31911] = 25'b0101000010011001001101100;
    rom[31912] = 25'b0101000010100001101110011;
    rom[31913] = 25'b0101000010101010001110110;
    rom[31914] = 25'b0101000010110010101110100;
    rom[31915] = 25'b0101000010111011001101111;
    rom[31916] = 25'b0101000011000011101100101;
    rom[31917] = 25'b0101000011001100001010111;
    rom[31918] = 25'b0101000011010100101000110;
    rom[31919] = 25'b0101000011011101000110000;
    rom[31920] = 25'b0101000011100101100010110;
    rom[31921] = 25'b0101000011101101111111000;
    rom[31922] = 25'b0101000011110110011010111;
    rom[31923] = 25'b0101000011111110110110001;
    rom[31924] = 25'b0101000100000111010000111;
    rom[31925] = 25'b0101000100001111101011001;
    rom[31926] = 25'b0101000100011000000100111;
    rom[31927] = 25'b0101000100100000011110000;
    rom[31928] = 25'b0101000100101000110110111;
    rom[31929] = 25'b0101000100110001001111000;
    rom[31930] = 25'b0101000100111001100110110;
    rom[31931] = 25'b0101000101000001111101111;
    rom[31932] = 25'b0101000101001010010100101;
    rom[31933] = 25'b0101000101010010101010111;
    rom[31934] = 25'b0101000101011011000000100;
    rom[31935] = 25'b0101000101100011010101110;
    rom[31936] = 25'b0101000101101011101010010;
    rom[31937] = 25'b0101000101110011111110011;
    rom[31938] = 25'b0101000101111100010010000;
    rom[31939] = 25'b0101000110000100100101001;
    rom[31940] = 25'b0101000110001100110111110;
    rom[31941] = 25'b0101000110010101001001111;
    rom[31942] = 25'b0101000110011101011011011;
    rom[31943] = 25'b0101000110100101101100100;
    rom[31944] = 25'b0101000110101101111101000;
    rom[31945] = 25'b0101000110110110001101000;
    rom[31946] = 25'b0101000110111110011100100;
    rom[31947] = 25'b0101000111000110101011100;
    rom[31948] = 25'b0101000111001110111010000;
    rom[31949] = 25'b0101000111010111001000000;
    rom[31950] = 25'b0101000111011111010101011;
    rom[31951] = 25'b0101000111100111100010010;
    rom[31952] = 25'b0101000111101111101110101;
    rom[31953] = 25'b0101000111110111111010100;
    rom[31954] = 25'b0101001000000000000101111;
    rom[31955] = 25'b0101001000001000010000110;
    rom[31956] = 25'b0101001000010000011011001;
    rom[31957] = 25'b0101001000011000100100111;
    rom[31958] = 25'b0101001000100000101110001;
    rom[31959] = 25'b0101001000101000110110111;
    rom[31960] = 25'b0101001000110000111111001;
    rom[31961] = 25'b0101001000111001000110110;
    rom[31962] = 25'b0101001001000001001101111;
    rom[31963] = 25'b0101001001001001010100101;
    rom[31964] = 25'b0101001001010001011010110;
    rom[31965] = 25'b0101001001011001100000011;
    rom[31966] = 25'b0101001001100001100101100;
    rom[31967] = 25'b0101001001101001101010001;
    rom[31968] = 25'b0101001001110001101110000;
    rom[31969] = 25'b0101001001111001110001101;
    rom[31970] = 25'b0101001010000001110100100;
    rom[31971] = 25'b0101001010001001110111000;
    rom[31972] = 25'b0101001010010001111000111;
    rom[31973] = 25'b0101001010011001111010011;
    rom[31974] = 25'b0101001010100001111011010;
    rom[31975] = 25'b0101001010101001111011101;
    rom[31976] = 25'b0101001010110001111011011;
    rom[31977] = 25'b0101001010111001111010101;
    rom[31978] = 25'b0101001011000001111001011;
    rom[31979] = 25'b0101001011001001110111101;
    rom[31980] = 25'b0101001011010001110101011;
    rom[31981] = 25'b0101001011011001110010100;
    rom[31982] = 25'b0101001011100001101111001;
    rom[31983] = 25'b0101001011101001101011001;
    rom[31984] = 25'b0101001011110001100110110;
    rom[31985] = 25'b0101001011111001100001111;
    rom[31986] = 25'b0101001100000001011100010;
    rom[31987] = 25'b0101001100001001010110010;
    rom[31988] = 25'b0101001100010001001111110;
    rom[31989] = 25'b0101001100011001001000101;
    rom[31990] = 25'b0101001100100001000001000;
    rom[31991] = 25'b0101001100101000111000110;
    rom[31992] = 25'b0101001100110000110000001;
    rom[31993] = 25'b0101001100111000100110111;
    rom[31994] = 25'b0101001101000000011101001;
    rom[31995] = 25'b0101001101001000010010110;
    rom[31996] = 25'b0101001101010000000111111;
    rom[31997] = 25'b0101001101010111111100100;
    rom[31998] = 25'b0101001101011111110000100;
    rom[31999] = 25'b0101001101100111100100000;
    rom[32000] = 25'b0101001101101111010111000;
    rom[32001] = 25'b0101001101110111001001100;
    rom[32002] = 25'b0101001101111110111011100;
    rom[32003] = 25'b0101001110000110101100111;
    rom[32004] = 25'b0101001110001110011101101;
    rom[32005] = 25'b0101001110010110001101111;
    rom[32006] = 25'b0101001110011101111101101;
    rom[32007] = 25'b0101001110100101101100111;
    rom[32008] = 25'b0101001110101101011011100;
    rom[32009] = 25'b0101001110110101001001101;
    rom[32010] = 25'b0101001110111100110111001;
    rom[32011] = 25'b0101001111000100100100010;
    rom[32012] = 25'b0101001111001100010000110;
    rom[32013] = 25'b0101001111010011111100101;
    rom[32014] = 25'b0101001111011011101000000;
    rom[32015] = 25'b0101001111100011010010111;
    rom[32016] = 25'b0101001111101010111101010;
    rom[32017] = 25'b0101001111110010100111000;
    rom[32018] = 25'b0101001111111010010000010;
    rom[32019] = 25'b0101010000000001111000111;
    rom[32020] = 25'b0101010000001001100001000;
    rom[32021] = 25'b0101010000010001001000101;
    rom[32022] = 25'b0101010000011000101111101;
    rom[32023] = 25'b0101010000100000010110001;
    rom[32024] = 25'b0101010000100111111100000;
    rom[32025] = 25'b0101010000101111100001011;
    rom[32026] = 25'b0101010000110111000110010;
    rom[32027] = 25'b0101010000111110101010100;
    rom[32028] = 25'b0101010001000110001110010;
    rom[32029] = 25'b0101010001001101110001011;
    rom[32030] = 25'b0101010001010101010100000;
    rom[32031] = 25'b0101010001011100110110001;
    rom[32032] = 25'b0101010001100100010111101;
    rom[32033] = 25'b0101010001101011111000101;
    rom[32034] = 25'b0101010001110011011001000;
    rom[32035] = 25'b0101010001111010111000111;
    rom[32036] = 25'b0101010010000010011000001;
    rom[32037] = 25'b0101010010001001110111000;
    rom[32038] = 25'b0101010010010001010101001;
    rom[32039] = 25'b0101010010011000110010110;
    rom[32040] = 25'b0101010010100000001111111;
    rom[32041] = 25'b0101010010100111101100011;
    rom[32042] = 25'b0101010010101111001000011;
    rom[32043] = 25'b0101010010110110100011111;
    rom[32044] = 25'b0101010010111101111110101;
    rom[32045] = 25'b0101010011000101011001000;
    rom[32046] = 25'b0101010011001100110010110;
    rom[32047] = 25'b0101010011010100001011111;
    rom[32048] = 25'b0101010011011011100100100;
    rom[32049] = 25'b0101010011100010111100101;
    rom[32050] = 25'b0101010011101010010100010;
    rom[32051] = 25'b0101010011110001101011001;
    rom[32052] = 25'b0101010011111001000001100;
    rom[32053] = 25'b0101010100000000010111011;
    rom[32054] = 25'b0101010100000111101100101;
    rom[32055] = 25'b0101010100001111000001011;
    rom[32056] = 25'b0101010100010110010101100;
    rom[32057] = 25'b0101010100011101101001001;
    rom[32058] = 25'b0101010100100100111100001;
    rom[32059] = 25'b0101010100101100001110101;
    rom[32060] = 25'b0101010100110011100000100;
    rom[32061] = 25'b0101010100111010110001111;
    rom[32062] = 25'b0101010101000010000010101;
    rom[32063] = 25'b0101010101001001010010111;
    rom[32064] = 25'b0101010101010000100010011;
    rom[32065] = 25'b0101010101010111110001100;
    rom[32066] = 25'b0101010101011111000000001;
    rom[32067] = 25'b0101010101100110001110000;
    rom[32068] = 25'b0101010101101101011011011;
    rom[32069] = 25'b0101010101110100101000001;
    rom[32070] = 25'b0101010101111011110100100;
    rom[32071] = 25'b0101010110000011000000001;
    rom[32072] = 25'b0101010110001010001011010;
    rom[32073] = 25'b0101010110010001010101111;
    rom[32074] = 25'b0101010110011000011111110;
    rom[32075] = 25'b0101010110011111101001010;
    rom[32076] = 25'b0101010110100110110010000;
    rom[32077] = 25'b0101010110101101111010011;
    rom[32078] = 25'b0101010110110101000010000;
    rom[32079] = 25'b0101010110111100001001001;
    rom[32080] = 25'b0101010111000011001111101;
    rom[32081] = 25'b0101010111001010010101110;
    rom[32082] = 25'b0101010111010001011011001;
    rom[32083] = 25'b0101010111011000100000000;
    rom[32084] = 25'b0101010111011111100100010;
    rom[32085] = 25'b0101010111100110100111111;
    rom[32086] = 25'b0101010111101101101011001;
    rom[32087] = 25'b0101010111110100101101101;
    rom[32088] = 25'b0101010111111011101111101;
    rom[32089] = 25'b0101011000000010110001000;
    rom[32090] = 25'b0101011000001001110001111;
    rom[32091] = 25'b0101011000010000110010001;
    rom[32092] = 25'b0101011000010111110001110;
    rom[32093] = 25'b0101011000011110110000111;
    rom[32094] = 25'b0101011000100101101111100;
    rom[32095] = 25'b0101011000101100101101011;
    rom[32096] = 25'b0101011000110011101010110;
    rom[32097] = 25'b0101011000111010100111101;
    rom[32098] = 25'b0101011001000001100011110;
    rom[32099] = 25'b0101011001001000011111100;
    rom[32100] = 25'b0101011001001111011010100;
    rom[32101] = 25'b0101011001010110010101000;
    rom[32102] = 25'b0101011001011101001110111;
    rom[32103] = 25'b0101011001100100001000010;
    rom[32104] = 25'b0101011001101011000001000;
    rom[32105] = 25'b0101011001110001111001001;
    rom[32106] = 25'b0101011001111000110000111;
    rom[32107] = 25'b0101011001111111100111111;
    rom[32108] = 25'b0101011010000110011110010;
    rom[32109] = 25'b0101011010001101010100001;
    rom[32110] = 25'b0101011010010100001001011;
    rom[32111] = 25'b0101011010011010111110000;
    rom[32112] = 25'b0101011010100001110010001;
    rom[32113] = 25'b0101011010101000100101101;
    rom[32114] = 25'b0101011010101111011000101;
    rom[32115] = 25'b0101011010110110001010111;
    rom[32116] = 25'b0101011010111100111100110;
    rom[32117] = 25'b0101011011000011101101111;
    rom[32118] = 25'b0101011011001010011110100;
    rom[32119] = 25'b0101011011010001001110100;
    rom[32120] = 25'b0101011011010111111110000;
    rom[32121] = 25'b0101011011011110101100110;
    rom[32122] = 25'b0101011011100101011011001;
    rom[32123] = 25'b0101011011101100001000110;
    rom[32124] = 25'b0101011011110010110101110;
    rom[32125] = 25'b0101011011111001100010011;
    rom[32126] = 25'b0101011100000000001110010;
    rom[32127] = 25'b0101011100000110111001101;
    rom[32128] = 25'b0101011100001101100100010;
    rom[32129] = 25'b0101011100010100001110100;
    rom[32130] = 25'b0101011100011010111000000;
    rom[32131] = 25'b0101011100100001100001000;
    rom[32132] = 25'b0101011100101000001001010;
    rom[32133] = 25'b0101011100101110110001001;
    rom[32134] = 25'b0101011100110101011000011;
    rom[32135] = 25'b0101011100111011111110111;
    rom[32136] = 25'b0101011101000010100100111;
    rom[32137] = 25'b0101011101001001001010011;
    rom[32138] = 25'b0101011101001111101111001;
    rom[32139] = 25'b0101011101010110010011011;
    rom[32140] = 25'b0101011101011100110111001;
    rom[32141] = 25'b0101011101100011011010001;
    rom[32142] = 25'b0101011101101001111100101;
    rom[32143] = 25'b0101011101110000011110100;
    rom[32144] = 25'b0101011101110110111111110;
    rom[32145] = 25'b0101011101111101100000011;
    rom[32146] = 25'b0101011110000100000000100;
    rom[32147] = 25'b0101011110001010100000000;
    rom[32148] = 25'b0101011110010000111110111;
    rom[32149] = 25'b0101011110010111011101010;
    rom[32150] = 25'b0101011110011101111010111;
    rom[32151] = 25'b0101011110100100011000000;
    rom[32152] = 25'b0101011110101010110100101;
    rom[32153] = 25'b0101011110110001010000011;
    rom[32154] = 25'b0101011110110111101011110;
    rom[32155] = 25'b0101011110111110000110100;
    rom[32156] = 25'b0101011111000100100000101;
    rom[32157] = 25'b0101011111001010111010001;
    rom[32158] = 25'b0101011111010001010011001;
    rom[32159] = 25'b0101011111010111101011011;
    rom[32160] = 25'b0101011111011110000011001;
    rom[32161] = 25'b0101011111100100011010010;
    rom[32162] = 25'b0101011111101010110000110;
    rom[32163] = 25'b0101011111110001000110101;
    rom[32164] = 25'b0101011111110111011100000;
    rom[32165] = 25'b0101011111111101110000110;
    rom[32166] = 25'b0101100000000100000100111;
    rom[32167] = 25'b0101100000001010011000011;
    rom[32168] = 25'b0101100000010000101011010;
    rom[32169] = 25'b0101100000010110111101101;
    rom[32170] = 25'b0101100000011101001111011;
    rom[32171] = 25'b0101100000100011100000011;
    rom[32172] = 25'b0101100000101001110001000;
    rom[32173] = 25'b0101100000110000000000111;
    rom[32174] = 25'b0101100000110110010000001;
    rom[32175] = 25'b0101100000111100011110111;
    rom[32176] = 25'b0101100001000010101101000;
    rom[32177] = 25'b0101100001001000111010011;
    rom[32178] = 25'b0101100001001111000111010;
    rom[32179] = 25'b0101100001010101010011101;
    rom[32180] = 25'b0101100001011011011111010;
    rom[32181] = 25'b0101100001100001101010011;
    rom[32182] = 25'b0101100001100111110100110;
    rom[32183] = 25'b0101100001101101111110101;
    rom[32184] = 25'b0101100001110100000111111;
    rom[32185] = 25'b0101100001111010010000100;
    rom[32186] = 25'b0101100010000000011000100;
    rom[32187] = 25'b0101100010000110100000000;
    rom[32188] = 25'b0101100010001100100110110;
    rom[32189] = 25'b0101100010010010101101000;
    rom[32190] = 25'b0101100010011000110010101;
    rom[32191] = 25'b0101100010011110110111100;
    rom[32192] = 25'b0101100010100100111100000;
    rom[32193] = 25'b0101100010101010111111101;
    rom[32194] = 25'b0101100010110001000010110;
    rom[32195] = 25'b0101100010110111000101011;
    rom[32196] = 25'b0101100010111101000111010;
    rom[32197] = 25'b0101100011000011001000101;
    rom[32198] = 25'b0101100011001001001001011;
    rom[32199] = 25'b0101100011001111001001100;
    rom[32200] = 25'b0101100011010101001000111;
    rom[32201] = 25'b0101100011011011000111110;
    rom[32202] = 25'b0101100011100001000110000;
    rom[32203] = 25'b0101100011100111000011101;
    rom[32204] = 25'b0101100011101101000000110;
    rom[32205] = 25'b0101100011110010111101001;
    rom[32206] = 25'b0101100011111000111000111;
    rom[32207] = 25'b0101100011111110110100001;
    rom[32208] = 25'b0101100100000100101110101;
    rom[32209] = 25'b0101100100001010101000100;
    rom[32210] = 25'b0101100100010000100001111;
    rom[32211] = 25'b0101100100010110011010101;
    rom[32212] = 25'b0101100100011100010010110;
    rom[32213] = 25'b0101100100100010001010010;
    rom[32214] = 25'b0101100100101000000001001;
    rom[32215] = 25'b0101100100101101110111011;
    rom[32216] = 25'b0101100100110011101101000;
    rom[32217] = 25'b0101100100111001100010000;
    rom[32218] = 25'b0101100100111111010110011;
    rom[32219] = 25'b0101100101000101001010010;
    rom[32220] = 25'b0101100101001010111101011;
    rom[32221] = 25'b0101100101010000101111111;
    rom[32222] = 25'b0101100101010110100001111;
    rom[32223] = 25'b0101100101011100010011001;
    rom[32224] = 25'b0101100101100010000011111;
    rom[32225] = 25'b0101100101100111110011111;
    rom[32226] = 25'b0101100101101101100011011;
    rom[32227] = 25'b0101100101110011010010001;
    rom[32228] = 25'b0101100101111001000000011;
    rom[32229] = 25'b0101100101111110101110000;
    rom[32230] = 25'b0101100110000100011010111;
    rom[32231] = 25'b0101100110001010000111010;
    rom[32232] = 25'b0101100110001111110011000;
    rom[32233] = 25'b0101100110010101011110000;
    rom[32234] = 25'b0101100110011011001000101;
    rom[32235] = 25'b0101100110100000110010011;
    rom[32236] = 25'b0101100110100110011011101;
    rom[32237] = 25'b0101100110101100000100010;
    rom[32238] = 25'b0101100110110001101100001;
    rom[32239] = 25'b0101100110110111010011100;
    rom[32240] = 25'b0101100110111100111010010;
    rom[32241] = 25'b0101100111000010100000011;
    rom[32242] = 25'b0101100111001000000101111;
    rom[32243] = 25'b0101100111001101101010101;
    rom[32244] = 25'b0101100111010011001110111;
    rom[32245] = 25'b0101100111011000110010100;
    rom[32246] = 25'b0101100111011110010101011;
    rom[32247] = 25'b0101100111100011110111111;
    rom[32248] = 25'b0101100111101001011001100;
    rom[32249] = 25'b0101100111101110111010101;
    rom[32250] = 25'b0101100111110100011011000;
    rom[32251] = 25'b0101100111111001111010111;
    rom[32252] = 25'b0101100111111111011010001;
    rom[32253] = 25'b0101101000000100111000110;
    rom[32254] = 25'b0101101000001010010110101;
    rom[32255] = 25'b0101101000001111110011111;
    rom[32256] = 25'b0101101000010101010000101;
    rom[32257] = 25'b0101101000011010101100101;
    rom[32258] = 25'b0101101000100000001000000;
    rom[32259] = 25'b0101101000100101100010111;
    rom[32260] = 25'b0101101000101010111101001;
    rom[32261] = 25'b0101101000110000010110101;
    rom[32262] = 25'b0101101000110101101111100;
    rom[32263] = 25'b0101101000111011000111110;
    rom[32264] = 25'b0101101001000000011111011;
    rom[32265] = 25'b0101101001000101110110011;
    rom[32266] = 25'b0101101001001011001100110;
    rom[32267] = 25'b0101101001010000100010100;
    rom[32268] = 25'b0101101001010101110111101;
    rom[32269] = 25'b0101101001011011001100001;
    rom[32270] = 25'b0101101001100000011111111;
    rom[32271] = 25'b0101101001100101110011010;
    rom[32272] = 25'b0101101001101011000101110;
    rom[32273] = 25'b0101101001110000010111101;
    rom[32274] = 25'b0101101001110101101001000;
    rom[32275] = 25'b0101101001111010111001101;
    rom[32276] = 25'b0101101010000000001001101;
    rom[32277] = 25'b0101101010000101011001000;
    rom[32278] = 25'b0101101010001010100111110;
    rom[32279] = 25'b0101101010001111110110000;
    rom[32280] = 25'b0101101010010101000011011;
    rom[32281] = 25'b0101101010011010010000010;
    rom[32282] = 25'b0101101010011111011100100;
    rom[32283] = 25'b0101101010100100101000000;
    rom[32284] = 25'b0101101010101001110011000;
    rom[32285] = 25'b0101101010101110111101011;
    rom[32286] = 25'b0101101010110100000111000;
    rom[32287] = 25'b0101101010111001010000000;
    rom[32288] = 25'b0101101010111110011000011;
    rom[32289] = 25'b0101101011000011100000001;
    rom[32290] = 25'b0101101011001000100111010;
    rom[32291] = 25'b0101101011001101101101110;
    rom[32292] = 25'b0101101011010010110011101;
    rom[32293] = 25'b0101101011010111111000110;
    rom[32294] = 25'b0101101011011100111101010;
    rom[32295] = 25'b0101101011100010000001010;
    rom[32296] = 25'b0101101011100111000100100;
    rom[32297] = 25'b0101101011101100000111001;
    rom[32298] = 25'b0101101011110001001001001;
    rom[32299] = 25'b0101101011110110001010011;
    rom[32300] = 25'b0101101011111011001011001;
    rom[32301] = 25'b0101101100000000001011001;
    rom[32302] = 25'b0101101100000101001010101;
    rom[32303] = 25'b0101101100001010001001011;
    rom[32304] = 25'b0101101100001111000111100;
    rom[32305] = 25'b0101101100010100000101000;
    rom[32306] = 25'b0101101100011001000001111;
    rom[32307] = 25'b0101101100011101111110000;
    rom[32308] = 25'b0101101100100010111001101;
    rom[32309] = 25'b0101101100100111110100100;
    rom[32310] = 25'b0101101100101100101110111;
    rom[32311] = 25'b0101101100110001101000011;
    rom[32312] = 25'b0101101100110110100001011;
    rom[32313] = 25'b0101101100111011011001110;
    rom[32314] = 25'b0101101101000000010001100;
    rom[32315] = 25'b0101101101000101001000100;
    rom[32316] = 25'b0101101101001001111110111;
    rom[32317] = 25'b0101101101001110110100101;
    rom[32318] = 25'b0101101101010011101001110;
    rom[32319] = 25'b0101101101011000011110010;
    rom[32320] = 25'b0101101101011101010010000;
    rom[32321] = 25'b0101101101100010000101001;
    rom[32322] = 25'b0101101101100110110111101;
    rom[32323] = 25'b0101101101101011101001100;
    rom[32324] = 25'b0101101101110000011010110;
    rom[32325] = 25'b0101101101110101001011010;
    rom[32326] = 25'b0101101101111001111011010;
    rom[32327] = 25'b0101101101111110101010100;
    rom[32328] = 25'b0101101110000011011001001;
    rom[32329] = 25'b0101101110001000000111001;
    rom[32330] = 25'b0101101110001100110100100;
    rom[32331] = 25'b0101101110010001100001001;
    rom[32332] = 25'b0101101110010110001101001;
    rom[32333] = 25'b0101101110011010111000100;
    rom[32334] = 25'b0101101110011111100011001;
    rom[32335] = 25'b0101101110100100001101010;
    rom[32336] = 25'b0101101110101000110110110;
    rom[32337] = 25'b0101101110101101011111100;
    rom[32338] = 25'b0101101110110010000111101;
    rom[32339] = 25'b0101101110110110101111000;
    rom[32340] = 25'b0101101110111011010101111;
    rom[32341] = 25'b0101101110111111111100000;
    rom[32342] = 25'b0101101111000100100001100;
    rom[32343] = 25'b0101101111001001000110011;
    rom[32344] = 25'b0101101111001101101010101;
    rom[32345] = 25'b0101101111010010001110001;
    rom[32346] = 25'b0101101111010110110001000;
    rom[32347] = 25'b0101101111011011010011010;
    rom[32348] = 25'b0101101111011111110100111;
    rom[32349] = 25'b0101101111100100010101110;
    rom[32350] = 25'b0101101111101000110110001;
    rom[32351] = 25'b0101101111101101010101101;
    rom[32352] = 25'b0101101111110001110100101;
    rom[32353] = 25'b0101101111110110010011000;
    rom[32354] = 25'b0101101111111010110000101;
    rom[32355] = 25'b0101101111111111001101101;
    rom[32356] = 25'b0101110000000011101010000;
    rom[32357] = 25'b0101110000001000000101101;
    rom[32358] = 25'b0101110000001100100000101;
    rom[32359] = 25'b0101110000010000111011001;
    rom[32360] = 25'b0101110000010101010100110;
    rom[32361] = 25'b0101110000011001101101111;
    rom[32362] = 25'b0101110000011110000110010;
    rom[32363] = 25'b0101110000100010011110000;
    rom[32364] = 25'b0101110000100110110101001;
    rom[32365] = 25'b0101110000101011001011100;
    rom[32366] = 25'b0101110000101111100001010;
    rom[32367] = 25'b0101110000110011110110011;
    rom[32368] = 25'b0101110000111000001010110;
    rom[32369] = 25'b0101110000111100011110101;
    rom[32370] = 25'b0101110001000000110001110;
    rom[32371] = 25'b0101110001000101000100010;
    rom[32372] = 25'b0101110001001001010110000;
    rom[32373] = 25'b0101110001001101100111010;
    rom[32374] = 25'b0101110001010001110111101;
    rom[32375] = 25'b0101110001010110000111100;
    rom[32376] = 25'b0101110001011010010110101;
    rom[32377] = 25'b0101110001011110100101010;
    rom[32378] = 25'b0101110001100010110011000;
    rom[32379] = 25'b0101110001100111000000010;
    rom[32380] = 25'b0101110001101011001100110;
    rom[32381] = 25'b0101110001101111011000101;
    rom[32382] = 25'b0101110001110011100011111;
    rom[32383] = 25'b0101110001110111101110011;
    rom[32384] = 25'b0101110001111011111000010;
    rom[32385] = 25'b0101110010000000000001100;
    rom[32386] = 25'b0101110010000100001010000;
    rom[32387] = 25'b0101110010001000010001111;
    rom[32388] = 25'b0101110010001100011001001;
    rom[32389] = 25'b0101110010010000011111110;
    rom[32390] = 25'b0101110010010100100101101;
    rom[32391] = 25'b0101110010011000101010111;
    rom[32392] = 25'b0101110010011100101111011;
    rom[32393] = 25'b0101110010100000110011010;
    rom[32394] = 25'b0101110010100100110110100;
    rom[32395] = 25'b0101110010101000111001001;
    rom[32396] = 25'b0101110010101100111011000;
    rom[32397] = 25'b0101110010110000111100010;
    rom[32398] = 25'b0101110010110100111100111;
    rom[32399] = 25'b0101110010111000111100110;
    rom[32400] = 25'b0101110010111100111100000;
    rom[32401] = 25'b0101110011000000111010101;
    rom[32402] = 25'b0101110011000100111000100;
    rom[32403] = 25'b0101110011001000110101110;
    rom[32404] = 25'b0101110011001100110010011;
    rom[32405] = 25'b0101110011010000101110010;
    rom[32406] = 25'b0101110011010100101001100;
    rom[32407] = 25'b0101110011011000100100001;
    rom[32408] = 25'b0101110011011100011110000;
    rom[32409] = 25'b0101110011100000010111010;
    rom[32410] = 25'b0101110011100100001111111;
    rom[32411] = 25'b0101110011101000000111110;
    rom[32412] = 25'b0101110011101011111111000;
    rom[32413] = 25'b0101110011101111110101100;
    rom[32414] = 25'b0101110011110011101011011;
    rom[32415] = 25'b0101110011110111100000101;
    rom[32416] = 25'b0101110011111011010101010;
    rom[32417] = 25'b0101110011111111001001000;
    rom[32418] = 25'b0101110100000010111100011;
    rom[32419] = 25'b0101110100000110101110111;
    rom[32420] = 25'b0101110100001010100000110;
    rom[32421] = 25'b0101110100001110010010000;
    rom[32422] = 25'b0101110100010010000010100;
    rom[32423] = 25'b0101110100010101110010011;
    rom[32424] = 25'b0101110100011001100001101;
    rom[32425] = 25'b0101110100011101010000001;
    rom[32426] = 25'b0101110100100000111110000;
    rom[32427] = 25'b0101110100100100101011001;
    rom[32428] = 25'b0101110100101000010111110;
    rom[32429] = 25'b0101110100101100000011100;
    rom[32430] = 25'b0101110100101111101110101;
    rom[32431] = 25'b0101110100110011011001001;
    rom[32432] = 25'b0101110100110111000011000;
    rom[32433] = 25'b0101110100111010101100001;
    rom[32434] = 25'b0101110100111110010100101;
    rom[32435] = 25'b0101110101000001111100011;
    rom[32436] = 25'b0101110101000101100011100;
    rom[32437] = 25'b0101110101001001001010000;
    rom[32438] = 25'b0101110101001100101111111;
    rom[32439] = 25'b0101110101010000010100111;
    rom[32440] = 25'b0101110101010011111001011;
    rom[32441] = 25'b0101110101010111011101001;
    rom[32442] = 25'b0101110101011011000000010;
    rom[32443] = 25'b0101110101011110100010101;
    rom[32444] = 25'b0101110101100010000100011;
    rom[32445] = 25'b0101110101100101100101011;
    rom[32446] = 25'b0101110101101001000101110;
    rom[32447] = 25'b0101110101101100100101100;
    rom[32448] = 25'b0101110101110000000100100;
    rom[32449] = 25'b0101110101110011100010111;
    rom[32450] = 25'b0101110101110111000000101;
    rom[32451] = 25'b0101110101111010011101101;
    rom[32452] = 25'b0101110101111101111010000;
    rom[32453] = 25'b0101110110000001010101101;
    rom[32454] = 25'b0101110110000100110000101;
    rom[32455] = 25'b0101110110001000001010111;
    rom[32456] = 25'b0101110110001011100100100;
    rom[32457] = 25'b0101110110001110111101100;
    rom[32458] = 25'b0101110110010010010101110;
    rom[32459] = 25'b0101110110010101101101010;
    rom[32460] = 25'b0101110110011001000100001;
    rom[32461] = 25'b0101110110011100011010011;
    rom[32462] = 25'b0101110110011111110000000;
    rom[32463] = 25'b0101110110100011000100111;
    rom[32464] = 25'b0101110110100110011001001;
    rom[32465] = 25'b0101110110101001101100101;
    rom[32466] = 25'b0101110110101100111111100;
    rom[32467] = 25'b0101110110110000010001101;
    rom[32468] = 25'b0101110110110011100011000;
    rom[32469] = 25'b0101110110110110110011111;
    rom[32470] = 25'b0101110110111010000100000;
    rom[32471] = 25'b0101110110111101010011100;
    rom[32472] = 25'b0101110111000000100010010;
    rom[32473] = 25'b0101110111000011110000010;
    rom[32474] = 25'b0101110111000110111101110;
    rom[32475] = 25'b0101110111001010001010100;
    rom[32476] = 25'b0101110111001101010110100;
    rom[32477] = 25'b0101110111010000100001111;
    rom[32478] = 25'b0101110111010011101100100;
    rom[32479] = 25'b0101110111010110110110100;
    rom[32480] = 25'b0101110111011001111111111;
    rom[32481] = 25'b0101110111011101001000100;
    rom[32482] = 25'b0101110111100000010000011;
    rom[32483] = 25'b0101110111100011010111110;
    rom[32484] = 25'b0101110111100110011110011;
    rom[32485] = 25'b0101110111101001100100010;
    rom[32486] = 25'b0101110111101100101001100;
    rom[32487] = 25'b0101110111101111101110000;
    rom[32488] = 25'b0101110111110010110001111;
    rom[32489] = 25'b0101110111110101110101001;
    rom[32490] = 25'b0101110111111000110111100;
    rom[32491] = 25'b0101110111111011111001011;
    rom[32492] = 25'b0101110111111110111010100;
    rom[32493] = 25'b0101111000000001111010111;
    rom[32494] = 25'b0101111000000100111010110;
    rom[32495] = 25'b0101111000000111111001110;
    rom[32496] = 25'b0101111000001010111000001;
    rom[32497] = 25'b0101111000001101110101111;
    rom[32498] = 25'b0101111000010000110010111;
    rom[32499] = 25'b0101111000010011101111010;
    rom[32500] = 25'b0101111000010110101010111;
    rom[32501] = 25'b0101111000011001100101111;
    rom[32502] = 25'b0101111000011100100000001;
    rom[32503] = 25'b0101111000011111011001110;
    rom[32504] = 25'b0101111000100010010010101;
    rom[32505] = 25'b0101111000100101001010111;
    rom[32506] = 25'b0101111000101000000010011;
    rom[32507] = 25'b0101111000101010111001010;
    rom[32508] = 25'b0101111000101101101111100;
    rom[32509] = 25'b0101111000110000100100111;
    rom[32510] = 25'b0101111000110011011001110;
    rom[32511] = 25'b0101111000110110001101111;
    rom[32512] = 25'b0101111000111001000001010;
    rom[32513] = 25'b0101111000111011110100000;
    rom[32514] = 25'b0101111000111110100110001;
    rom[32515] = 25'b0101111001000001010111011;
    rom[32516] = 25'b0101111001000100001000001;
    rom[32517] = 25'b0101111001000110111000001;
    rom[32518] = 25'b0101111001001001100111100;
    rom[32519] = 25'b0101111001001100010110001;
    rom[32520] = 25'b0101111001001111000100000;
    rom[32521] = 25'b0101111001010001110001010;
    rom[32522] = 25'b0101111001010100011101110;
    rom[32523] = 25'b0101111001010111001001101;
    rom[32524] = 25'b0101111001011001110100110;
    rom[32525] = 25'b0101111001011100011111010;
    rom[32526] = 25'b0101111001011111001001001;
    rom[32527] = 25'b0101111001100001110010010;
    rom[32528] = 25'b0101111001100100011010101;
    rom[32529] = 25'b0101111001100111000010011;
    rom[32530] = 25'b0101111001101001101001100;
    rom[32531] = 25'b0101111001101100001111110;
    rom[32532] = 25'b0101111001101110110101100;
    rom[32533] = 25'b0101111001110001011010100;
    rom[32534] = 25'b0101111001110011111110110;
    rom[32535] = 25'b0101111001110110100010011;
    rom[32536] = 25'b0101111001111001000101010;
    rom[32537] = 25'b0101111001111011100111100;
    rom[32538] = 25'b0101111001111110001001000;
    rom[32539] = 25'b0101111010000000101001111;
    rom[32540] = 25'b0101111010000011001010000;
    rom[32541] = 25'b0101111010000101101001011;
    rom[32542] = 25'b0101111010001000001000001;
    rom[32543] = 25'b0101111010001010100110010;
    rom[32544] = 25'b0101111010001101000011101;
    rom[32545] = 25'b0101111010001111100000010;
    rom[32546] = 25'b0101111010010001111100011;
    rom[32547] = 25'b0101111010010100010111101;
    rom[32548] = 25'b0101111010010110110010010;
    rom[32549] = 25'b0101111010011001001100010;
    rom[32550] = 25'b0101111010011011100101100;
    rom[32551] = 25'b0101111010011101111110000;
    rom[32552] = 25'b0101111010100000010101110;
    rom[32553] = 25'b0101111010100010101101000;
    rom[32554] = 25'b0101111010100101000011100;
    rom[32555] = 25'b0101111010100111011001010;
    rom[32556] = 25'b0101111010101001101110010;
    rom[32557] = 25'b0101111010101100000010101;
    rom[32558] = 25'b0101111010101110010110011;
    rom[32559] = 25'b0101111010110000101001011;
    rom[32560] = 25'b0101111010110010111011101;
    rom[32561] = 25'b0101111010110101001101011;
    rom[32562] = 25'b0101111010110111011110010;
    rom[32563] = 25'b0101111010111001101110100;
    rom[32564] = 25'b0101111010111011111110000;
    rom[32565] = 25'b0101111010111110001100110;
    rom[32566] = 25'b0101111011000000011011000;
    rom[32567] = 25'b0101111011000010101000011;
    rom[32568] = 25'b0101111011000100110101010;
    rom[32569] = 25'b0101111011000111000001010;
    rom[32570] = 25'b0101111011001001001100101;
    rom[32571] = 25'b0101111011001011010111011;
    rom[32572] = 25'b0101111011001101100001010;
    rom[32573] = 25'b0101111011001111101010100;
    rom[32574] = 25'b0101111011010001110011001;
    rom[32575] = 25'b0101111011010011111011000;
    rom[32576] = 25'b0101111011010110000010010;
    rom[32577] = 25'b0101111011011000001000110;
    rom[32578] = 25'b0101111011011010001110100;
    rom[32579] = 25'b0101111011011100010011110;
    rom[32580] = 25'b0101111011011110011000001;
    rom[32581] = 25'b0101111011100000011011111;
    rom[32582] = 25'b0101111011100010011110111;
    rom[32583] = 25'b0101111011100100100001010;
    rom[32584] = 25'b0101111011100110100010111;
    rom[32585] = 25'b0101111011101000100011110;
    rom[32586] = 25'b0101111011101010100100000;
    rom[32587] = 25'b0101111011101100100011101;
    rom[32588] = 25'b0101111011101110100010011;
    rom[32589] = 25'b0101111011110000100000101;
    rom[32590] = 25'b0101111011110010011110001;
    rom[32591] = 25'b0101111011110100011010111;
    rom[32592] = 25'b0101111011110110010110111;
    rom[32593] = 25'b0101111011111000010010010;
    rom[32594] = 25'b0101111011111010001101000;
    rom[32595] = 25'b0101111011111100000110111;
    rom[32596] = 25'b0101111011111110000000010;
    rom[32597] = 25'b0101111011111111111000110;
    rom[32598] = 25'b0101111100000001110000110;
    rom[32599] = 25'b0101111100000011100111111;
    rom[32600] = 25'b0101111100000101011110011;
    rom[32601] = 25'b0101111100000111010100001;
    rom[32602] = 25'b0101111100001001001001010;
    rom[32603] = 25'b0101111100001010111101110;
    rom[32604] = 25'b0101111100001100110001011;
    rom[32605] = 25'b0101111100001110100100011;
    rom[32606] = 25'b0101111100010000010110101;
    rom[32607] = 25'b0101111100010010001000010;
    rom[32608] = 25'b0101111100010011111001010;
    rom[32609] = 25'b0101111100010101101001011;
    rom[32610] = 25'b0101111100010111011000111;
    rom[32611] = 25'b0101111100011001000111110;
    rom[32612] = 25'b0101111100011010110101111;
    rom[32613] = 25'b0101111100011100100011010;
    rom[32614] = 25'b0101111100011110010000000;
    rom[32615] = 25'b0101111100011111111100000;
    rom[32616] = 25'b0101111100100001100111010;
    rom[32617] = 25'b0101111100100011010001111;
    rom[32618] = 25'b0101111100100100111011110;
    rom[32619] = 25'b0101111100100110100101000;
    rom[32620] = 25'b0101111100101000001101100;
    rom[32621] = 25'b0101111100101001110101011;
    rom[32622] = 25'b0101111100101011011100100;
    rom[32623] = 25'b0101111100101101000010111;
    rom[32624] = 25'b0101111100101110101000101;
    rom[32625] = 25'b0101111100110000001101101;
    rom[32626] = 25'b0101111100110001110010000;
    rom[32627] = 25'b0101111100110011010101101;
    rom[32628] = 25'b0101111100110100111000100;
    rom[32629] = 25'b0101111100110110011010110;
    rom[32630] = 25'b0101111100110111111100010;
    rom[32631] = 25'b0101111100111001011101001;
    rom[32632] = 25'b0101111100111010111101010;
    rom[32633] = 25'b0101111100111100011100101;
    rom[32634] = 25'b0101111100111101111011011;
    rom[32635] = 25'b0101111100111111011001011;
    rom[32636] = 25'b0101111101000000110110101;
    rom[32637] = 25'b0101111101000010010011010;
    rom[32638] = 25'b0101111101000011101111010;
    rom[32639] = 25'b0101111101000101001010011;
    rom[32640] = 25'b0101111101000110100100111;
    rom[32641] = 25'b0101111101000111111110110;
    rom[32642] = 25'b0101111101001001010111111;
    rom[32643] = 25'b0101111101001010110000010;
    rom[32644] = 25'b0101111101001100001000000;
    rom[32645] = 25'b0101111101001101011111000;
    rom[32646] = 25'b0101111101001110110101010;
    rom[32647] = 25'b0101111101010000001010111;
    rom[32648] = 25'b0101111101010001011111111;
    rom[32649] = 25'b0101111101010010110100000;
    rom[32650] = 25'b0101111101010100000111100;
    rom[32651] = 25'b0101111101010101011010010;
    rom[32652] = 25'b0101111101010110101100011;
    rom[32653] = 25'b0101111101010111111101111;
    rom[32654] = 25'b0101111101011001001110100;
    rom[32655] = 25'b0101111101011010011110100;
    rom[32656] = 25'b0101111101011011101101110;
    rom[32657] = 25'b0101111101011100111100011;
    rom[32658] = 25'b0101111101011110001010010;
    rom[32659] = 25'b0101111101011111010111011;
    rom[32660] = 25'b0101111101100000100011111;
    rom[32661] = 25'b0101111101100001101111101;
    rom[32662] = 25'b0101111101100010111010101;
    rom[32663] = 25'b0101111101100100000101001;
    rom[32664] = 25'b0101111101100101001110110;
    rom[32665] = 25'b0101111101100110010111110;
    rom[32666] = 25'b0101111101100111011111111;
    rom[32667] = 25'b0101111101101000100111100;
    rom[32668] = 25'b0101111101101001101110011;
    rom[32669] = 25'b0101111101101010110100100;
    rom[32670] = 25'b0101111101101011111010000;
    rom[32671] = 25'b0101111101101100111110101;
    rom[32672] = 25'b0101111101101110000010110;
    rom[32673] = 25'b0101111101101111000110001;
    rom[32674] = 25'b0101111101110000001000110;
    rom[32675] = 25'b0101111101110001001010110;
    rom[32676] = 25'b0101111101110010001011111;
    rom[32677] = 25'b0101111101110011001100011;
    rom[32678] = 25'b0101111101110100001100010;
    rom[32679] = 25'b0101111101110101001011011;
    rom[32680] = 25'b0101111101110110001001110;
    rom[32681] = 25'b0101111101110111000111100;
    rom[32682] = 25'b0101111101111000000100100;
    rom[32683] = 25'b0101111101111001000000110;
    rom[32684] = 25'b0101111101111001111100011;
    rom[32685] = 25'b0101111101111010110111010;
    rom[32686] = 25'b0101111101111011110001100;
    rom[32687] = 25'b0101111101111100101011000;
    rom[32688] = 25'b0101111101111101100011110;
    rom[32689] = 25'b0101111101111110011011110;
    rom[32690] = 25'b0101111101111111010011001;
    rom[32691] = 25'b0101111110000000001001111;
    rom[32692] = 25'b0101111110000000111111111;
    rom[32693] = 25'b0101111110000001110101001;
    rom[32694] = 25'b0101111110000010101001101;
    rom[32695] = 25'b0101111110000011011101100;
    rom[32696] = 25'b0101111110000100010000101;
    rom[32697] = 25'b0101111110000101000011001;
    rom[32698] = 25'b0101111110000101110100111;
    rom[32699] = 25'b0101111110000110100101111;
    rom[32700] = 25'b0101111110000111010110001;
    rom[32701] = 25'b0101111110001000000101110;
    rom[32702] = 25'b0101111110001000110100110;
    rom[32703] = 25'b0101111110001001100010111;
    rom[32704] = 25'b0101111110001010010000100;
    rom[32705] = 25'b0101111110001010111101011;
    rom[32706] = 25'b0101111110001011101001011;
    rom[32707] = 25'b0101111110001100010100111;
    rom[32708] = 25'b0101111110001100111111100;
    rom[32709] = 25'b0101111110001101101001011;
    rom[32710] = 25'b0101111110001110010010110;
    rom[32711] = 25'b0101111110001110111011011;
    rom[32712] = 25'b0101111110001111100011010;
    rom[32713] = 25'b0101111110010000001010011;
    rom[32714] = 25'b0101111110010000110000110;
    rom[32715] = 25'b0101111110010001010110100;
    rom[32716] = 25'b0101111110010001111011101;
    rom[32717] = 25'b0101111110010010100000000;
    rom[32718] = 25'b0101111110010011000011101;
    rom[32719] = 25'b0101111110010011100110100;
    rom[32720] = 25'b0101111110010100001000111;
    rom[32721] = 25'b0101111110010100101010011;
    rom[32722] = 25'b0101111110010101001011001;
    rom[32723] = 25'b0101111110010101101011010;
    rom[32724] = 25'b0101111110010110001010101;
    rom[32725] = 25'b0101111110010110101001011;
    rom[32726] = 25'b0101111110010111000111011;
    rom[32727] = 25'b0101111110010111100100101;
    rom[32728] = 25'b0101111110011000000001010;
    rom[32729] = 25'b0101111110011000011101001;
    rom[32730] = 25'b0101111110011000111000011;
    rom[32731] = 25'b0101111110011001010010110;
    rom[32732] = 25'b0101111110011001101100100;
    rom[32733] = 25'b0101111110011010000101100;
    rom[32734] = 25'b0101111110011010011101111;
    rom[32735] = 25'b0101111110011010110101100;
    rom[32736] = 25'b0101111110011011001100100;
    rom[32737] = 25'b0101111110011011100010110;
    rom[32738] = 25'b0101111110011011111000011;
    rom[32739] = 25'b0101111110011100001101001;
    rom[32740] = 25'b0101111110011100100001010;
    rom[32741] = 25'b0101111110011100110100101;
    rom[32742] = 25'b0101111110011101000111011;
    rom[32743] = 25'b0101111110011101011001011;
    rom[32744] = 25'b0101111110011101101010101;
    rom[32745] = 25'b0101111110011101111011010;
    rom[32746] = 25'b0101111110011110001011001;
    rom[32747] = 25'b0101111110011110011010011;
    rom[32748] = 25'b0101111110011110101000111;
    rom[32749] = 25'b0101111110011110110110100;
    rom[32750] = 25'b0101111110011111000011101;
    rom[32751] = 25'b0101111110011111010000000;
    rom[32752] = 25'b0101111110011111011011101;
    rom[32753] = 25'b0101111110011111100110100;
    rom[32754] = 25'b0101111110011111110000111;
    rom[32755] = 25'b0101111110011111111010011;
    rom[32756] = 25'b0101111110100000000011001;
    rom[32757] = 25'b0101111110100000001011010;
    rom[32758] = 25'b0101111110100000010010101;
    rom[32759] = 25'b0101111110100000011001011;
    rom[32760] = 25'b0101111110100000011111011;
    rom[32761] = 25'b0101111110100000100100101;
    rom[32762] = 25'b0101111110100000101001010;
    rom[32763] = 25'b0101111110100000101101001;
    rom[32764] = 25'b0101111110100000110000011;
    rom[32765] = 25'b0101111110100000110010110;
    rom[32766] = 25'b0101111110100000110100100;
    rom[32767] = 25'b0101111110100000110101101;
    rom[32768] = 25'b0101111110100000110101111;
    rom[32769] = 25'b0101111110100000110101101;
    rom[32770] = 25'b0101111110100000110100100;
    rom[32771] = 25'b0101111110100000110010110;
    rom[32772] = 25'b0101111110100000110000011;
    rom[32773] = 25'b0101111110100000101101001;
    rom[32774] = 25'b0101111110100000101001010;
    rom[32775] = 25'b0101111110100000100100101;
    rom[32776] = 25'b0101111110100000011111011;
    rom[32777] = 25'b0101111110100000011001011;
    rom[32778] = 25'b0101111110100000010010101;
    rom[32779] = 25'b0101111110100000001011010;
    rom[32780] = 25'b0101111110100000000011001;
    rom[32781] = 25'b0101111110011111111010011;
    rom[32782] = 25'b0101111110011111110000111;
    rom[32783] = 25'b0101111110011111100110100;
    rom[32784] = 25'b0101111110011111011011101;
    rom[32785] = 25'b0101111110011111010000000;
    rom[32786] = 25'b0101111110011111000011101;
    rom[32787] = 25'b0101111110011110110110100;
    rom[32788] = 25'b0101111110011110101000111;
    rom[32789] = 25'b0101111110011110011010011;
    rom[32790] = 25'b0101111110011110001011001;
    rom[32791] = 25'b0101111110011101111011010;
    rom[32792] = 25'b0101111110011101101010101;
    rom[32793] = 25'b0101111110011101011001011;
    rom[32794] = 25'b0101111110011101000111011;
    rom[32795] = 25'b0101111110011100110100101;
    rom[32796] = 25'b0101111110011100100001010;
    rom[32797] = 25'b0101111110011100001101001;
    rom[32798] = 25'b0101111110011011111000011;
    rom[32799] = 25'b0101111110011011100010110;
    rom[32800] = 25'b0101111110011011001100100;
    rom[32801] = 25'b0101111110011010110101100;
    rom[32802] = 25'b0101111110011010011101111;
    rom[32803] = 25'b0101111110011010000101100;
    rom[32804] = 25'b0101111110011001101100100;
    rom[32805] = 25'b0101111110011001010010110;
    rom[32806] = 25'b0101111110011000111000011;
    rom[32807] = 25'b0101111110011000011101001;
    rom[32808] = 25'b0101111110011000000001010;
    rom[32809] = 25'b0101111110010111100100101;
    rom[32810] = 25'b0101111110010111000111011;
    rom[32811] = 25'b0101111110010110101001011;
    rom[32812] = 25'b0101111110010110001010101;
    rom[32813] = 25'b0101111110010101101011010;
    rom[32814] = 25'b0101111110010101001011001;
    rom[32815] = 25'b0101111110010100101010011;
    rom[32816] = 25'b0101111110010100001000111;
    rom[32817] = 25'b0101111110010011100110100;
    rom[32818] = 25'b0101111110010011000011101;
    rom[32819] = 25'b0101111110010010100000000;
    rom[32820] = 25'b0101111110010001111011101;
    rom[32821] = 25'b0101111110010001010110100;
    rom[32822] = 25'b0101111110010000110000110;
    rom[32823] = 25'b0101111110010000001010011;
    rom[32824] = 25'b0101111110001111100011010;
    rom[32825] = 25'b0101111110001110111011011;
    rom[32826] = 25'b0101111110001110010010110;
    rom[32827] = 25'b0101111110001101101001011;
    rom[32828] = 25'b0101111110001100111111100;
    rom[32829] = 25'b0101111110001100010100111;
    rom[32830] = 25'b0101111110001011101001011;
    rom[32831] = 25'b0101111110001010111101011;
    rom[32832] = 25'b0101111110001010010000100;
    rom[32833] = 25'b0101111110001001100010111;
    rom[32834] = 25'b0101111110001000110100110;
    rom[32835] = 25'b0101111110001000000101110;
    rom[32836] = 25'b0101111110000111010110001;
    rom[32837] = 25'b0101111110000110100101111;
    rom[32838] = 25'b0101111110000101110100111;
    rom[32839] = 25'b0101111110000101000011001;
    rom[32840] = 25'b0101111110000100010000101;
    rom[32841] = 25'b0101111110000011011101100;
    rom[32842] = 25'b0101111110000010101001101;
    rom[32843] = 25'b0101111110000001110101001;
    rom[32844] = 25'b0101111110000000111111111;
    rom[32845] = 25'b0101111110000000001001111;
    rom[32846] = 25'b0101111101111111010011001;
    rom[32847] = 25'b0101111101111110011011110;
    rom[32848] = 25'b0101111101111101100011110;
    rom[32849] = 25'b0101111101111100101011000;
    rom[32850] = 25'b0101111101111011110001100;
    rom[32851] = 25'b0101111101111010110111010;
    rom[32852] = 25'b0101111101111001111100011;
    rom[32853] = 25'b0101111101111001000000110;
    rom[32854] = 25'b0101111101111000000100100;
    rom[32855] = 25'b0101111101110111000111100;
    rom[32856] = 25'b0101111101110110001001110;
    rom[32857] = 25'b0101111101110101001011011;
    rom[32858] = 25'b0101111101110100001100010;
    rom[32859] = 25'b0101111101110011001100011;
    rom[32860] = 25'b0101111101110010001011111;
    rom[32861] = 25'b0101111101110001001010110;
    rom[32862] = 25'b0101111101110000001000110;
    rom[32863] = 25'b0101111101101111000110001;
    rom[32864] = 25'b0101111101101110000010110;
    rom[32865] = 25'b0101111101101100111110101;
    rom[32866] = 25'b0101111101101011111010000;
    rom[32867] = 25'b0101111101101010110100100;
    rom[32868] = 25'b0101111101101001101110011;
    rom[32869] = 25'b0101111101101000100111100;
    rom[32870] = 25'b0101111101100111011111111;
    rom[32871] = 25'b0101111101100110010111110;
    rom[32872] = 25'b0101111101100101001110110;
    rom[32873] = 25'b0101111101100100000101001;
    rom[32874] = 25'b0101111101100010111010101;
    rom[32875] = 25'b0101111101100001101111101;
    rom[32876] = 25'b0101111101100000100011111;
    rom[32877] = 25'b0101111101011111010111011;
    rom[32878] = 25'b0101111101011110001010010;
    rom[32879] = 25'b0101111101011100111100011;
    rom[32880] = 25'b0101111101011011101101110;
    rom[32881] = 25'b0101111101011010011110100;
    rom[32882] = 25'b0101111101011001001110100;
    rom[32883] = 25'b0101111101010111111101111;
    rom[32884] = 25'b0101111101010110101100011;
    rom[32885] = 25'b0101111101010101011010010;
    rom[32886] = 25'b0101111101010100000111100;
    rom[32887] = 25'b0101111101010010110100000;
    rom[32888] = 25'b0101111101010001011111111;
    rom[32889] = 25'b0101111101010000001010111;
    rom[32890] = 25'b0101111101001110110101010;
    rom[32891] = 25'b0101111101001101011111000;
    rom[32892] = 25'b0101111101001100001000000;
    rom[32893] = 25'b0101111101001010110000010;
    rom[32894] = 25'b0101111101001001010111111;
    rom[32895] = 25'b0101111101000111111110110;
    rom[32896] = 25'b0101111101000110100100111;
    rom[32897] = 25'b0101111101000101001010011;
    rom[32898] = 25'b0101111101000011101111010;
    rom[32899] = 25'b0101111101000010010011010;
    rom[32900] = 25'b0101111101000000110110101;
    rom[32901] = 25'b0101111100111111011001011;
    rom[32902] = 25'b0101111100111101111011011;
    rom[32903] = 25'b0101111100111100011100101;
    rom[32904] = 25'b0101111100111010111101010;
    rom[32905] = 25'b0101111100111001011101001;
    rom[32906] = 25'b0101111100110111111100010;
    rom[32907] = 25'b0101111100110110011010110;
    rom[32908] = 25'b0101111100110100111000100;
    rom[32909] = 25'b0101111100110011010101101;
    rom[32910] = 25'b0101111100110001110010000;
    rom[32911] = 25'b0101111100110000001101101;
    rom[32912] = 25'b0101111100101110101000101;
    rom[32913] = 25'b0101111100101101000010111;
    rom[32914] = 25'b0101111100101011011100100;
    rom[32915] = 25'b0101111100101001110101011;
    rom[32916] = 25'b0101111100101000001101100;
    rom[32917] = 25'b0101111100100110100101000;
    rom[32918] = 25'b0101111100100100111011110;
    rom[32919] = 25'b0101111100100011010001111;
    rom[32920] = 25'b0101111100100001100111010;
    rom[32921] = 25'b0101111100011111111100000;
    rom[32922] = 25'b0101111100011110010000000;
    rom[32923] = 25'b0101111100011100100011010;
    rom[32924] = 25'b0101111100011010110101111;
    rom[32925] = 25'b0101111100011001000111110;
    rom[32926] = 25'b0101111100010111011000111;
    rom[32927] = 25'b0101111100010101101001011;
    rom[32928] = 25'b0101111100010011111001010;
    rom[32929] = 25'b0101111100010010001000010;
    rom[32930] = 25'b0101111100010000010110101;
    rom[32931] = 25'b0101111100001110100100011;
    rom[32932] = 25'b0101111100001100110001011;
    rom[32933] = 25'b0101111100001010111101110;
    rom[32934] = 25'b0101111100001001001001010;
    rom[32935] = 25'b0101111100000111010100001;
    rom[32936] = 25'b0101111100000101011110011;
    rom[32937] = 25'b0101111100000011100111111;
    rom[32938] = 25'b0101111100000001110000110;
    rom[32939] = 25'b0101111011111111111000110;
    rom[32940] = 25'b0101111011111110000000010;
    rom[32941] = 25'b0101111011111100000110111;
    rom[32942] = 25'b0101111011111010001101000;
    rom[32943] = 25'b0101111011111000010010010;
    rom[32944] = 25'b0101111011110110010110111;
    rom[32945] = 25'b0101111011110100011010111;
    rom[32946] = 25'b0101111011110010011110001;
    rom[32947] = 25'b0101111011110000100000101;
    rom[32948] = 25'b0101111011101110100010011;
    rom[32949] = 25'b0101111011101100100011101;
    rom[32950] = 25'b0101111011101010100100000;
    rom[32951] = 25'b0101111011101000100011110;
    rom[32952] = 25'b0101111011100110100010111;
    rom[32953] = 25'b0101111011100100100001010;
    rom[32954] = 25'b0101111011100010011110111;
    rom[32955] = 25'b0101111011100000011011111;
    rom[32956] = 25'b0101111011011110011000001;
    rom[32957] = 25'b0101111011011100010011110;
    rom[32958] = 25'b0101111011011010001110100;
    rom[32959] = 25'b0101111011011000001000110;
    rom[32960] = 25'b0101111011010110000010010;
    rom[32961] = 25'b0101111011010011111011000;
    rom[32962] = 25'b0101111011010001110011001;
    rom[32963] = 25'b0101111011001111101010100;
    rom[32964] = 25'b0101111011001101100001010;
    rom[32965] = 25'b0101111011001011010111011;
    rom[32966] = 25'b0101111011001001001100101;
    rom[32967] = 25'b0101111011000111000001010;
    rom[32968] = 25'b0101111011000100110101010;
    rom[32969] = 25'b0101111011000010101000011;
    rom[32970] = 25'b0101111011000000011011000;
    rom[32971] = 25'b0101111010111110001100110;
    rom[32972] = 25'b0101111010111011111110000;
    rom[32973] = 25'b0101111010111001101110100;
    rom[32974] = 25'b0101111010110111011110010;
    rom[32975] = 25'b0101111010110101001101011;
    rom[32976] = 25'b0101111010110010111011101;
    rom[32977] = 25'b0101111010110000101001011;
    rom[32978] = 25'b0101111010101110010110011;
    rom[32979] = 25'b0101111010101100000010101;
    rom[32980] = 25'b0101111010101001101110010;
    rom[32981] = 25'b0101111010100111011001010;
    rom[32982] = 25'b0101111010100101000011100;
    rom[32983] = 25'b0101111010100010101101000;
    rom[32984] = 25'b0101111010100000010101110;
    rom[32985] = 25'b0101111010011101111110000;
    rom[32986] = 25'b0101111010011011100101100;
    rom[32987] = 25'b0101111010011001001100010;
    rom[32988] = 25'b0101111010010110110010010;
    rom[32989] = 25'b0101111010010100010111101;
    rom[32990] = 25'b0101111010010001111100011;
    rom[32991] = 25'b0101111010001111100000010;
    rom[32992] = 25'b0101111010001101000011101;
    rom[32993] = 25'b0101111010001010100110010;
    rom[32994] = 25'b0101111010001000001000001;
    rom[32995] = 25'b0101111010000101101001011;
    rom[32996] = 25'b0101111010000011001010000;
    rom[32997] = 25'b0101111010000000101001111;
    rom[32998] = 25'b0101111001111110001001000;
    rom[32999] = 25'b0101111001111011100111100;
    rom[33000] = 25'b0101111001111001000101010;
    rom[33001] = 25'b0101111001110110100010011;
    rom[33002] = 25'b0101111001110011111110110;
    rom[33003] = 25'b0101111001110001011010100;
    rom[33004] = 25'b0101111001101110110101100;
    rom[33005] = 25'b0101111001101100001111110;
    rom[33006] = 25'b0101111001101001101001100;
    rom[33007] = 25'b0101111001100111000010011;
    rom[33008] = 25'b0101111001100100011010101;
    rom[33009] = 25'b0101111001100001110010010;
    rom[33010] = 25'b0101111001011111001001001;
    rom[33011] = 25'b0101111001011100011111010;
    rom[33012] = 25'b0101111001011001110100110;
    rom[33013] = 25'b0101111001010111001001101;
    rom[33014] = 25'b0101111001010100011101110;
    rom[33015] = 25'b0101111001010001110001010;
    rom[33016] = 25'b0101111001001111000100000;
    rom[33017] = 25'b0101111001001100010110001;
    rom[33018] = 25'b0101111001001001100111100;
    rom[33019] = 25'b0101111001000110111000001;
    rom[33020] = 25'b0101111001000100001000001;
    rom[33021] = 25'b0101111001000001010111011;
    rom[33022] = 25'b0101111000111110100110001;
    rom[33023] = 25'b0101111000111011110100000;
    rom[33024] = 25'b0101111000111001000001010;
    rom[33025] = 25'b0101111000110110001101111;
    rom[33026] = 25'b0101111000110011011001110;
    rom[33027] = 25'b0101111000110000100100111;
    rom[33028] = 25'b0101111000101101101111100;
    rom[33029] = 25'b0101111000101010111001010;
    rom[33030] = 25'b0101111000101000000010011;
    rom[33031] = 25'b0101111000100101001010111;
    rom[33032] = 25'b0101111000100010010010101;
    rom[33033] = 25'b0101111000011111011001110;
    rom[33034] = 25'b0101111000011100100000001;
    rom[33035] = 25'b0101111000011001100101111;
    rom[33036] = 25'b0101111000010110101010111;
    rom[33037] = 25'b0101111000010011101111010;
    rom[33038] = 25'b0101111000010000110010111;
    rom[33039] = 25'b0101111000001101110101111;
    rom[33040] = 25'b0101111000001010111000001;
    rom[33041] = 25'b0101111000000111111001110;
    rom[33042] = 25'b0101111000000100111010110;
    rom[33043] = 25'b0101111000000001111010111;
    rom[33044] = 25'b0101110111111110111010100;
    rom[33045] = 25'b0101110111111011111001011;
    rom[33046] = 25'b0101110111111000110111100;
    rom[33047] = 25'b0101110111110101110101001;
    rom[33048] = 25'b0101110111110010110001111;
    rom[33049] = 25'b0101110111101111101110000;
    rom[33050] = 25'b0101110111101100101001100;
    rom[33051] = 25'b0101110111101001100100010;
    rom[33052] = 25'b0101110111100110011110011;
    rom[33053] = 25'b0101110111100011010111110;
    rom[33054] = 25'b0101110111100000010000011;
    rom[33055] = 25'b0101110111011101001000100;
    rom[33056] = 25'b0101110111011001111111111;
    rom[33057] = 25'b0101110111010110110110100;
    rom[33058] = 25'b0101110111010011101100100;
    rom[33059] = 25'b0101110111010000100001111;
    rom[33060] = 25'b0101110111001101010110100;
    rom[33061] = 25'b0101110111001010001010100;
    rom[33062] = 25'b0101110111000110111101110;
    rom[33063] = 25'b0101110111000011110000010;
    rom[33064] = 25'b0101110111000000100010010;
    rom[33065] = 25'b0101110110111101010011100;
    rom[33066] = 25'b0101110110111010000100000;
    rom[33067] = 25'b0101110110110110110011111;
    rom[33068] = 25'b0101110110110011100011000;
    rom[33069] = 25'b0101110110110000010001101;
    rom[33070] = 25'b0101110110101100111111100;
    rom[33071] = 25'b0101110110101001101100101;
    rom[33072] = 25'b0101110110100110011001001;
    rom[33073] = 25'b0101110110100011000100111;
    rom[33074] = 25'b0101110110011111110000000;
    rom[33075] = 25'b0101110110011100011010011;
    rom[33076] = 25'b0101110110011001000100001;
    rom[33077] = 25'b0101110110010101101101010;
    rom[33078] = 25'b0101110110010010010101110;
    rom[33079] = 25'b0101110110001110111101100;
    rom[33080] = 25'b0101110110001011100100100;
    rom[33081] = 25'b0101110110001000001010111;
    rom[33082] = 25'b0101110110000100110000101;
    rom[33083] = 25'b0101110110000001010101101;
    rom[33084] = 25'b0101110101111101111010000;
    rom[33085] = 25'b0101110101111010011101101;
    rom[33086] = 25'b0101110101110111000000101;
    rom[33087] = 25'b0101110101110011100010111;
    rom[33088] = 25'b0101110101110000000100100;
    rom[33089] = 25'b0101110101101100100101100;
    rom[33090] = 25'b0101110101101001000101110;
    rom[33091] = 25'b0101110101100101100101011;
    rom[33092] = 25'b0101110101100010000100011;
    rom[33093] = 25'b0101110101011110100010101;
    rom[33094] = 25'b0101110101011011000000010;
    rom[33095] = 25'b0101110101010111011101001;
    rom[33096] = 25'b0101110101010011111001011;
    rom[33097] = 25'b0101110101010000010100111;
    rom[33098] = 25'b0101110101001100101111111;
    rom[33099] = 25'b0101110101001001001010000;
    rom[33100] = 25'b0101110101000101100011100;
    rom[33101] = 25'b0101110101000001111100011;
    rom[33102] = 25'b0101110100111110010100101;
    rom[33103] = 25'b0101110100111010101100001;
    rom[33104] = 25'b0101110100110111000011000;
    rom[33105] = 25'b0101110100110011011001001;
    rom[33106] = 25'b0101110100101111101110101;
    rom[33107] = 25'b0101110100101100000011100;
    rom[33108] = 25'b0101110100101000010111110;
    rom[33109] = 25'b0101110100100100101011001;
    rom[33110] = 25'b0101110100100000111110000;
    rom[33111] = 25'b0101110100011101010000001;
    rom[33112] = 25'b0101110100011001100001101;
    rom[33113] = 25'b0101110100010101110010011;
    rom[33114] = 25'b0101110100010010000010100;
    rom[33115] = 25'b0101110100001110010010000;
    rom[33116] = 25'b0101110100001010100000110;
    rom[33117] = 25'b0101110100000110101110111;
    rom[33118] = 25'b0101110100000010111100011;
    rom[33119] = 25'b0101110011111111001001000;
    rom[33120] = 25'b0101110011111011010101010;
    rom[33121] = 25'b0101110011110111100000101;
    rom[33122] = 25'b0101110011110011101011011;
    rom[33123] = 25'b0101110011101111110101100;
    rom[33124] = 25'b0101110011101011111111000;
    rom[33125] = 25'b0101110011101000000111110;
    rom[33126] = 25'b0101110011100100001111111;
    rom[33127] = 25'b0101110011100000010111010;
    rom[33128] = 25'b0101110011011100011110000;
    rom[33129] = 25'b0101110011011000100100001;
    rom[33130] = 25'b0101110011010100101001100;
    rom[33131] = 25'b0101110011010000101110010;
    rom[33132] = 25'b0101110011001100110010011;
    rom[33133] = 25'b0101110011001000110101110;
    rom[33134] = 25'b0101110011000100111000100;
    rom[33135] = 25'b0101110011000000111010101;
    rom[33136] = 25'b0101110010111100111100000;
    rom[33137] = 25'b0101110010111000111100110;
    rom[33138] = 25'b0101110010110100111100111;
    rom[33139] = 25'b0101110010110000111100010;
    rom[33140] = 25'b0101110010101100111011000;
    rom[33141] = 25'b0101110010101000111001001;
    rom[33142] = 25'b0101110010100100110110100;
    rom[33143] = 25'b0101110010100000110011010;
    rom[33144] = 25'b0101110010011100101111011;
    rom[33145] = 25'b0101110010011000101010111;
    rom[33146] = 25'b0101110010010100100101101;
    rom[33147] = 25'b0101110010010000011111110;
    rom[33148] = 25'b0101110010001100011001001;
    rom[33149] = 25'b0101110010001000010001111;
    rom[33150] = 25'b0101110010000100001010000;
    rom[33151] = 25'b0101110010000000000001100;
    rom[33152] = 25'b0101110001111011111000010;
    rom[33153] = 25'b0101110001110111101110011;
    rom[33154] = 25'b0101110001110011100011111;
    rom[33155] = 25'b0101110001101111011000101;
    rom[33156] = 25'b0101110001101011001100110;
    rom[33157] = 25'b0101110001100111000000010;
    rom[33158] = 25'b0101110001100010110011000;
    rom[33159] = 25'b0101110001011110100101010;
    rom[33160] = 25'b0101110001011010010110101;
    rom[33161] = 25'b0101110001010110000111100;
    rom[33162] = 25'b0101110001010001110111101;
    rom[33163] = 25'b0101110001001101100111010;
    rom[33164] = 25'b0101110001001001010110000;
    rom[33165] = 25'b0101110001000101000100010;
    rom[33166] = 25'b0101110001000000110001110;
    rom[33167] = 25'b0101110000111100011110101;
    rom[33168] = 25'b0101110000111000001010110;
    rom[33169] = 25'b0101110000110011110110011;
    rom[33170] = 25'b0101110000101111100001010;
    rom[33171] = 25'b0101110000101011001011100;
    rom[33172] = 25'b0101110000100110110101001;
    rom[33173] = 25'b0101110000100010011110000;
    rom[33174] = 25'b0101110000011110000110010;
    rom[33175] = 25'b0101110000011001101101111;
    rom[33176] = 25'b0101110000010101010100110;
    rom[33177] = 25'b0101110000010000111011001;
    rom[33178] = 25'b0101110000001100100000101;
    rom[33179] = 25'b0101110000001000000101101;
    rom[33180] = 25'b0101110000000011101010000;
    rom[33181] = 25'b0101101111111111001101101;
    rom[33182] = 25'b0101101111111010110000101;
    rom[33183] = 25'b0101101111110110010011000;
    rom[33184] = 25'b0101101111110001110100101;
    rom[33185] = 25'b0101101111101101010101101;
    rom[33186] = 25'b0101101111101000110110001;
    rom[33187] = 25'b0101101111100100010101110;
    rom[33188] = 25'b0101101111011111110100111;
    rom[33189] = 25'b0101101111011011010011010;
    rom[33190] = 25'b0101101111010110110001000;
    rom[33191] = 25'b0101101111010010001110001;
    rom[33192] = 25'b0101101111001101101010101;
    rom[33193] = 25'b0101101111001001000110011;
    rom[33194] = 25'b0101101111000100100001100;
    rom[33195] = 25'b0101101110111111111100000;
    rom[33196] = 25'b0101101110111011010101111;
    rom[33197] = 25'b0101101110110110101111000;
    rom[33198] = 25'b0101101110110010000111101;
    rom[33199] = 25'b0101101110101101011111100;
    rom[33200] = 25'b0101101110101000110110110;
    rom[33201] = 25'b0101101110100100001101010;
    rom[33202] = 25'b0101101110011111100011001;
    rom[33203] = 25'b0101101110011010111000100;
    rom[33204] = 25'b0101101110010110001101001;
    rom[33205] = 25'b0101101110010001100001001;
    rom[33206] = 25'b0101101110001100110100100;
    rom[33207] = 25'b0101101110001000000111001;
    rom[33208] = 25'b0101101110000011011001001;
    rom[33209] = 25'b0101101101111110101010100;
    rom[33210] = 25'b0101101101111001111011010;
    rom[33211] = 25'b0101101101110101001011010;
    rom[33212] = 25'b0101101101110000011010110;
    rom[33213] = 25'b0101101101101011101001100;
    rom[33214] = 25'b0101101101100110110111101;
    rom[33215] = 25'b0101101101100010000101001;
    rom[33216] = 25'b0101101101011101010010000;
    rom[33217] = 25'b0101101101011000011110010;
    rom[33218] = 25'b0101101101010011101001110;
    rom[33219] = 25'b0101101101001110110100101;
    rom[33220] = 25'b0101101101001001111110111;
    rom[33221] = 25'b0101101101000101001000100;
    rom[33222] = 25'b0101101101000000010001100;
    rom[33223] = 25'b0101101100111011011001110;
    rom[33224] = 25'b0101101100110110100001011;
    rom[33225] = 25'b0101101100110001101000011;
    rom[33226] = 25'b0101101100101100101110111;
    rom[33227] = 25'b0101101100100111110100100;
    rom[33228] = 25'b0101101100100010111001101;
    rom[33229] = 25'b0101101100011101111110000;
    rom[33230] = 25'b0101101100011001000001111;
    rom[33231] = 25'b0101101100010100000101000;
    rom[33232] = 25'b0101101100001111000111100;
    rom[33233] = 25'b0101101100001010001001011;
    rom[33234] = 25'b0101101100000101001010101;
    rom[33235] = 25'b0101101100000000001011001;
    rom[33236] = 25'b0101101011111011001011001;
    rom[33237] = 25'b0101101011110110001010011;
    rom[33238] = 25'b0101101011110001001001001;
    rom[33239] = 25'b0101101011101100000111001;
    rom[33240] = 25'b0101101011100111000100100;
    rom[33241] = 25'b0101101011100010000001010;
    rom[33242] = 25'b0101101011011100111101010;
    rom[33243] = 25'b0101101011010111111000110;
    rom[33244] = 25'b0101101011010010110011101;
    rom[33245] = 25'b0101101011001101101101110;
    rom[33246] = 25'b0101101011001000100111010;
    rom[33247] = 25'b0101101011000011100000001;
    rom[33248] = 25'b0101101010111110011000011;
    rom[33249] = 25'b0101101010111001010000000;
    rom[33250] = 25'b0101101010110100000111000;
    rom[33251] = 25'b0101101010101110111101011;
    rom[33252] = 25'b0101101010101001110011000;
    rom[33253] = 25'b0101101010100100101000000;
    rom[33254] = 25'b0101101010011111011100100;
    rom[33255] = 25'b0101101010011010010000010;
    rom[33256] = 25'b0101101010010101000011011;
    rom[33257] = 25'b0101101010001111110110000;
    rom[33258] = 25'b0101101010001010100111110;
    rom[33259] = 25'b0101101010000101011001000;
    rom[33260] = 25'b0101101010000000001001101;
    rom[33261] = 25'b0101101001111010111001101;
    rom[33262] = 25'b0101101001110101101001000;
    rom[33263] = 25'b0101101001110000010111101;
    rom[33264] = 25'b0101101001101011000101110;
    rom[33265] = 25'b0101101001100101110011010;
    rom[33266] = 25'b0101101001100000011111111;
    rom[33267] = 25'b0101101001011011001100001;
    rom[33268] = 25'b0101101001010101110111101;
    rom[33269] = 25'b0101101001010000100010100;
    rom[33270] = 25'b0101101001001011001100110;
    rom[33271] = 25'b0101101001000101110110011;
    rom[33272] = 25'b0101101001000000011111011;
    rom[33273] = 25'b0101101000111011000111110;
    rom[33274] = 25'b0101101000110101101111100;
    rom[33275] = 25'b0101101000110000010110101;
    rom[33276] = 25'b0101101000101010111101001;
    rom[33277] = 25'b0101101000100101100010111;
    rom[33278] = 25'b0101101000100000001000000;
    rom[33279] = 25'b0101101000011010101100101;
    rom[33280] = 25'b0101101000010101010000101;
    rom[33281] = 25'b0101101000001111110011111;
    rom[33282] = 25'b0101101000001010010110101;
    rom[33283] = 25'b0101101000000100111000110;
    rom[33284] = 25'b0101100111111111011010001;
    rom[33285] = 25'b0101100111111001111010111;
    rom[33286] = 25'b0101100111110100011011000;
    rom[33287] = 25'b0101100111101110111010101;
    rom[33288] = 25'b0101100111101001011001100;
    rom[33289] = 25'b0101100111100011110111111;
    rom[33290] = 25'b0101100111011110010101011;
    rom[33291] = 25'b0101100111011000110010100;
    rom[33292] = 25'b0101100111010011001110111;
    rom[33293] = 25'b0101100111001101101010101;
    rom[33294] = 25'b0101100111001000000101111;
    rom[33295] = 25'b0101100111000010100000011;
    rom[33296] = 25'b0101100110111100111010010;
    rom[33297] = 25'b0101100110110111010011100;
    rom[33298] = 25'b0101100110110001101100001;
    rom[33299] = 25'b0101100110101100000100010;
    rom[33300] = 25'b0101100110100110011011101;
    rom[33301] = 25'b0101100110100000110010011;
    rom[33302] = 25'b0101100110011011001000101;
    rom[33303] = 25'b0101100110010101011110000;
    rom[33304] = 25'b0101100110001111110011000;
    rom[33305] = 25'b0101100110001010000111010;
    rom[33306] = 25'b0101100110000100011010111;
    rom[33307] = 25'b0101100101111110101110000;
    rom[33308] = 25'b0101100101111001000000011;
    rom[33309] = 25'b0101100101110011010010001;
    rom[33310] = 25'b0101100101101101100011011;
    rom[33311] = 25'b0101100101100111110011111;
    rom[33312] = 25'b0101100101100010000011111;
    rom[33313] = 25'b0101100101011100010011001;
    rom[33314] = 25'b0101100101010110100001111;
    rom[33315] = 25'b0101100101010000101111111;
    rom[33316] = 25'b0101100101001010111101011;
    rom[33317] = 25'b0101100101000101001010010;
    rom[33318] = 25'b0101100100111111010110011;
    rom[33319] = 25'b0101100100111001100010000;
    rom[33320] = 25'b0101100100110011101101000;
    rom[33321] = 25'b0101100100101101110111011;
    rom[33322] = 25'b0101100100101000000001001;
    rom[33323] = 25'b0101100100100010001010010;
    rom[33324] = 25'b0101100100011100010010110;
    rom[33325] = 25'b0101100100010110011010101;
    rom[33326] = 25'b0101100100010000100001111;
    rom[33327] = 25'b0101100100001010101000100;
    rom[33328] = 25'b0101100100000100101110101;
    rom[33329] = 25'b0101100011111110110100001;
    rom[33330] = 25'b0101100011111000111000111;
    rom[33331] = 25'b0101100011110010111101001;
    rom[33332] = 25'b0101100011101101000000110;
    rom[33333] = 25'b0101100011100111000011101;
    rom[33334] = 25'b0101100011100001000110000;
    rom[33335] = 25'b0101100011011011000111110;
    rom[33336] = 25'b0101100011010101001000111;
    rom[33337] = 25'b0101100011001111001001100;
    rom[33338] = 25'b0101100011001001001001011;
    rom[33339] = 25'b0101100011000011001000101;
    rom[33340] = 25'b0101100010111101000111010;
    rom[33341] = 25'b0101100010110111000101011;
    rom[33342] = 25'b0101100010110001000010110;
    rom[33343] = 25'b0101100010101010111111101;
    rom[33344] = 25'b0101100010100100111100000;
    rom[33345] = 25'b0101100010011110110111100;
    rom[33346] = 25'b0101100010011000110010101;
    rom[33347] = 25'b0101100010010010101101000;
    rom[33348] = 25'b0101100010001100100110110;
    rom[33349] = 25'b0101100010000110100000000;
    rom[33350] = 25'b0101100010000000011000100;
    rom[33351] = 25'b0101100001111010010000100;
    rom[33352] = 25'b0101100001110100000111111;
    rom[33353] = 25'b0101100001101101111110101;
    rom[33354] = 25'b0101100001100111110100110;
    rom[33355] = 25'b0101100001100001101010011;
    rom[33356] = 25'b0101100001011011011111010;
    rom[33357] = 25'b0101100001010101010011101;
    rom[33358] = 25'b0101100001001111000111010;
    rom[33359] = 25'b0101100001001000111010011;
    rom[33360] = 25'b0101100001000010101101000;
    rom[33361] = 25'b0101100000111100011110111;
    rom[33362] = 25'b0101100000110110010000001;
    rom[33363] = 25'b0101100000110000000000111;
    rom[33364] = 25'b0101100000101001110001000;
    rom[33365] = 25'b0101100000100011100000011;
    rom[33366] = 25'b0101100000011101001111011;
    rom[33367] = 25'b0101100000010110111101101;
    rom[33368] = 25'b0101100000010000101011010;
    rom[33369] = 25'b0101100000001010011000011;
    rom[33370] = 25'b0101100000000100000100111;
    rom[33371] = 25'b0101011111111101110000110;
    rom[33372] = 25'b0101011111110111011100000;
    rom[33373] = 25'b0101011111110001000110101;
    rom[33374] = 25'b0101011111101010110000110;
    rom[33375] = 25'b0101011111100100011010010;
    rom[33376] = 25'b0101011111011110000011001;
    rom[33377] = 25'b0101011111010111101011011;
    rom[33378] = 25'b0101011111010001010011001;
    rom[33379] = 25'b0101011111001010111010001;
    rom[33380] = 25'b0101011111000100100000101;
    rom[33381] = 25'b0101011110111110000110100;
    rom[33382] = 25'b0101011110110111101011110;
    rom[33383] = 25'b0101011110110001010000011;
    rom[33384] = 25'b0101011110101010110100101;
    rom[33385] = 25'b0101011110100100011000000;
    rom[33386] = 25'b0101011110011101111010111;
    rom[33387] = 25'b0101011110010111011101010;
    rom[33388] = 25'b0101011110010000111110111;
    rom[33389] = 25'b0101011110001010100000000;
    rom[33390] = 25'b0101011110000100000000100;
    rom[33391] = 25'b0101011101111101100000011;
    rom[33392] = 25'b0101011101110110111111110;
    rom[33393] = 25'b0101011101110000011110100;
    rom[33394] = 25'b0101011101101001111100101;
    rom[33395] = 25'b0101011101100011011010001;
    rom[33396] = 25'b0101011101011100110111001;
    rom[33397] = 25'b0101011101010110010011011;
    rom[33398] = 25'b0101011101001111101111001;
    rom[33399] = 25'b0101011101001001001010011;
    rom[33400] = 25'b0101011101000010100100111;
    rom[33401] = 25'b0101011100111011111110111;
    rom[33402] = 25'b0101011100110101011000011;
    rom[33403] = 25'b0101011100101110110001001;
    rom[33404] = 25'b0101011100101000001001010;
    rom[33405] = 25'b0101011100100001100001000;
    rom[33406] = 25'b0101011100011010111000000;
    rom[33407] = 25'b0101011100010100001110100;
    rom[33408] = 25'b0101011100001101100100010;
    rom[33409] = 25'b0101011100000110111001101;
    rom[33410] = 25'b0101011100000000001110010;
    rom[33411] = 25'b0101011011111001100010011;
    rom[33412] = 25'b0101011011110010110101110;
    rom[33413] = 25'b0101011011101100001000110;
    rom[33414] = 25'b0101011011100101011011001;
    rom[33415] = 25'b0101011011011110101100110;
    rom[33416] = 25'b0101011011010111111110000;
    rom[33417] = 25'b0101011011010001001110100;
    rom[33418] = 25'b0101011011001010011110100;
    rom[33419] = 25'b0101011011000011101101111;
    rom[33420] = 25'b0101011010111100111100110;
    rom[33421] = 25'b0101011010110110001010111;
    rom[33422] = 25'b0101011010101111011000101;
    rom[33423] = 25'b0101011010101000100101101;
    rom[33424] = 25'b0101011010100001110010001;
    rom[33425] = 25'b0101011010011010111110000;
    rom[33426] = 25'b0101011010010100001001011;
    rom[33427] = 25'b0101011010001101010100001;
    rom[33428] = 25'b0101011010000110011110010;
    rom[33429] = 25'b0101011001111111100111111;
    rom[33430] = 25'b0101011001111000110000111;
    rom[33431] = 25'b0101011001110001111001001;
    rom[33432] = 25'b0101011001101011000001000;
    rom[33433] = 25'b0101011001100100001000010;
    rom[33434] = 25'b0101011001011101001110111;
    rom[33435] = 25'b0101011001010110010101000;
    rom[33436] = 25'b0101011001001111011010100;
    rom[33437] = 25'b0101011001001000011111100;
    rom[33438] = 25'b0101011001000001100011110;
    rom[33439] = 25'b0101011000111010100111101;
    rom[33440] = 25'b0101011000110011101010110;
    rom[33441] = 25'b0101011000101100101101011;
    rom[33442] = 25'b0101011000100101101111100;
    rom[33443] = 25'b0101011000011110110000111;
    rom[33444] = 25'b0101011000010111110001110;
    rom[33445] = 25'b0101011000010000110010001;
    rom[33446] = 25'b0101011000001001110001111;
    rom[33447] = 25'b0101011000000010110001000;
    rom[33448] = 25'b0101010111111011101111101;
    rom[33449] = 25'b0101010111110100101101101;
    rom[33450] = 25'b0101010111101101101011001;
    rom[33451] = 25'b0101010111100110100111111;
    rom[33452] = 25'b0101010111011111100100010;
    rom[33453] = 25'b0101010111011000100000000;
    rom[33454] = 25'b0101010111010001011011001;
    rom[33455] = 25'b0101010111001010010101110;
    rom[33456] = 25'b0101010111000011001111101;
    rom[33457] = 25'b0101010110111100001001001;
    rom[33458] = 25'b0101010110110101000010000;
    rom[33459] = 25'b0101010110101101111010011;
    rom[33460] = 25'b0101010110100110110010000;
    rom[33461] = 25'b0101010110011111101001010;
    rom[33462] = 25'b0101010110011000011111110;
    rom[33463] = 25'b0101010110010001010101111;
    rom[33464] = 25'b0101010110001010001011010;
    rom[33465] = 25'b0101010110000011000000001;
    rom[33466] = 25'b0101010101111011110100100;
    rom[33467] = 25'b0101010101110100101000001;
    rom[33468] = 25'b0101010101101101011011011;
    rom[33469] = 25'b0101010101100110001110000;
    rom[33470] = 25'b0101010101011111000000001;
    rom[33471] = 25'b0101010101010111110001100;
    rom[33472] = 25'b0101010101010000100010011;
    rom[33473] = 25'b0101010101001001010010111;
    rom[33474] = 25'b0101010101000010000010101;
    rom[33475] = 25'b0101010100111010110001111;
    rom[33476] = 25'b0101010100110011100000100;
    rom[33477] = 25'b0101010100101100001110101;
    rom[33478] = 25'b0101010100100100111100001;
    rom[33479] = 25'b0101010100011101101001001;
    rom[33480] = 25'b0101010100010110010101100;
    rom[33481] = 25'b0101010100001111000001011;
    rom[33482] = 25'b0101010100000111101100101;
    rom[33483] = 25'b0101010100000000010111011;
    rom[33484] = 25'b0101010011111001000001100;
    rom[33485] = 25'b0101010011110001101011001;
    rom[33486] = 25'b0101010011101010010100010;
    rom[33487] = 25'b0101010011100010111100101;
    rom[33488] = 25'b0101010011011011100100100;
    rom[33489] = 25'b0101010011010100001011111;
    rom[33490] = 25'b0101010011001100110010110;
    rom[33491] = 25'b0101010011000101011001000;
    rom[33492] = 25'b0101010010111101111110101;
    rom[33493] = 25'b0101010010110110100011111;
    rom[33494] = 25'b0101010010101111001000011;
    rom[33495] = 25'b0101010010100111101100011;
    rom[33496] = 25'b0101010010100000001111111;
    rom[33497] = 25'b0101010010011000110010110;
    rom[33498] = 25'b0101010010010001010101001;
    rom[33499] = 25'b0101010010001001110111000;
    rom[33500] = 25'b0101010010000010011000001;
    rom[33501] = 25'b0101010001111010111000111;
    rom[33502] = 25'b0101010001110011011001000;
    rom[33503] = 25'b0101010001101011111000101;
    rom[33504] = 25'b0101010001100100010111101;
    rom[33505] = 25'b0101010001011100110110001;
    rom[33506] = 25'b0101010001010101010100000;
    rom[33507] = 25'b0101010001001101110001011;
    rom[33508] = 25'b0101010001000110001110010;
    rom[33509] = 25'b0101010000111110101010100;
    rom[33510] = 25'b0101010000110111000110010;
    rom[33511] = 25'b0101010000101111100001011;
    rom[33512] = 25'b0101010000100111111100000;
    rom[33513] = 25'b0101010000100000010110001;
    rom[33514] = 25'b0101010000011000101111101;
    rom[33515] = 25'b0101010000010001001000101;
    rom[33516] = 25'b0101010000001001100001000;
    rom[33517] = 25'b0101010000000001111000111;
    rom[33518] = 25'b0101001111111010010000010;
    rom[33519] = 25'b0101001111110010100111000;
    rom[33520] = 25'b0101001111101010111101010;
    rom[33521] = 25'b0101001111100011010010111;
    rom[33522] = 25'b0101001111011011101000000;
    rom[33523] = 25'b0101001111010011111100101;
    rom[33524] = 25'b0101001111001100010000110;
    rom[33525] = 25'b0101001111000100100100010;
    rom[33526] = 25'b0101001110111100110111001;
    rom[33527] = 25'b0101001110110101001001101;
    rom[33528] = 25'b0101001110101101011011100;
    rom[33529] = 25'b0101001110100101101100111;
    rom[33530] = 25'b0101001110011101111101101;
    rom[33531] = 25'b0101001110010110001101111;
    rom[33532] = 25'b0101001110001110011101101;
    rom[33533] = 25'b0101001110000110101100111;
    rom[33534] = 25'b0101001101111110111011100;
    rom[33535] = 25'b0101001101110111001001100;
    rom[33536] = 25'b0101001101101111010111000;
    rom[33537] = 25'b0101001101100111100100000;
    rom[33538] = 25'b0101001101011111110000100;
    rom[33539] = 25'b0101001101010111111100100;
    rom[33540] = 25'b0101001101010000000111111;
    rom[33541] = 25'b0101001101001000010010110;
    rom[33542] = 25'b0101001101000000011101001;
    rom[33543] = 25'b0101001100111000100110111;
    rom[33544] = 25'b0101001100110000110000001;
    rom[33545] = 25'b0101001100101000111000110;
    rom[33546] = 25'b0101001100100001000001000;
    rom[33547] = 25'b0101001100011001001000101;
    rom[33548] = 25'b0101001100010001001111110;
    rom[33549] = 25'b0101001100001001010110010;
    rom[33550] = 25'b0101001100000001011100010;
    rom[33551] = 25'b0101001011111001100001111;
    rom[33552] = 25'b0101001011110001100110110;
    rom[33553] = 25'b0101001011101001101011001;
    rom[33554] = 25'b0101001011100001101111001;
    rom[33555] = 25'b0101001011011001110010100;
    rom[33556] = 25'b0101001011010001110101011;
    rom[33557] = 25'b0101001011001001110111101;
    rom[33558] = 25'b0101001011000001111001011;
    rom[33559] = 25'b0101001010111001111010101;
    rom[33560] = 25'b0101001010110001111011011;
    rom[33561] = 25'b0101001010101001111011101;
    rom[33562] = 25'b0101001010100001111011010;
    rom[33563] = 25'b0101001010011001111010011;
    rom[33564] = 25'b0101001010010001111000111;
    rom[33565] = 25'b0101001010001001110111000;
    rom[33566] = 25'b0101001010000001110100100;
    rom[33567] = 25'b0101001001111001110001101;
    rom[33568] = 25'b0101001001110001101110000;
    rom[33569] = 25'b0101001001101001101010001;
    rom[33570] = 25'b0101001001100001100101100;
    rom[33571] = 25'b0101001001011001100000011;
    rom[33572] = 25'b0101001001010001011010110;
    rom[33573] = 25'b0101001001001001010100101;
    rom[33574] = 25'b0101001001000001001101111;
    rom[33575] = 25'b0101001000111001000110110;
    rom[33576] = 25'b0101001000110000111111001;
    rom[33577] = 25'b0101001000101000110110111;
    rom[33578] = 25'b0101001000100000101110001;
    rom[33579] = 25'b0101001000011000100100111;
    rom[33580] = 25'b0101001000010000011011001;
    rom[33581] = 25'b0101001000001000010000110;
    rom[33582] = 25'b0101001000000000000101111;
    rom[33583] = 25'b0101000111110111111010100;
    rom[33584] = 25'b0101000111101111101110101;
    rom[33585] = 25'b0101000111100111100010010;
    rom[33586] = 25'b0101000111011111010101011;
    rom[33587] = 25'b0101000111010111001000000;
    rom[33588] = 25'b0101000111001110111010000;
    rom[33589] = 25'b0101000111000110101011100;
    rom[33590] = 25'b0101000110111110011100100;
    rom[33591] = 25'b0101000110110110001101000;
    rom[33592] = 25'b0101000110101101111101000;
    rom[33593] = 25'b0101000110100101101100100;
    rom[33594] = 25'b0101000110011101011011011;
    rom[33595] = 25'b0101000110010101001001111;
    rom[33596] = 25'b0101000110001100110111110;
    rom[33597] = 25'b0101000110000100100101001;
    rom[33598] = 25'b0101000101111100010010000;
    rom[33599] = 25'b0101000101110011111110011;
    rom[33600] = 25'b0101000101101011101010010;
    rom[33601] = 25'b0101000101100011010101110;
    rom[33602] = 25'b0101000101011011000000100;
    rom[33603] = 25'b0101000101010010101010111;
    rom[33604] = 25'b0101000101001010010100101;
    rom[33605] = 25'b0101000101000001111101111;
    rom[33606] = 25'b0101000100111001100110110;
    rom[33607] = 25'b0101000100110001001111000;
    rom[33608] = 25'b0101000100101000110110111;
    rom[33609] = 25'b0101000100100000011110000;
    rom[33610] = 25'b0101000100011000000100111;
    rom[33611] = 25'b0101000100001111101011001;
    rom[33612] = 25'b0101000100000111010000111;
    rom[33613] = 25'b0101000011111110110110001;
    rom[33614] = 25'b0101000011110110011010111;
    rom[33615] = 25'b0101000011101101111111000;
    rom[33616] = 25'b0101000011100101100010110;
    rom[33617] = 25'b0101000011011101000110000;
    rom[33618] = 25'b0101000011010100101000110;
    rom[33619] = 25'b0101000011001100001010111;
    rom[33620] = 25'b0101000011000011101100101;
    rom[33621] = 25'b0101000010111011001101111;
    rom[33622] = 25'b0101000010110010101110100;
    rom[33623] = 25'b0101000010101010001110110;
    rom[33624] = 25'b0101000010100001101110011;
    rom[33625] = 25'b0101000010011001001101100;
    rom[33626] = 25'b0101000010010000101100010;
    rom[33627] = 25'b0101000010001000001010100;
    rom[33628] = 25'b0101000001111111101000001;
    rom[33629] = 25'b0101000001110111000101010;
    rom[33630] = 25'b0101000001101110100010000;
    rom[33631] = 25'b0101000001100101111110001;
    rom[33632] = 25'b0101000001011101011001111;
    rom[33633] = 25'b0101000001010100110101000;
    rom[33634] = 25'b0101000001001100001111110;
    rom[33635] = 25'b0101000001000011101010000;
    rom[33636] = 25'b0101000000111011000011101;
    rom[33637] = 25'b0101000000110010011100111;
    rom[33638] = 25'b0101000000101001110101101;
    rom[33639] = 25'b0101000000100001001101110;
    rom[33640] = 25'b0101000000011000100101100;
    rom[33641] = 25'b0101000000001111111100110;
    rom[33642] = 25'b0101000000000111010011100;
    rom[33643] = 25'b0100111111111110101001110;
    rom[33644] = 25'b0100111111110101111111100;
    rom[33645] = 25'b0100111111101101010100101;
    rom[33646] = 25'b0100111111100100101001100;
    rom[33647] = 25'b0100111111011011111101110;
    rom[33648] = 25'b0100111111010011010001100;
    rom[33649] = 25'b0100111111001010100100110;
    rom[33650] = 25'b0100111111000001110111101;
    rom[33651] = 25'b0100111110111001001001111;
    rom[33652] = 25'b0100111110110000011011110;
    rom[33653] = 25'b0100111110100111101101000;
    rom[33654] = 25'b0100111110011110111101111;
    rom[33655] = 25'b0100111110010110001110001;
    rom[33656] = 25'b0100111110001101011110000;
    rom[33657] = 25'b0100111110000100101101011;
    rom[33658] = 25'b0100111101111011111100010;
    rom[33659] = 25'b0100111101110011001010101;
    rom[33660] = 25'b0100111101101010011000100;
    rom[33661] = 25'b0100111101100001100110000;
    rom[33662] = 25'b0100111101011000110011000;
    rom[33663] = 25'b0100111101001111111111011;
    rom[33664] = 25'b0100111101000111001011011;
    rom[33665] = 25'b0100111100111110010110111;
    rom[33666] = 25'b0100111100110101100001111;
    rom[33667] = 25'b0100111100101100101100011;
    rom[33668] = 25'b0100111100100011110110011;
    rom[33669] = 25'b0100111100011011000000000;
    rom[33670] = 25'b0100111100010010001001001;
    rom[33671] = 25'b0100111100001001010001101;
    rom[33672] = 25'b0100111100000000011001110;
    rom[33673] = 25'b0100111011110111100001011;
    rom[33674] = 25'b0100111011101110101000101;
    rom[33675] = 25'b0100111011100101101111010;
    rom[33676] = 25'b0100111011011100110101100;
    rom[33677] = 25'b0100111011010011111011010;
    rom[33678] = 25'b0100111011001011000000100;
    rom[33679] = 25'b0100111011000010000101010;
    rom[33680] = 25'b0100111010111001001001100;
    rom[33681] = 25'b0100111010110000001101010;
    rom[33682] = 25'b0100111010100111010000101;
    rom[33683] = 25'b0100111010011110010011100;
    rom[33684] = 25'b0100111010010101010101111;
    rom[33685] = 25'b0100111010001100010111110;
    rom[33686] = 25'b0100111010000011011001010;
    rom[33687] = 25'b0100111001111010011010010;
    rom[33688] = 25'b0100111001110001011010101;
    rom[33689] = 25'b0100111001101000011010110;
    rom[33690] = 25'b0100111001011111011010010;
    rom[33691] = 25'b0100111001010110011001011;
    rom[33692] = 25'b0100111001001101011000000;
    rom[33693] = 25'b0100111001000100010110001;
    rom[33694] = 25'b0100111000111011010011110;
    rom[33695] = 25'b0100111000110010010001000;
    rom[33696] = 25'b0100111000101001001101110;
    rom[33697] = 25'b0100111000100000001010000;
    rom[33698] = 25'b0100111000010111000101110;
    rom[33699] = 25'b0100111000001110000001000;
    rom[33700] = 25'b0100111000000100111011111;
    rom[33701] = 25'b0100110111111011110110010;
    rom[33702] = 25'b0100110111110010110000010;
    rom[33703] = 25'b0100110111101001101001110;
    rom[33704] = 25'b0100110111100000100010110;
    rom[33705] = 25'b0100110111010111011011010;
    rom[33706] = 25'b0100110111001110010011011;
    rom[33707] = 25'b0100110111000101001010111;
    rom[33708] = 25'b0100110110111100000010000;
    rom[33709] = 25'b0100110110110010111000110;
    rom[33710] = 25'b0100110110101001101111000;
    rom[33711] = 25'b0100110110100000100100101;
    rom[33712] = 25'b0100110110010111011010000;
    rom[33713] = 25'b0100110110001110001110110;
    rom[33714] = 25'b0100110110000101000011010;
    rom[33715] = 25'b0100110101111011110111000;
    rom[33716] = 25'b0100110101110010101010100;
    rom[33717] = 25'b0100110101101001011101100;
    rom[33718] = 25'b0100110101100000010000001;
    rom[33719] = 25'b0100110101010111000010001;
    rom[33720] = 25'b0100110101001101110011110;
    rom[33721] = 25'b0100110101000100100100111;
    rom[33722] = 25'b0100110100111011010101100;
    rom[33723] = 25'b0100110100110010000101110;
    rom[33724] = 25'b0100110100101000110101101;
    rom[33725] = 25'b0100110100011111100101000;
    rom[33726] = 25'b0100110100010110010011110;
    rom[33727] = 25'b0100110100001101000010010;
    rom[33728] = 25'b0100110100000011110000001;
    rom[33729] = 25'b0100110011111010011101110;
    rom[33730] = 25'b0100110011110001001010110;
    rom[33731] = 25'b0100110011100111110111011;
    rom[33732] = 25'b0100110011011110100011100;
    rom[33733] = 25'b0100110011010101001111010;
    rom[33734] = 25'b0100110011001011111010100;
    rom[33735] = 25'b0100110011000010100101011;
    rom[33736] = 25'b0100110010111001001111101;
    rom[33737] = 25'b0100110010101111111001101;
    rom[33738] = 25'b0100110010100110100011001;
    rom[33739] = 25'b0100110010011101001100001;
    rom[33740] = 25'b0100110010010011110100101;
    rom[33741] = 25'b0100110010001010011100110;
    rom[33742] = 25'b0100110010000001000100011;
    rom[33743] = 25'b0100110001110111101011101;
    rom[33744] = 25'b0100110001101110010010011;
    rom[33745] = 25'b0100110001100100111000110;
    rom[33746] = 25'b0100110001011011011110101;
    rom[33747] = 25'b0100110001010010000100000;
    rom[33748] = 25'b0100110001001000101001000;
    rom[33749] = 25'b0100110000111111001101101;
    rom[33750] = 25'b0100110000110101110001101;
    rom[33751] = 25'b0100110000101100010101011;
    rom[33752] = 25'b0100110000100010111000101;
    rom[33753] = 25'b0100110000011001011011011;
    rom[33754] = 25'b0100110000001111111101110;
    rom[33755] = 25'b0100110000000110011111101;
    rom[33756] = 25'b0100101111111101000001001;
    rom[33757] = 25'b0100101111110011100010001;
    rom[33758] = 25'b0100101111101010000010101;
    rom[33759] = 25'b0100101111100000100010111;
    rom[33760] = 25'b0100101111010111000010100;
    rom[33761] = 25'b0100101111001101100001110;
    rom[33762] = 25'b0100101111000100000000101;
    rom[33763] = 25'b0100101110111010011111000;
    rom[33764] = 25'b0100101110110000111101000;
    rom[33765] = 25'b0100101110100111011010100;
    rom[33766] = 25'b0100101110011101110111101;
    rom[33767] = 25'b0100101110010100010100010;
    rom[33768] = 25'b0100101110001010110000011;
    rom[33769] = 25'b0100101110000001001100010;
    rom[33770] = 25'b0100101101110111100111100;
    rom[33771] = 25'b0100101101101110000010100;
    rom[33772] = 25'b0100101101100100011101000;
    rom[33773] = 25'b0100101101011010110111001;
    rom[33774] = 25'b0100101101010001010000110;
    rom[33775] = 25'b0100101101000111101001111;
    rom[33776] = 25'b0100101100111110000010101;
    rom[33777] = 25'b0100101100110100011011000;
    rom[33778] = 25'b0100101100101010110010111;
    rom[33779] = 25'b0100101100100001001010011;
    rom[33780] = 25'b0100101100010111100001011;
    rom[33781] = 25'b0100101100001101111000000;
    rom[33782] = 25'b0100101100000100001110010;
    rom[33783] = 25'b0100101011111010100100000;
    rom[33784] = 25'b0100101011110000111001011;
    rom[33785] = 25'b0100101011100111001110010;
    rom[33786] = 25'b0100101011011101100010110;
    rom[33787] = 25'b0100101011010011110110110;
    rom[33788] = 25'b0100101011001010001010100;
    rom[33789] = 25'b0100101011000000011101101;
    rom[33790] = 25'b0100101010110110110000011;
    rom[33791] = 25'b0100101010101101000010111;
    rom[33792] = 25'b0100101010100011010100110;
    rom[33793] = 25'b0100101010011001100110010;
    rom[33794] = 25'b0100101010001111110111011;
    rom[33795] = 25'b0100101010000110001000001;
    rom[33796] = 25'b0100101001111100011000010;
    rom[33797] = 25'b0100101001110010101000001;
    rom[33798] = 25'b0100101001101000110111101;
    rom[33799] = 25'b0100101001011111000110100;
    rom[33800] = 25'b0100101001010101010101001;
    rom[33801] = 25'b0100101001001011100011011;
    rom[33802] = 25'b0100101001000001110001001;
    rom[33803] = 25'b0100101000110111111110100;
    rom[33804] = 25'b0100101000101110001011011;
    rom[33805] = 25'b0100101000100100010111111;
    rom[33806] = 25'b0100101000011010100100000;
    rom[33807] = 25'b0100101000010000101111101;
    rom[33808] = 25'b0100101000000110111010111;
    rom[33809] = 25'b0100100111111101000101110;
    rom[33810] = 25'b0100100111110011010000010;
    rom[33811] = 25'b0100100111101001011010010;
    rom[33812] = 25'b0100100111011111100011110;
    rom[33813] = 25'b0100100111010101101101000;
    rom[33814] = 25'b0100100111001011110101111;
    rom[33815] = 25'b0100100111000001111110001;
    rom[33816] = 25'b0100100110111000000110001;
    rom[33817] = 25'b0100100110101110001101110;
    rom[33818] = 25'b0100100110100100010100111;
    rom[33819] = 25'b0100100110011010011011101;
    rom[33820] = 25'b0100100110010000100010000;
    rom[33821] = 25'b0100100110000110100111111;
    rom[33822] = 25'b0100100101111100101101011;
    rom[33823] = 25'b0100100101110010110010100;
    rom[33824] = 25'b0100100101101000110111010;
    rom[33825] = 25'b0100100101011110111011100;
    rom[33826] = 25'b0100100101010100111111011;
    rom[33827] = 25'b0100100101001011000010111;
    rom[33828] = 25'b0100100101000001000110000;
    rom[33829] = 25'b0100100100110111001000101;
    rom[33830] = 25'b0100100100101101001010111;
    rom[33831] = 25'b0100100100100011001100111;
    rom[33832] = 25'b0100100100011001001110011;
    rom[33833] = 25'b0100100100001111001111011;
    rom[33834] = 25'b0100100100000101010000000;
    rom[33835] = 25'b0100100011111011010000011;
    rom[33836] = 25'b0100100011110001010000001;
    rom[33837] = 25'b0100100011100111001111101;
    rom[33838] = 25'b0100100011011101001110110;
    rom[33839] = 25'b0100100011010011001101100;
    rom[33840] = 25'b0100100011001001001011101;
    rom[33841] = 25'b0100100010111111001001101;
    rom[33842] = 25'b0100100010110101000111001;
    rom[33843] = 25'b0100100010101011000100001;
    rom[33844] = 25'b0100100010100001000000111;
    rom[33845] = 25'b0100100010010110111101010;
    rom[33846] = 25'b0100100010001100111001001;
    rom[33847] = 25'b0100100010000010110100101;
    rom[33848] = 25'b0100100001111000101111110;
    rom[33849] = 25'b0100100001101110101010100;
    rom[33850] = 25'b0100100001100100100100111;
    rom[33851] = 25'b0100100001011010011110110;
    rom[33852] = 25'b0100100001010000011000010;
    rom[33853] = 25'b0100100001000110010001100;
    rom[33854] = 25'b0100100000111100001010010;
    rom[33855] = 25'b0100100000110010000010101;
    rom[33856] = 25'b0100100000100111111010101;
    rom[33857] = 25'b0100100000011101110010001;
    rom[33858] = 25'b0100100000010011101001011;
    rom[33859] = 25'b0100100000001001100000010;
    rom[33860] = 25'b0100011111111111010110101;
    rom[33861] = 25'b0100011111110101001100110;
    rom[33862] = 25'b0100011111101011000010100;
    rom[33863] = 25'b0100011111100000110111110;
    rom[33864] = 25'b0100011111010110101100101;
    rom[33865] = 25'b0100011111001100100001001;
    rom[33866] = 25'b0100011111000010010101010;
    rom[33867] = 25'b0100011110111000001001000;
    rom[33868] = 25'b0100011110101101111100011;
    rom[33869] = 25'b0100011110100011101111010;
    rom[33870] = 25'b0100011110011001100010000;
    rom[33871] = 25'b0100011110001111010100001;
    rom[33872] = 25'b0100011110000101000110000;
    rom[33873] = 25'b0100011101111010110111011;
    rom[33874] = 25'b0100011101110000101000100;
    rom[33875] = 25'b0100011101100110011001010;
    rom[33876] = 25'b0100011101011100001001100;
    rom[33877] = 25'b0100011101010001111001100;
    rom[33878] = 25'b0100011101000111101001000;
    rom[33879] = 25'b0100011100111101011000001;
    rom[33880] = 25'b0100011100110011000111000;
    rom[33881] = 25'b0100011100101000110101011;
    rom[33882] = 25'b0100011100011110100011100;
    rom[33883] = 25'b0100011100010100010001001;
    rom[33884] = 25'b0100011100001001111110011;
    rom[33885] = 25'b0100011011111111101011011;
    rom[33886] = 25'b0100011011110101010111111;
    rom[33887] = 25'b0100011011101011000100001;
    rom[33888] = 25'b0100011011100000110000000;
    rom[33889] = 25'b0100011011010110011011011;
    rom[33890] = 25'b0100011011001100000110100;
    rom[33891] = 25'b0100011011000001110001001;
    rom[33892] = 25'b0100011010110111011011011;
    rom[33893] = 25'b0100011010101101000101011;
    rom[33894] = 25'b0100011010100010101111000;
    rom[33895] = 25'b0100011010011000011000010;
    rom[33896] = 25'b0100011010001110000001001;
    rom[33897] = 25'b0100011010000011101001101;
    rom[33898] = 25'b0100011001111001010001110;
    rom[33899] = 25'b0100011001101110111001100;
    rom[33900] = 25'b0100011001100100100000110;
    rom[33901] = 25'b0100011001011010000111111;
    rom[33902] = 25'b0100011001001111101110100;
    rom[33903] = 25'b0100011001000101010100110;
    rom[33904] = 25'b0100011000111010111010110;
    rom[33905] = 25'b0100011000110000100000010;
    rom[33906] = 25'b0100011000100110000101100;
    rom[33907] = 25'b0100011000011011101010010;
    rom[33908] = 25'b0100011000010001001110111;
    rom[33909] = 25'b0100011000000110110010111;
    rom[33910] = 25'b0100010111111100010110101;
    rom[33911] = 25'b0100010111110001111010001;
    rom[33912] = 25'b0100010111100111011101001;
    rom[33913] = 25'b0100010111011100111111110;
    rom[33914] = 25'b0100010111010010100010001;
    rom[33915] = 25'b0100010111001000000100000;
    rom[33916] = 25'b0100010110111101100101101;
    rom[33917] = 25'b0100010110110011000110111;
    rom[33918] = 25'b0100010110101000100111110;
    rom[33919] = 25'b0100010110011110001000010;
    rom[33920] = 25'b0100010110010011101000100;
    rom[33921] = 25'b0100010110001001001000010;
    rom[33922] = 25'b0100010101111110100111110;
    rom[33923] = 25'b0100010101110100000110111;
    rom[33924] = 25'b0100010101101001100101101;
    rom[33925] = 25'b0100010101011111000100000;
    rom[33926] = 25'b0100010101010100100010001;
    rom[33927] = 25'b0100010101001001111111110;
    rom[33928] = 25'b0100010100111111011101001;
    rom[33929] = 25'b0100010100110100111010001;
    rom[33930] = 25'b0100010100101010010110111;
    rom[33931] = 25'b0100010100011111110011001;
    rom[33932] = 25'b0100010100010101001111001;
    rom[33933] = 25'b0100010100001010101010101;
    rom[33934] = 25'b0100010100000000000101111;
    rom[33935] = 25'b0100010011110101100000111;
    rom[33936] = 25'b0100010011101010111011011;
    rom[33937] = 25'b0100010011100000010101101;
    rom[33938] = 25'b0100010011010101101111100;
    rom[33939] = 25'b0100010011001011001001001;
    rom[33940] = 25'b0100010011000000100010010;
    rom[33941] = 25'b0100010010110101111011000;
    rom[33942] = 25'b0100010010101011010011101;
    rom[33943] = 25'b0100010010100000101011110;
    rom[33944] = 25'b0100010010010110000011101;
    rom[33945] = 25'b0100010010001011011011000;
    rom[33946] = 25'b0100010010000000110010001;
    rom[33947] = 25'b0100010001110110001000111;
    rom[33948] = 25'b0100010001101011011111011;
    rom[33949] = 25'b0100010001100000110101100;
    rom[33950] = 25'b0100010001010110001011010;
    rom[33951] = 25'b0100010001001011100000110;
    rom[33952] = 25'b0100010001000000110101110;
    rom[33953] = 25'b0100010000110110001010100;
    rom[33954] = 25'b0100010000101011011111000;
    rom[33955] = 25'b0100010000100000110011000;
    rom[33956] = 25'b0100010000010110000110110;
    rom[33957] = 25'b0100010000001011011010010;
    rom[33958] = 25'b0100010000000000101101010;
    rom[33959] = 25'b0100001111110110000000000;
    rom[33960] = 25'b0100001111101011010010011;
    rom[33961] = 25'b0100001111100000100100100;
    rom[33962] = 25'b0100001111010101110110010;
    rom[33963] = 25'b0100001111001011000111101;
    rom[33964] = 25'b0100001111000000011000110;
    rom[33965] = 25'b0100001110110101101001100;
    rom[33966] = 25'b0100001110101010111001111;
    rom[33967] = 25'b0100001110100000001010000;
    rom[33968] = 25'b0100001110010101011001110;
    rom[33969] = 25'b0100001110001010101001001;
    rom[33970] = 25'b0100001101111111111000010;
    rom[33971] = 25'b0100001101110101000111001;
    rom[33972] = 25'b0100001101101010010101100;
    rom[33973] = 25'b0100001101011111100011100;
    rom[33974] = 25'b0100001101010100110001011;
    rom[33975] = 25'b0100001101001001111110111;
    rom[33976] = 25'b0100001100111111001100000;
    rom[33977] = 25'b0100001100110100011000110;
    rom[33978] = 25'b0100001100101001100101011;
    rom[33979] = 25'b0100001100011110110001100;
    rom[33980] = 25'b0100001100010011111101011;
    rom[33981] = 25'b0100001100001001001000111;
    rom[33982] = 25'b0100001011111110010100000;
    rom[33983] = 25'b0100001011110011011111000;
    rom[33984] = 25'b0100001011101000101001100;
    rom[33985] = 25'b0100001011011101110011110;
    rom[33986] = 25'b0100001011010010111101110;
    rom[33987] = 25'b0100001011001000000111011;
    rom[33988] = 25'b0100001010111101010000101;
    rom[33989] = 25'b0100001010110010011001101;
    rom[33990] = 25'b0100001010100111100010010;
    rom[33991] = 25'b0100001010011100101010101;
    rom[33992] = 25'b0100001010010001110010101;
    rom[33993] = 25'b0100001010000110111010011;
    rom[33994] = 25'b0100001001111100000001110;
    rom[33995] = 25'b0100001001110001001000110;
    rom[33996] = 25'b0100001001100110001111100;
    rom[33997] = 25'b0100001001011011010110000;
    rom[33998] = 25'b0100001001010000011100001;
    rom[33999] = 25'b0100001001000101100010000;
    rom[34000] = 25'b0100001000111010100111100;
    rom[34001] = 25'b0100001000101111101100110;
    rom[34002] = 25'b0100001000100100110001101;
    rom[34003] = 25'b0100001000011001110110001;
    rom[34004] = 25'b0100001000001110111010100;
    rom[34005] = 25'b0100001000000011111110100;
    rom[34006] = 25'b0100000111111001000010001;
    rom[34007] = 25'b0100000111101110000101100;
    rom[34008] = 25'b0100000111100011001000100;
    rom[34009] = 25'b0100000111011000001011010;
    rom[34010] = 25'b0100000111001101001101101;
    rom[34011] = 25'b0100000111000010001111110;
    rom[34012] = 25'b0100000110110111010001101;
    rom[34013] = 25'b0100000110101100010011001;
    rom[34014] = 25'b0100000110100001010100011;
    rom[34015] = 25'b0100000110010110010101010;
    rom[34016] = 25'b0100000110001011010101111;
    rom[34017] = 25'b0100000110000000010110010;
    rom[34018] = 25'b0100000101110101010110010;
    rom[34019] = 25'b0100000101101010010101111;
    rom[34020] = 25'b0100000101011111010101011;
    rom[34021] = 25'b0100000101010100010100011;
    rom[34022] = 25'b0100000101001001010011010;
    rom[34023] = 25'b0100000100111110010001110;
    rom[34024] = 25'b0100000100110011010000000;
    rom[34025] = 25'b0100000100101000001101111;
    rom[34026] = 25'b0100000100011101001011100;
    rom[34027] = 25'b0100000100010010001000110;
    rom[34028] = 25'b0100000100000111000101110;
    rom[34029] = 25'b0100000011111100000010100;
    rom[34030] = 25'b0100000011110000111111000;
    rom[34031] = 25'b0100000011100101111011001;
    rom[34032] = 25'b0100000011011010110110111;
    rom[34033] = 25'b0100000011001111110010100;
    rom[34034] = 25'b0100000011000100101101110;
    rom[34035] = 25'b0100000010111001101000110;
    rom[34036] = 25'b0100000010101110100011011;
    rom[34037] = 25'b0100000010100011011101110;
    rom[34038] = 25'b0100000010011000010111111;
    rom[34039] = 25'b0100000010001101010001101;
    rom[34040] = 25'b0100000010000010001011001;
    rom[34041] = 25'b0100000001110111000100011;
    rom[34042] = 25'b0100000001101011111101011;
    rom[34043] = 25'b0100000001100000110110000;
    rom[34044] = 25'b0100000001010101101110011;
    rom[34045] = 25'b0100000001001010100110011;
    rom[34046] = 25'b0100000000111111011110010;
    rom[34047] = 25'b0100000000110100010101110;
    rom[34048] = 25'b0100000000101001001101000;
    rom[34049] = 25'b0100000000011110000100000;
    rom[34050] = 25'b0100000000010010111010101;
    rom[34051] = 25'b0100000000000111110000111;
    rom[34052] = 25'b0011111111111100100111000;
    rom[34053] = 25'b0011111111110001011100111;
    rom[34054] = 25'b0011111111100110010010011;
    rom[34055] = 25'b0011111111011011000111101;
    rom[34056] = 25'b0011111111001111111100101;
    rom[34057] = 25'b0011111111000100110001010;
    rom[34058] = 25'b0011111110111001100101110;
    rom[34059] = 25'b0011111110101110011001110;
    rom[34060] = 25'b0011111110100011001101101;
    rom[34061] = 25'b0011111110011000000001010;
    rom[34062] = 25'b0011111110001100110100100;
    rom[34063] = 25'b0011111110000001100111101;
    rom[34064] = 25'b0011111101110110011010010;
    rom[34065] = 25'b0011111101101011001100110;
    rom[34066] = 25'b0011111101011111111111000;
    rom[34067] = 25'b0011111101010100110000111;
    rom[34068] = 25'b0011111101001001100010100;
    rom[34069] = 25'b0011111100111110010011111;
    rom[34070] = 25'b0011111100110011000101000;
    rom[34071] = 25'b0011111100100111110101111;
    rom[34072] = 25'b0011111100011100100110011;
    rom[34073] = 25'b0011111100010001010110110;
    rom[34074] = 25'b0011111100000110000110110;
    rom[34075] = 25'b0011111011111010110110100;
    rom[34076] = 25'b0011111011101111100110000;
    rom[34077] = 25'b0011111011100100010101010;
    rom[34078] = 25'b0011111011011001000100001;
    rom[34079] = 25'b0011111011001101110010111;
    rom[34080] = 25'b0011111011000010100001010;
    rom[34081] = 25'b0011111010110111001111011;
    rom[34082] = 25'b0011111010101011111101010;
    rom[34083] = 25'b0011111010100000101010111;
    rom[34084] = 25'b0011111010010101011000010;
    rom[34085] = 25'b0011111010001010000101010;
    rom[34086] = 25'b0011111001111110110010001;
    rom[34087] = 25'b0011111001110011011110110;
    rom[34088] = 25'b0011111001101000001011000;
    rom[34089] = 25'b0011111001011100110111000;
    rom[34090] = 25'b0011111001010001100010111;
    rom[34091] = 25'b0011111001000110001110011;
    rom[34092] = 25'b0011111000111010111001101;
    rom[34093] = 25'b0011111000101111100100101;
    rom[34094] = 25'b0011111000100100001111011;
    rom[34095] = 25'b0011111000011000111001111;
    rom[34096] = 25'b0011111000001101100100001;
    rom[34097] = 25'b0011111000000010001110000;
    rom[34098] = 25'b0011110111110110110111110;
    rom[34099] = 25'b0011110111101011100001010;
    rom[34100] = 25'b0011110111100000001010100;
    rom[34101] = 25'b0011110111010100110011011;
    rom[34102] = 25'b0011110111001001011100000;
    rom[34103] = 25'b0011110110111110000100101;
    rom[34104] = 25'b0011110110110010101100110;
    rom[34105] = 25'b0011110110100111010100101;
    rom[34106] = 25'b0011110110011011111100011;
    rom[34107] = 25'b0011110110010000100011111;
    rom[34108] = 25'b0011110110000101001011000;
    rom[34109] = 25'b0011110101111001110001111;
    rom[34110] = 25'b0011110101101110011000101;
    rom[34111] = 25'b0011110101100010111111001;
    rom[34112] = 25'b0011110101010111100101010;
    rom[34113] = 25'b0011110101001100001011001;
    rom[34114] = 25'b0011110101000000110000111;
    rom[34115] = 25'b0011110100110101010110010;
    rom[34116] = 25'b0011110100101001111011100;
    rom[34117] = 25'b0011110100011110100000100;
    rom[34118] = 25'b0011110100010011000101010;
    rom[34119] = 25'b0011110100000111101001101;
    rom[34120] = 25'b0011110011111100001101111;
    rom[34121] = 25'b0011110011110000110001111;
    rom[34122] = 25'b0011110011100101010101101;
    rom[34123] = 25'b0011110011011001111001001;
    rom[34124] = 25'b0011110011001110011100011;
    rom[34125] = 25'b0011110011000010111111011;
    rom[34126] = 25'b0011110010110111100010001;
    rom[34127] = 25'b0011110010101100000100101;
    rom[34128] = 25'b0011110010100000100111000;
    rom[34129] = 25'b0011110010010101001001001;
    rom[34130] = 25'b0011110010001001101010111;
    rom[34131] = 25'b0011110001111110001100100;
    rom[34132] = 25'b0011110001110010101101110;
    rom[34133] = 25'b0011110001100111001110111;
    rom[34134] = 25'b0011110001011011101111110;
    rom[34135] = 25'b0011110001010000010000100;
    rom[34136] = 25'b0011110001000100110000111;
    rom[34137] = 25'b0011110000111001010001000;
    rom[34138] = 25'b0011110000101101110001000;
    rom[34139] = 25'b0011110000100010010000101;
    rom[34140] = 25'b0011110000010110110000001;
    rom[34141] = 25'b0011110000001011001111011;
    rom[34142] = 25'b0011101111111111101110011;
    rom[34143] = 25'b0011101111110100001101001;
    rom[34144] = 25'b0011101111101000101011110;
    rom[34145] = 25'b0011101111011101001010000;
    rom[34146] = 25'b0011101111010001101000001;
    rom[34147] = 25'b0011101111000110000110000;
    rom[34148] = 25'b0011101110111010100011101;
    rom[34149] = 25'b0011101110101111000001001;
    rom[34150] = 25'b0011101110100011011110010;
    rom[34151] = 25'b0011101110010111111011010;
    rom[34152] = 25'b0011101110001100010111111;
    rom[34153] = 25'b0011101110000000110100100;
    rom[34154] = 25'b0011101101110101010000110;
    rom[34155] = 25'b0011101101101001101100111;
    rom[34156] = 25'b0011101101011110001000101;
    rom[34157] = 25'b0011101101010010100100010;
    rom[34158] = 25'b0011101101000110111111101;
    rom[34159] = 25'b0011101100111011011010110;
    rom[34160] = 25'b0011101100101111110101110;
    rom[34161] = 25'b0011101100100100010000100;
    rom[34162] = 25'b0011101100011000101011000;
    rom[34163] = 25'b0011101100001101000101011;
    rom[34164] = 25'b0011101100000001011111011;
    rom[34165] = 25'b0011101011110101111001010;
    rom[34166] = 25'b0011101011101010010010111;
    rom[34167] = 25'b0011101011011110101100011;
    rom[34168] = 25'b0011101011010011000101100;
    rom[34169] = 25'b0011101011000111011110100;
    rom[34170] = 25'b0011101010111011110111011;
    rom[34171] = 25'b0011101010110000001111111;
    rom[34172] = 25'b0011101010100100101000010;
    rom[34173] = 25'b0011101010011001000000011;
    rom[34174] = 25'b0011101010001101011000011;
    rom[34175] = 25'b0011101010000001110000000;
    rom[34176] = 25'b0011101001110110000111100;
    rom[34177] = 25'b0011101001101010011110111;
    rom[34178] = 25'b0011101001011110110101111;
    rom[34179] = 25'b0011101001010011001100110;
    rom[34180] = 25'b0011101001000111100011100;
    rom[34181] = 25'b0011101000111011111010000;
    rom[34182] = 25'b0011101000110000010000001;
    rom[34183] = 25'b0011101000100100100110010;
    rom[34184] = 25'b0011101000011000111100000;
    rom[34185] = 25'b0011101000001101010001110;
    rom[34186] = 25'b0011101000000001100111001;
    rom[34187] = 25'b0011100111110101111100011;
    rom[34188] = 25'b0011100111101010010001011;
    rom[34189] = 25'b0011100111011110100110001;
    rom[34190] = 25'b0011100111010010111010110;
    rom[34191] = 25'b0011100111000111001111010;
    rom[34192] = 25'b0011100110111011100011100;
    rom[34193] = 25'b0011100110101111110111011;
    rom[34194] = 25'b0011100110100100001011010;
    rom[34195] = 25'b0011100110011000011110110;
    rom[34196] = 25'b0011100110001100110010010;
    rom[34197] = 25'b0011100110000001000101100;
    rom[34198] = 25'b0011100101110101011000100;
    rom[34199] = 25'b0011100101101001101011010;
    rom[34200] = 25'b0011100101011101111101111;
    rom[34201] = 25'b0011100101010010010000010;
    rom[34202] = 25'b0011100101000110100010100;
    rom[34203] = 25'b0011100100111010110100101;
    rom[34204] = 25'b0011100100101111000110011;
    rom[34205] = 25'b0011100100100011011000000;
    rom[34206] = 25'b0011100100010111101001100;
    rom[34207] = 25'b0011100100001011111010101;
    rom[34208] = 25'b0011100100000000001011110;
    rom[34209] = 25'b0011100011110100011100101;
    rom[34210] = 25'b0011100011101000101101011;
    rom[34211] = 25'b0011100011011100111101110;
    rom[34212] = 25'b0011100011010001001110001;
    rom[34213] = 25'b0011100011000101011110001;
    rom[34214] = 25'b0011100010111001101110001;
    rom[34215] = 25'b0011100010101101111101111;
    rom[34216] = 25'b0011100010100010001101011;
    rom[34217] = 25'b0011100010010110011100110;
    rom[34218] = 25'b0011100010001010101011111;
    rom[34219] = 25'b0011100001111110111010111;
    rom[34220] = 25'b0011100001110011001001101;
    rom[34221] = 25'b0011100001100111011000010;
    rom[34222] = 25'b0011100001011011100110101;
    rom[34223] = 25'b0011100001001111110100111;
    rom[34224] = 25'b0011100001000100000011000;
    rom[34225] = 25'b0011100000111000010000110;
    rom[34226] = 25'b0011100000101100011110100;
    rom[34227] = 25'b0011100000100000101100000;
    rom[34228] = 25'b0011100000010100111001011;
    rom[34229] = 25'b0011100000001001000110100;
    rom[34230] = 25'b0011011111111101010011100;
    rom[34231] = 25'b0011011111110001100000010;
    rom[34232] = 25'b0011011111100101101100111;
    rom[34233] = 25'b0011011111011001111001010;
    rom[34234] = 25'b0011011111001110000101100;
    rom[34235] = 25'b0011011111000010010001101;
    rom[34236] = 25'b0011011110110110011101100;
    rom[34237] = 25'b0011011110101010101001010;
    rom[34238] = 25'b0011011110011110110100110;
    rom[34239] = 25'b0011011110010011000000001;
    rom[34240] = 25'b0011011110000111001011011;
    rom[34241] = 25'b0011011101111011010110011;
    rom[34242] = 25'b0011011101101111100001010;
    rom[34243] = 25'b0011011101100011101100000;
    rom[34244] = 25'b0011011101010111110110011;
    rom[34245] = 25'b0011011101001100000000110;
    rom[34246] = 25'b0011011101000000001010111;
    rom[34247] = 25'b0011011100110100010101000;
    rom[34248] = 25'b0011011100101000011110110;
    rom[34249] = 25'b0011011100011100101000100;
    rom[34250] = 25'b0011011100010000110010000;
    rom[34251] = 25'b0011011100000100111011011;
    rom[34252] = 25'b0011011011111001000100100;
    rom[34253] = 25'b0011011011101101001101011;
    rom[34254] = 25'b0011011011100001010110010;
    rom[34255] = 25'b0011011011010101011110111;
    rom[34256] = 25'b0011011011001001100111011;
    rom[34257] = 25'b0011011010111101101111110;
    rom[34258] = 25'b0011011010110001110111111;
    rom[34259] = 25'b0011011010100101111111111;
    rom[34260] = 25'b0011011010011010000111111;
    rom[34261] = 25'b0011011010001110001111100;
    rom[34262] = 25'b0011011010000010010111000;
    rom[34263] = 25'b0011011001110110011110011;
    rom[34264] = 25'b0011011001101010100101101;
    rom[34265] = 25'b0011011001011110101100101;
    rom[34266] = 25'b0011011001010010110011101;
    rom[34267] = 25'b0011011001000110111010010;
    rom[34268] = 25'b0011011000111011000000111;
    rom[34269] = 25'b0011011000101111000111010;
    rom[34270] = 25'b0011011000100011001101100;
    rom[34271] = 25'b0011011000010111010011101;
    rom[34272] = 25'b0011011000001011011001101;
    rom[34273] = 25'b0011010111111111011111011;
    rom[34274] = 25'b0011010111110011100101000;
    rom[34275] = 25'b0011010111100111101010100;
    rom[34276] = 25'b0011010111011011101111111;
    rom[34277] = 25'b0011010111001111110101000;
    rom[34278] = 25'b0011010111000011111010001;
    rom[34279] = 25'b0011010110110111111110111;
    rom[34280] = 25'b0011010110101100000011101;
    rom[34281] = 25'b0011010110100000001000010;
    rom[34282] = 25'b0011010110010100001100110;
    rom[34283] = 25'b0011010110001000010001000;
    rom[34284] = 25'b0011010101111100010101001;
    rom[34285] = 25'b0011010101110000011001001;
    rom[34286] = 25'b0011010101100100011100111;
    rom[34287] = 25'b0011010101011000100000101;
    rom[34288] = 25'b0011010101001100100100001;
    rom[34289] = 25'b0011010101000000100111101;
    rom[34290] = 25'b0011010100110100101010111;
    rom[34291] = 25'b0011010100101000101101111;
    rom[34292] = 25'b0011010100011100110000111;
    rom[34293] = 25'b0011010100010000110011110;
    rom[34294] = 25'b0011010100000100110110100;
    rom[34295] = 25'b0011010011111000111001000;
    rom[34296] = 25'b0011010011101100111011011;
    rom[34297] = 25'b0011010011100000111101101;
    rom[34298] = 25'b0011010011010100111111110;
    rom[34299] = 25'b0011010011001001000001110;
    rom[34300] = 25'b0011010010111101000011101;
    rom[34301] = 25'b0011010010110001000101010;
    rom[34302] = 25'b0011010010100101000110111;
    rom[34303] = 25'b0011010010011001001000011;
    rom[34304] = 25'b0011010010001101001001101;
    rom[34305] = 25'b0011010010000001001010110;
    rom[34306] = 25'b0011010001110101001011110;
    rom[34307] = 25'b0011010001101001001100101;
    rom[34308] = 25'b0011010001011101001101011;
    rom[34309] = 25'b0011010001010001001110000;
    rom[34310] = 25'b0011010001000101001110101;
    rom[34311] = 25'b0011010000111001001111000;
    rom[34312] = 25'b0011010000101101001111001;
    rom[34313] = 25'b0011010000100001001111010;
    rom[34314] = 25'b0011010000010101001111001;
    rom[34315] = 25'b0011010000001001001111001;
    rom[34316] = 25'b0011001111111101001110110;
    rom[34317] = 25'b0011001111110001001110010;
    rom[34318] = 25'b0011001111100101001101111;
    rom[34319] = 25'b0011001111011001001101001;
    rom[34320] = 25'b0011001111001101001100010;
    rom[34321] = 25'b0011001111000001001011011;
    rom[34322] = 25'b0011001110110101001010010;
    rom[34323] = 25'b0011001110101001001001001;
    rom[34324] = 25'b0011001110011101000111111;
    rom[34325] = 25'b0011001110010001000110011;
    rom[34326] = 25'b0011001110000101000100111;
    rom[34327] = 25'b0011001101111001000011010;
    rom[34328] = 25'b0011001101101101000001011;
    rom[34329] = 25'b0011001101100000111111100;
    rom[34330] = 25'b0011001101010100111101011;
    rom[34331] = 25'b0011001101001000111011010;
    rom[34332] = 25'b0011001100111100111001000;
    rom[34333] = 25'b0011001100110000110110101;
    rom[34334] = 25'b0011001100100100110100001;
    rom[34335] = 25'b0011001100011000110001100;
    rom[34336] = 25'b0011001100001100101110101;
    rom[34337] = 25'b0011001100000000101011111;
    rom[34338] = 25'b0011001011110100101000111;
    rom[34339] = 25'b0011001011101000100101110;
    rom[34340] = 25'b0011001011011100100010100;
    rom[34341] = 25'b0011001011010000011111001;
    rom[34342] = 25'b0011001011000100011011101;
    rom[34343] = 25'b0011001010111000011000010;
    rom[34344] = 25'b0011001010101100010100100;
    rom[34345] = 25'b0011001010100000010000110;
    rom[34346] = 25'b0011001010010100001100110;
    rom[34347] = 25'b0011001010001000001000111;
    rom[34348] = 25'b0011001001111100000100110;
    rom[34349] = 25'b0011001001110000000000100;
    rom[34350] = 25'b0011001001100011111100001;
    rom[34351] = 25'b0011001001010111110111110;
    rom[34352] = 25'b0011001001001011110011001;
    rom[34353] = 25'b0011001000111111101110100;
    rom[34354] = 25'b0011001000110011101001110;
    rom[34355] = 25'b0011001000100111100100111;
    rom[34356] = 25'b0011001000011011011111111;
    rom[34357] = 25'b0011001000001111011010110;
    rom[34358] = 25'b0011001000000011010101101;
    rom[34359] = 25'b0011000111110111010000011;
    rom[34360] = 25'b0011000111101011001010111;
    rom[34361] = 25'b0011000111011111000101011;
    rom[34362] = 25'b0011000111010010111111110;
    rom[34363] = 25'b0011000111000110111010001;
    rom[34364] = 25'b0011000110111010110100011;
    rom[34365] = 25'b0011000110101110101110011;
    rom[34366] = 25'b0011000110100010101000011;
    rom[34367] = 25'b0011000110010110100010010;
    rom[34368] = 25'b0011000110001010011100001;
    rom[34369] = 25'b0011000101111110010101111;
    rom[34370] = 25'b0011000101110010001111011;
    rom[34371] = 25'b0011000101100110001000111;
    rom[34372] = 25'b0011000101011010000010011;
    rom[34373] = 25'b0011000101001101111011101;
    rom[34374] = 25'b0011000101000001110100111;
    rom[34375] = 25'b0011000100110101101110000;
    rom[34376] = 25'b0011000100101001100111000;
    rom[34377] = 25'b0011000100011101011111111;
    rom[34378] = 25'b0011000100010001011000111;
    rom[34379] = 25'b0011000100000101010001100;
    rom[34380] = 25'b0011000011111001001010010;
    rom[34381] = 25'b0011000011101101000010111;
    rom[34382] = 25'b0011000011100000111011010;
    rom[34383] = 25'b0011000011010100110011101;
    rom[34384] = 25'b0011000011001000101100000;
    rom[34385] = 25'b0011000010111100100100010;
    rom[34386] = 25'b0011000010110000011100010;
    rom[34387] = 25'b0011000010100100010100011;
    rom[34388] = 25'b0011000010011000001100010;
    rom[34389] = 25'b0011000010001100000100001;
    rom[34390] = 25'b0011000001111111111011111;
    rom[34391] = 25'b0011000001110011110011101;
    rom[34392] = 25'b0011000001100111101011010;
    rom[34393] = 25'b0011000001011011100010110;
    rom[34394] = 25'b0011000001001111011010010;
    rom[34395] = 25'b0011000001000011010001100;
    rom[34396] = 25'b0011000000110111001000111;
    rom[34397] = 25'b0011000000101011000000000;
    rom[34398] = 25'b0011000000011110110111001;
    rom[34399] = 25'b0011000000010010101110001;
    rom[34400] = 25'b0011000000000110100101001;
    rom[34401] = 25'b0010111111111010011100000;
    rom[34402] = 25'b0010111111101110010010111;
    rom[34403] = 25'b0010111111100010001001100;
    rom[34404] = 25'b0010111111010110000000001;
    rom[34405] = 25'b0010111111001001110110110;
    rom[34406] = 25'b0010111110111101101101010;
    rom[34407] = 25'b0010111110110001100011101;
    rom[34408] = 25'b0010111110100101011010000;
    rom[34409] = 25'b0010111110011001010000010;
    rom[34410] = 25'b0010111110001101000110011;
    rom[34411] = 25'b0010111110000000111100100;
    rom[34412] = 25'b0010111101110100110010101;
    rom[34413] = 25'b0010111101101000101000101;
    rom[34414] = 25'b0010111101011100011110100;
    rom[34415] = 25'b0010111101010000010100010;
    rom[34416] = 25'b0010111101000100001010000;
    rom[34417] = 25'b0010111100110111111111110;
    rom[34418] = 25'b0010111100101011110101011;
    rom[34419] = 25'b0010111100011111101010111;
    rom[34420] = 25'b0010111100010011100000011;
    rom[34421] = 25'b0010111100000111010101111;
    rom[34422] = 25'b0010111011111011001011001;
    rom[34423] = 25'b0010111011101111000000011;
    rom[34424] = 25'b0010111011100010110101101;
    rom[34425] = 25'b0010111011010110101010111;
    rom[34426] = 25'b0010111011001010011111111;
    rom[34427] = 25'b0010111010111110010100111;
    rom[34428] = 25'b0010111010110010001001110;
    rom[34429] = 25'b0010111010100101111110110;
    rom[34430] = 25'b0010111010011001110011100;
    rom[34431] = 25'b0010111010001101101000011;
    rom[34432] = 25'b0010111010000001011101000;
    rom[34433] = 25'b0010111001110101010001110;
    rom[34434] = 25'b0010111001101001000110010;
    rom[34435] = 25'b0010111001011100111010110;
    rom[34436] = 25'b0010111001010000101111010;
    rom[34437] = 25'b0010111001000100100011110;
    rom[34438] = 25'b0010111000111000011000001;
    rom[34439] = 25'b0010111000101100001100011;
    rom[34440] = 25'b0010111000100000000000101;
    rom[34441] = 25'b0010111000010011110100110;
    rom[34442] = 25'b0010111000000111101001000;
    rom[34443] = 25'b0010110111111011011101000;
    rom[34444] = 25'b0010110111101111010001000;
    rom[34445] = 25'b0010110111100011000101000;
    rom[34446] = 25'b0010110111010110111000111;
    rom[34447] = 25'b0010110111001010101100110;
    rom[34448] = 25'b0010110110111110100000101;
    rom[34449] = 25'b0010110110110010010100011;
    rom[34450] = 25'b0010110110100110001000001;
    rom[34451] = 25'b0010110110011001111011110;
    rom[34452] = 25'b0010110110001101101111011;
    rom[34453] = 25'b0010110110000001100010111;
    rom[34454] = 25'b0010110101110101010110100;
    rom[34455] = 25'b0010110101101001001001111;
    rom[34456] = 25'b0010110101011100111101010;
    rom[34457] = 25'b0010110101010000110000101;
    rom[34458] = 25'b0010110101000100100100000;
    rom[34459] = 25'b0010110100111000010111010;
    rom[34460] = 25'b0010110100101100001010100;
    rom[34461] = 25'b0010110100011111111101110;
    rom[34462] = 25'b0010110100010011110000111;
    rom[34463] = 25'b0010110100000111100100000;
    rom[34464] = 25'b0010110011111011010111000;
    rom[34465] = 25'b0010110011101111001010001;
    rom[34466] = 25'b0010110011100010111101000;
    rom[34467] = 25'b0010110011010110110000000;
    rom[34468] = 25'b0010110011001010100011000;
    rom[34469] = 25'b0010110010111110010101110;
    rom[34470] = 25'b0010110010110010001000101;
    rom[34471] = 25'b0010110010100101111011011;
    rom[34472] = 25'b0010110010011001101110001;
    rom[34473] = 25'b0010110010001101100000111;
    rom[34474] = 25'b0010110010000001010011100;
    rom[34475] = 25'b0010110001110101000110010;
    rom[34476] = 25'b0010110001101000111000110;
    rom[34477] = 25'b0010110001011100101011011;
    rom[34478] = 25'b0010110001010000011101111;
    rom[34479] = 25'b0010110001000100010000011;
    rom[34480] = 25'b0010110000111000000010110;
    rom[34481] = 25'b0010110000101011110101010;
    rom[34482] = 25'b0010110000011111100111101;
    rom[34483] = 25'b0010110000010011011010000;
    rom[34484] = 25'b0010110000000111001100011;
    rom[34485] = 25'b0010101111111010111110110;
    rom[34486] = 25'b0010101111101110110001000;
    rom[34487] = 25'b0010101111100010100011010;
    rom[34488] = 25'b0010101111010110010101100;
    rom[34489] = 25'b0010101111001010000111101;
    rom[34490] = 25'b0010101110111101111001111;
    rom[34491] = 25'b0010101110110001101100000;
    rom[34492] = 25'b0010101110100101011110001;
    rom[34493] = 25'b0010101110011001010000001;
    rom[34494] = 25'b0010101110001101000010010;
    rom[34495] = 25'b0010101110000000110100010;
    rom[34496] = 25'b0010101101110100100110011;
    rom[34497] = 25'b0010101101101000011000011;
    rom[34498] = 25'b0010101101011100001010010;
    rom[34499] = 25'b0010101101001111111100010;
    rom[34500] = 25'b0010101101000011101110001;
    rom[34501] = 25'b0010101100110111100000000;
    rom[34502] = 25'b0010101100101011010001111;
    rom[34503] = 25'b0010101100011111000011111;
    rom[34504] = 25'b0010101100010010110101110;
    rom[34505] = 25'b0010101100000110100111100;
    rom[34506] = 25'b0010101011111010011001011;
    rom[34507] = 25'b0010101011101110001011001;
    rom[34508] = 25'b0010101011100001111101000;
    rom[34509] = 25'b0010101011010101101110101;
    rom[34510] = 25'b0010101011001001100000100;
    rom[34511] = 25'b0010101010111101010010001;
    rom[34512] = 25'b0010101010110001000011111;
    rom[34513] = 25'b0010101010100100110101101;
    rom[34514] = 25'b0010101010011000100111010;
    rom[34515] = 25'b0010101010001100011000111;
    rom[34516] = 25'b0010101010000000001010101;
    rom[34517] = 25'b0010101001110011111100011;
    rom[34518] = 25'b0010101001100111101101111;
    rom[34519] = 25'b0010101001011011011111100;
    rom[34520] = 25'b0010101001001111010001010;
    rom[34521] = 25'b0010101001000011000010111;
    rom[34522] = 25'b0010101000110110110100011;
    rom[34523] = 25'b0010101000101010100110000;
    rom[34524] = 25'b0010101000011110010111101;
    rom[34525] = 25'b0010101000010010001001001;
    rom[34526] = 25'b0010101000000101111010110;
    rom[34527] = 25'b0010100111111001101100011;
    rom[34528] = 25'b0010100111101101011101111;
    rom[34529] = 25'b0010100111100001001111100;
    rom[34530] = 25'b0010100111010101000001001;
    rom[34531] = 25'b0010100111001000110010101;
    rom[34532] = 25'b0010100110111100100100001;
    rom[34533] = 25'b0010100110110000010101110;
    rom[34534] = 25'b0010100110100100000111010;
    rom[34535] = 25'b0010100110010111111000110;
    rom[34536] = 25'b0010100110001011101010011;
    rom[34537] = 25'b0010100101111111011011111;
    rom[34538] = 25'b0010100101110011001101011;
    rom[34539] = 25'b0010100101100110111111000;
    rom[34540] = 25'b0010100101011010110000100;
    rom[34541] = 25'b0010100101001110100010000;
    rom[34542] = 25'b0010100101000010010011101;
    rom[34543] = 25'b0010100100110110000101001;
    rom[34544] = 25'b0010100100101001110110110;
    rom[34545] = 25'b0010100100011101101000011;
    rom[34546] = 25'b0010100100010001011001111;
    rom[34547] = 25'b0010100100000101001011100;
    rom[34548] = 25'b0010100011111000111101001;
    rom[34549] = 25'b0010100011101100101110110;
    rom[34550] = 25'b0010100011100000100000010;
    rom[34551] = 25'b0010100011010100010001111;
    rom[34552] = 25'b0010100011001000000011100;
    rom[34553] = 25'b0010100010111011110101001;
    rom[34554] = 25'b0010100010101111100110110;
    rom[34555] = 25'b0010100010100011011000011;
    rom[34556] = 25'b0010100010010111001010001;
    rom[34557] = 25'b0010100010001010111011110;
    rom[34558] = 25'b0010100001111110101101011;
    rom[34559] = 25'b0010100001110010011111001;
    rom[34560] = 25'b0010100001100110010000110;
    rom[34561] = 25'b0010100001011010000010101;
    rom[34562] = 25'b0010100001001101110100010;
    rom[34563] = 25'b0010100001000001100110001;
    rom[34564] = 25'b0010100000110101010111110;
    rom[34565] = 25'b0010100000101001001001101;
    rom[34566] = 25'b0010100000011100111011011;
    rom[34567] = 25'b0010100000010000101101010;
    rom[34568] = 25'b0010100000000100011111000;
    rom[34569] = 25'b0010011111111000010000111;
    rom[34570] = 25'b0010011111101100000010110;
    rom[34571] = 25'b0010011111011111110100110;
    rom[34572] = 25'b0010011111010011100110101;
    rom[34573] = 25'b0010011111000111011000100;
    rom[34574] = 25'b0010011110111011001010011;
    rom[34575] = 25'b0010011110101110111100011;
    rom[34576] = 25'b0010011110100010101110100;
    rom[34577] = 25'b0010011110010110100000100;
    rom[34578] = 25'b0010011110001010010010100;
    rom[34579] = 25'b0010011101111110000100101;
    rom[34580] = 25'b0010011101110001110110101;
    rom[34581] = 25'b0010011101100101101000111;
    rom[34582] = 25'b0010011101011001011010111;
    rom[34583] = 25'b0010011101001101001101001;
    rom[34584] = 25'b0010011101000000111111011;
    rom[34585] = 25'b0010011100110100110001101;
    rom[34586] = 25'b0010011100101000100011111;
    rom[34587] = 25'b0010011100011100010110001;
    rom[34588] = 25'b0010011100010000001000100;
    rom[34589] = 25'b0010011100000011111010110;
    rom[34590] = 25'b0010011011110111101101001;
    rom[34591] = 25'b0010011011101011011111100;
    rom[34592] = 25'b0010011011011111010010000;
    rom[34593] = 25'b0010011011010011000100100;
    rom[34594] = 25'b0010011011000110110110111;
    rom[34595] = 25'b0010011010111010101001100;
    rom[34596] = 25'b0010011010101110011100000;
    rom[34597] = 25'b0010011010100010001110101;
    rom[34598] = 25'b0010011010010110000001010;
    rom[34599] = 25'b0010011010001001110100000;
    rom[34600] = 25'b0010011001111101100110110;
    rom[34601] = 25'b0010011001110001011001011;
    rom[34602] = 25'b0010011001100101001100001;
    rom[34603] = 25'b0010011001011000111111001;
    rom[34604] = 25'b0010011001001100110001111;
    rom[34605] = 25'b0010011001000000100100110;
    rom[34606] = 25'b0010011000110100010111110;
    rom[34607] = 25'b0010011000101000001010110;
    rom[34608] = 25'b0010011000011011111101110;
    rom[34609] = 25'b0010011000001111110000111;
    rom[34610] = 25'b0010011000000011100011111;
    rom[34611] = 25'b0010010111110111010111000;
    rom[34612] = 25'b0010010111101011001010010;
    rom[34613] = 25'b0010010111011110111101100;
    rom[34614] = 25'b0010010111010010110000110;
    rom[34615] = 25'b0010010111000110100100000;
    rom[34616] = 25'b0010010110111010010111011;
    rom[34617] = 25'b0010010110101110001010110;
    rom[34618] = 25'b0010010110100001111110010;
    rom[34619] = 25'b0010010110010101110001111;
    rom[34620] = 25'b0010010110001001100101011;
    rom[34621] = 25'b0010010101111101011001000;
    rom[34622] = 25'b0010010101110001001100101;
    rom[34623] = 25'b0010010101100101000000010;
    rom[34624] = 25'b0010010101011000110100000;
    rom[34625] = 25'b0010010101001100100111111;
    rom[34626] = 25'b0010010101000000011011110;
    rom[34627] = 25'b0010010100110100001111101;
    rom[34628] = 25'b0010010100101000000011101;
    rom[34629] = 25'b0010010100011011110111100;
    rom[34630] = 25'b0010010100001111101011101;
    rom[34631] = 25'b0010010100000011011111110;
    rom[34632] = 25'b0010010011110111010011111;
    rom[34633] = 25'b0010010011101011001000001;
    rom[34634] = 25'b0010010011011110111100100;
    rom[34635] = 25'b0010010011010010110000110;
    rom[34636] = 25'b0010010011000110100101001;
    rom[34637] = 25'b0010010010111010011001101;
    rom[34638] = 25'b0010010010101110001110001;
    rom[34639] = 25'b0010010010100010000010101;
    rom[34640] = 25'b0010010010010101110111010;
    rom[34641] = 25'b0010010010001001101100000;
    rom[34642] = 25'b0010010001111101100000110;
    rom[34643] = 25'b0010010001110001010101100;
    rom[34644] = 25'b0010010001100101001010011;
    rom[34645] = 25'b0010010001011000111111011;
    rom[34646] = 25'b0010010001001100110100010;
    rom[34647] = 25'b0010010001000000101001011;
    rom[34648] = 25'b0010010000110100011110011;
    rom[34649] = 25'b0010010000101000010011101;
    rom[34650] = 25'b0010010000011100001000111;
    rom[34651] = 25'b0010010000001111111110001;
    rom[34652] = 25'b0010010000000011110011101;
    rom[34653] = 25'b0010001111110111101001000;
    rom[34654] = 25'b0010001111101011011110100;
    rom[34655] = 25'b0010001111011111010100001;
    rom[34656] = 25'b0010001111010011001001110;
    rom[34657] = 25'b0010001111000110111111011;
    rom[34658] = 25'b0010001110111010110101010;
    rom[34659] = 25'b0010001110101110101011000;
    rom[34660] = 25'b0010001110100010100000111;
    rom[34661] = 25'b0010001110010110010110111;
    rom[34662] = 25'b0010001110001010001101000;
    rom[34663] = 25'b0010001101111110000011001;
    rom[34664] = 25'b0010001101110001111001011;
    rom[34665] = 25'b0010001101100101101111101;
    rom[34666] = 25'b0010001101011001100110000;
    rom[34667] = 25'b0010001101001101011100011;
    rom[34668] = 25'b0010001101000001010010111;
    rom[34669] = 25'b0010001100110101001001100;
    rom[34670] = 25'b0010001100101001000000001;
    rom[34671] = 25'b0010001100011100110110111;
    rom[34672] = 25'b0010001100010000101101101;
    rom[34673] = 25'b0010001100000100100100100;
    rom[34674] = 25'b0010001011111000011011100;
    rom[34675] = 25'b0010001011101100010010100;
    rom[34676] = 25'b0010001011100000001001101;
    rom[34677] = 25'b0010001011010100000000110;
    rom[34678] = 25'b0010001011000111111000001;
    rom[34679] = 25'b0010001010111011101111011;
    rom[34680] = 25'b0010001010101111100110111;
    rom[34681] = 25'b0010001010100011011110011;
    rom[34682] = 25'b0010001010010111010110000;
    rom[34683] = 25'b0010001010001011001101101;
    rom[34684] = 25'b0010001001111111000101011;
    rom[34685] = 25'b0010001001110010111101010;
    rom[34686] = 25'b0010001001100110110101010;
    rom[34687] = 25'b0010001001011010101101010;
    rom[34688] = 25'b0010001001001110100101010;
    rom[34689] = 25'b0010001001000010011101100;
    rom[34690] = 25'b0010001000110110010101110;
    rom[34691] = 25'b0010001000101010001110001;
    rom[34692] = 25'b0010001000011110000110101;
    rom[34693] = 25'b0010001000010001111111001;
    rom[34694] = 25'b0010001000000101110111111;
    rom[34695] = 25'b0010000111111001110000100;
    rom[34696] = 25'b0010000111101101101001010;
    rom[34697] = 25'b0010000111100001100010010;
    rom[34698] = 25'b0010000111010101011011001;
    rom[34699] = 25'b0010000111001001010100010;
    rom[34700] = 25'b0010000110111101001101100;
    rom[34701] = 25'b0010000110110001000110110;
    rom[34702] = 25'b0010000110100101000000001;
    rom[34703] = 25'b0010000110011000111001101;
    rom[34704] = 25'b0010000110001100110011001;
    rom[34705] = 25'b0010000110000000101100110;
    rom[34706] = 25'b0010000101110100100110100;
    rom[34707] = 25'b0010000101101000100000010;
    rom[34708] = 25'b0010000101011100011010010;
    rom[34709] = 25'b0010000101010000010100011;
    rom[34710] = 25'b0010000101000100001110011;
    rom[34711] = 25'b0010000100111000001000101;
    rom[34712] = 25'b0010000100101100000011000;
    rom[34713] = 25'b0010000100011111111101011;
    rom[34714] = 25'b0010000100010011111000000;
    rom[34715] = 25'b0010000100000111110010100;
    rom[34716] = 25'b0010000011111011101101010;
    rom[34717] = 25'b0010000011101111101000001;
    rom[34718] = 25'b0010000011100011100011001;
    rom[34719] = 25'b0010000011010111011110001;
    rom[34720] = 25'b0010000011001011011001010;
    rom[34721] = 25'b0010000010111111010100100;
    rom[34722] = 25'b0010000010110011001111110;
    rom[34723] = 25'b0010000010100111001011010;
    rom[34724] = 25'b0010000010011011000110110;
    rom[34725] = 25'b0010000010001111000010100;
    rom[34726] = 25'b0010000010000010111110010;
    rom[34727] = 25'b0010000001110110111010001;
    rom[34728] = 25'b0010000001101010110110001;
    rom[34729] = 25'b0010000001011110110010001;
    rom[34730] = 25'b0010000001010010101110011;
    rom[34731] = 25'b0010000001000110101010101;
    rom[34732] = 25'b0010000000111010100111001;
    rom[34733] = 25'b0010000000101110100011101;
    rom[34734] = 25'b0010000000100010100000010;
    rom[34735] = 25'b0010000000010110011101000;
    rom[34736] = 25'b0010000000001010011001111;
    rom[34737] = 25'b0001111111111110010110111;
    rom[34738] = 25'b0001111111110010010100000;
    rom[34739] = 25'b0001111111100110010001001;
    rom[34740] = 25'b0001111111011010001110011;
    rom[34741] = 25'b0001111111001110001011111;
    rom[34742] = 25'b0001111111000010001001011;
    rom[34743] = 25'b0001111110110110000111001;
    rom[34744] = 25'b0001111110101010000100111;
    rom[34745] = 25'b0001111110011110000010110;
    rom[34746] = 25'b0001111110010010000000110;
    rom[34747] = 25'b0001111110000101111110111;
    rom[34748] = 25'b0001111101111001111101001;
    rom[34749] = 25'b0001111101101101111011100;
    rom[34750] = 25'b0001111101100001111010000;
    rom[34751] = 25'b0001111101010101111000101;
    rom[34752] = 25'b0001111101001001110111011;
    rom[34753] = 25'b0001111100111101110110010;
    rom[34754] = 25'b0001111100110001110101001;
    rom[34755] = 25'b0001111100100101110100010;
    rom[34756] = 25'b0001111100011001110011100;
    rom[34757] = 25'b0001111100001101110010110;
    rom[34758] = 25'b0001111100000001110010011;
    rom[34759] = 25'b0001111011110101110001111;
    rom[34760] = 25'b0001111011101001110001100;
    rom[34761] = 25'b0001111011011101110001011;
    rom[34762] = 25'b0001111011010001110001011;
    rom[34763] = 25'b0001111011000101110001100;
    rom[34764] = 25'b0001111010111001110001101;
    rom[34765] = 25'b0001111010101101110010000;
    rom[34766] = 25'b0001111010100001110010100;
    rom[34767] = 25'b0001111010010101110011001;
    rom[34768] = 25'b0001111010001001110011111;
    rom[34769] = 25'b0001111001111101110100101;
    rom[34770] = 25'b0001111001110001110101101;
    rom[34771] = 25'b0001111001100101110110110;
    rom[34772] = 25'b0001111001011001111000001;
    rom[34773] = 25'b0001111001001101111001100;
    rom[34774] = 25'b0001111001000001111011000;
    rom[34775] = 25'b0001111000110101111100101;
    rom[34776] = 25'b0001111000101001111110100;
    rom[34777] = 25'b0001111000011110000000011;
    rom[34778] = 25'b0001111000010010000010011;
    rom[34779] = 25'b0001111000000110000100101;
    rom[34780] = 25'b0001110111111010000110111;
    rom[34781] = 25'b0001110111101110001001011;
    rom[34782] = 25'b0001110111100010001100000;
    rom[34783] = 25'b0001110111010110001110110;
    rom[34784] = 25'b0001110111001010010001101;
    rom[34785] = 25'b0001110110111110010100100;
    rom[34786] = 25'b0001110110110010010111110;
    rom[34787] = 25'b0001110110100110011011001;
    rom[34788] = 25'b0001110110011010011110100;
    rom[34789] = 25'b0001110110001110100010000;
    rom[34790] = 25'b0001110110000010100101110;
    rom[34791] = 25'b0001110101110110101001101;
    rom[34792] = 25'b0001110101101010101101101;
    rom[34793] = 25'b0001110101011110110001110;
    rom[34794] = 25'b0001110101010010110110000;
    rom[34795] = 25'b0001110101000110111010011;
    rom[34796] = 25'b0001110100111010111111001;
    rom[34797] = 25'b0001110100101111000011110;
    rom[34798] = 25'b0001110100100011001000101;
    rom[34799] = 25'b0001110100010111001101101;
    rom[34800] = 25'b0001110100001011010010110;
    rom[34801] = 25'b0001110011111111011000000;
    rom[34802] = 25'b0001110011110011011101100;
    rom[34803] = 25'b0001110011100111100011001;
    rom[34804] = 25'b0001110011011011101000111;
    rom[34805] = 25'b0001110011001111101110110;
    rom[34806] = 25'b0001110011000011110100110;
    rom[34807] = 25'b0001110010110111111011000;
    rom[34808] = 25'b0001110010101100000001010;
    rom[34809] = 25'b0001110010100000000111111;
    rom[34810] = 25'b0001110010010100001110011;
    rom[34811] = 25'b0001110010001000010101010;
    rom[34812] = 25'b0001110001111100011100010;
    rom[34813] = 25'b0001110001110000100011010;
    rom[34814] = 25'b0001110001100100101010101;
    rom[34815] = 25'b0001110001011000110010000;
    rom[34816] = 25'b0001110001001100111001101;
    rom[34817] = 25'b0001110001000001000001010;
    rom[34818] = 25'b0001110000110101001001001;
    rom[34819] = 25'b0001110000101001010001001;
    rom[34820] = 25'b0001110000011101011001011;
    rom[34821] = 25'b0001110000010001100001110;
    rom[34822] = 25'b0001110000000101101010010;
    rom[34823] = 25'b0001101111111001110010111;
    rom[34824] = 25'b0001101111101101111011101;
    rom[34825] = 25'b0001101111100010000100110;
    rom[34826] = 25'b0001101111010110001101111;
    rom[34827] = 25'b0001101111001010010111001;
    rom[34828] = 25'b0001101110111110100000101;
    rom[34829] = 25'b0001101110110010101010010;
    rom[34830] = 25'b0001101110100110110100000;
    rom[34831] = 25'b0001101110011010111110000;
    rom[34832] = 25'b0001101110001111001000000;
    rom[34833] = 25'b0001101110000011010010011;
    rom[34834] = 25'b0001101101110111011100111;
    rom[34835] = 25'b0001101101101011100111011;
    rom[34836] = 25'b0001101101011111110010010;
    rom[34837] = 25'b0001101101010011111101001;
    rom[34838] = 25'b0001101101001000001000010;
    rom[34839] = 25'b0001101100111100010011100;
    rom[34840] = 25'b0001101100110000011111000;
    rom[34841] = 25'b0001101100100100101010100;
    rom[34842] = 25'b0001101100011000110110010;
    rom[34843] = 25'b0001101100001101000010010;
    rom[34844] = 25'b0001101100000001001110011;
    rom[34845] = 25'b0001101011110101011010101;
    rom[34846] = 25'b0001101011101001100111000;
    rom[34847] = 25'b0001101011011101110011110;
    rom[34848] = 25'b0001101011010010000000100;
    rom[34849] = 25'b0001101011000110001101100;
    rom[34850] = 25'b0001101010111010011010101;
    rom[34851] = 25'b0001101010101110101000000;
    rom[34852] = 25'b0001101010100010110101011;
    rom[34853] = 25'b0001101010010111000011001;
    rom[34854] = 25'b0001101010001011010000111;
    rom[34855] = 25'b0001101001111111011110111;
    rom[34856] = 25'b0001101001110011101101001;
    rom[34857] = 25'b0001101001100111111011100;
    rom[34858] = 25'b0001101001011100001010000;
    rom[34859] = 25'b0001101001010000011000110;
    rom[34860] = 25'b0001101001000100100111101;
    rom[34861] = 25'b0001101000111000110110110;
    rom[34862] = 25'b0001101000101101000101111;
    rom[34863] = 25'b0001101000100001010101011;
    rom[34864] = 25'b0001101000010101100101000;
    rom[34865] = 25'b0001101000001001110100110;
    rom[34866] = 25'b0001100111111110000100110;
    rom[34867] = 25'b0001100111110010010101000;
    rom[34868] = 25'b0001100111100110100101010;
    rom[34869] = 25'b0001100111011010110101110;
    rom[34870] = 25'b0001100111001111000110100;
    rom[34871] = 25'b0001100111000011010111011;
    rom[34872] = 25'b0001100110110111101000100;
    rom[34873] = 25'b0001100110101011111001101;
    rom[34874] = 25'b0001100110100000001011001;
    rom[34875] = 25'b0001100110010100011100110;
    rom[34876] = 25'b0001100110001000101110100;
    rom[34877] = 25'b0001100101111101000000100;
    rom[34878] = 25'b0001100101110001010010110;
    rom[34879] = 25'b0001100101100101100101000;
    rom[34880] = 25'b0001100101011001110111101;
    rom[34881] = 25'b0001100101001110001010011;
    rom[34882] = 25'b0001100101000010011101010;
    rom[34883] = 25'b0001100100110110110000011;
    rom[34884] = 25'b0001100100101011000011110;
    rom[34885] = 25'b0001100100011111010111010;
    rom[34886] = 25'b0001100100010011101010111;
    rom[34887] = 25'b0001100100000111111110110;
    rom[34888] = 25'b0001100011111100010010111;
    rom[34889] = 25'b0001100011110000100111001;
    rom[34890] = 25'b0001100011100100111011101;
    rom[34891] = 25'b0001100011011001010000010;
    rom[34892] = 25'b0001100011001101100101001;
    rom[34893] = 25'b0001100011000001111010001;
    rom[34894] = 25'b0001100010110110001111011;
    rom[34895] = 25'b0001100010101010100100111;
    rom[34896] = 25'b0001100010011110111010100;
    rom[34897] = 25'b0001100010010011010000010;
    rom[34898] = 25'b0001100010000111100110011;
    rom[34899] = 25'b0001100001111011111100100;
    rom[34900] = 25'b0001100001110000010011000;
    rom[34901] = 25'b0001100001100100101001100;
    rom[34902] = 25'b0001100001011001000000011;
    rom[34903] = 25'b0001100001001101010111011;
    rom[34904] = 25'b0001100001000001101110101;
    rom[34905] = 25'b0001100000110110000110000;
    rom[34906] = 25'b0001100000101010011101101;
    rom[34907] = 25'b0001100000011110110101011;
    rom[34908] = 25'b0001100000010011001101100;
    rom[34909] = 25'b0001100000000111100101101;
    rom[34910] = 25'b0001011111111011111110001;
    rom[34911] = 25'b0001011111110000010110110;
    rom[34912] = 25'b0001011111100100101111101;
    rom[34913] = 25'b0001011111011001001000101;
    rom[34914] = 25'b0001011111001101100001111;
    rom[34915] = 25'b0001011111000001111011010;
    rom[34916] = 25'b0001011110110110010101000;
    rom[34917] = 25'b0001011110101010101110110;
    rom[34918] = 25'b0001011110011111001001000;
    rom[34919] = 25'b0001011110010011100011001;
    rom[34920] = 25'b0001011110000111111101101;
    rom[34921] = 25'b0001011101111100011000011;
    rom[34922] = 25'b0001011101110000110011010;
    rom[34923] = 25'b0001011101100101001110011;
    rom[34924] = 25'b0001011101011001101001101;
    rom[34925] = 25'b0001011101001110000101010;
    rom[34926] = 25'b0001011101000010100001000;
    rom[34927] = 25'b0001011100110110111100111;
    rom[34928] = 25'b0001011100101011011001001;
    rom[34929] = 25'b0001011100011111110101100;
    rom[34930] = 25'b0001011100010100010010000;
    rom[34931] = 25'b0001011100001000101110111;
    rom[34932] = 25'b0001011011111101001011111;
    rom[34933] = 25'b0001011011110001101001001;
    rom[34934] = 25'b0001011011100110000110100;
    rom[34935] = 25'b0001011011011010100100010;
    rom[34936] = 25'b0001011011001111000010001;
    rom[34937] = 25'b0001011011000011100000010;
    rom[34938] = 25'b0001011010110111111110100;
    rom[34939] = 25'b0001011010101100011101000;
    rom[34940] = 25'b0001011010100000111011110;
    rom[34941] = 25'b0001011010010101011010110;
    rom[34942] = 25'b0001011010001001111010000;
    rom[34943] = 25'b0001011001111110011001011;
    rom[34944] = 25'b0001011001110010111001000;
    rom[34945] = 25'b0001011001100111011000110;
    rom[34946] = 25'b0001011001011011111000111;
    rom[34947] = 25'b0001011001010000011001010;
    rom[34948] = 25'b0001011001000100111001110;
    rom[34949] = 25'b0001011000111001011010011;
    rom[34950] = 25'b0001011000101101111011011;
    rom[34951] = 25'b0001011000100010011100100;
    rom[34952] = 25'b0001011000010110111110000;
    rom[34953] = 25'b0001011000001011011111101;
    rom[34954] = 25'b0001011000000000000001011;
    rom[34955] = 25'b0001010111110100100011011;
    rom[34956] = 25'b0001010111101001000101110;
    rom[34957] = 25'b0001010111011101101000011;
    rom[34958] = 25'b0001010111010010001011000;
    rom[34959] = 25'b0001010111000110101110000;
    rom[34960] = 25'b0001010110111011010001010;
    rom[34961] = 25'b0001010110101111110100110;
    rom[34962] = 25'b0001010110100100011000011;
    rom[34963] = 25'b0001010110011000111100010;
    rom[34964] = 25'b0001010110001101100000011;
    rom[34965] = 25'b0001010110000010000100110;
    rom[34966] = 25'b0001010101110110101001010;
    rom[34967] = 25'b0001010101101011001110001;
    rom[34968] = 25'b0001010101011111110011010;
    rom[34969] = 25'b0001010101010100011000011;
    rom[34970] = 25'b0001010101001000111110000;
    rom[34971] = 25'b0001010100111101100011101;
    rom[34972] = 25'b0001010100110010001001101;
    rom[34973] = 25'b0001010100100110101111111;
    rom[34974] = 25'b0001010100011011010110010;
    rom[34975] = 25'b0001010100001111111101000;
    rom[34976] = 25'b0001010100000100100011111;
    rom[34977] = 25'b0001010011111001001011001;
    rom[34978] = 25'b0001010011101101110010011;
    rom[34979] = 25'b0001010011100010011010001;
    rom[34980] = 25'b0001010011010111000001111;
    rom[34981] = 25'b0001010011001011101010000;
    rom[34982] = 25'b0001010011000000010010011;
    rom[34983] = 25'b0001010010110100111010111;
    rom[34984] = 25'b0001010010101001100011110;
    rom[34985] = 25'b0001010010011110001100110;
    rom[34986] = 25'b0001010010010010110110000;
    rom[34987] = 25'b0001010010000111011111101;
    rom[34988] = 25'b0001010001111100001001011;
    rom[34989] = 25'b0001010001110000110011011;
    rom[34990] = 25'b0001010001100101011101110;
    rom[34991] = 25'b0001010001011010001000001;
    rom[34992] = 25'b0001010001001110110011000;
    rom[34993] = 25'b0001010001000011011101111;
    rom[34994] = 25'b0001010000111000001001001;
    rom[34995] = 25'b0001010000101100110100101;
    rom[34996] = 25'b0001010000100001100000010;
    rom[34997] = 25'b0001010000010110001100010;
    rom[34998] = 25'b0001010000001010111000100;
    rom[34999] = 25'b0001001111111111100101000;
    rom[35000] = 25'b0001001111110100010001101;
    rom[35001] = 25'b0001001111101000111110101;
    rom[35002] = 25'b0001001111011101101011111;
    rom[35003] = 25'b0001001111010010011001010;
    rom[35004] = 25'b0001001111000111000111000;
    rom[35005] = 25'b0001001110111011110100111;
    rom[35006] = 25'b0001001110110000100011001;
    rom[35007] = 25'b0001001110100101010001100;
    rom[35008] = 25'b0001001110011010000000010;
    rom[35009] = 25'b0001001110001110101111001;
    rom[35010] = 25'b0001001110000011011110011;
    rom[35011] = 25'b0001001101111000001101111;
    rom[35012] = 25'b0001001101101100111101100;
    rom[35013] = 25'b0001001101100001101101100;
    rom[35014] = 25'b0001001101010110011101101;
    rom[35015] = 25'b0001001101001011001110001;
    rom[35016] = 25'b0001001100111111111110111;
    rom[35017] = 25'b0001001100110100101111111;
    rom[35018] = 25'b0001001100101001100001001;
    rom[35019] = 25'b0001001100011110010010101;
    rom[35020] = 25'b0001001100010011000100011;
    rom[35021] = 25'b0001001100000111110110010;
    rom[35022] = 25'b0001001011111100101000100;
    rom[35023] = 25'b0001001011110001011011000;
    rom[35024] = 25'b0001001011100110001101110;
    rom[35025] = 25'b0001001011011011000000111;
    rom[35026] = 25'b0001001011001111110100001;
    rom[35027] = 25'b0001001011000100100111101;
    rom[35028] = 25'b0001001010111001011011100;
    rom[35029] = 25'b0001001010101110001111100;
    rom[35030] = 25'b0001001010100011000011111;
    rom[35031] = 25'b0001001010010111111000011;
    rom[35032] = 25'b0001001010001100101101010;
    rom[35033] = 25'b0001001010000001100010011;
    rom[35034] = 25'b0001001001110110010111110;
    rom[35035] = 25'b0001001001101011001101011;
    rom[35036] = 25'b0001001001100000000011010;
    rom[35037] = 25'b0001001001010100111001011;
    rom[35038] = 25'b0001001001001001101111111;
    rom[35039] = 25'b0001001000111110100110100;
    rom[35040] = 25'b0001001000110011011101100;
    rom[35041] = 25'b0001001000101000010100110;
    rom[35042] = 25'b0001001000011101001100010;
    rom[35043] = 25'b0001001000010010000100000;
    rom[35044] = 25'b0001001000000110111100000;
    rom[35045] = 25'b0001000111111011110100010;
    rom[35046] = 25'b0001000111110000101100110;
    rom[35047] = 25'b0001000111100101100101101;
    rom[35048] = 25'b0001000111011010011110110;
    rom[35049] = 25'b0001000111001111011000001;
    rom[35050] = 25'b0001000111000100010001110;
    rom[35051] = 25'b0001000110111001001011101;
    rom[35052] = 25'b0001000110101110000101111;
    rom[35053] = 25'b0001000110100011000000010;
    rom[35054] = 25'b0001000110010111111010111;
    rom[35055] = 25'b0001000110001100110101111;
    rom[35056] = 25'b0001000110000001110001010;
    rom[35057] = 25'b0001000101110110101100110;
    rom[35058] = 25'b0001000101101011101000100;
    rom[35059] = 25'b0001000101100000100100101;
    rom[35060] = 25'b0001000101010101100001000;
    rom[35061] = 25'b0001000101001010011101101;
    rom[35062] = 25'b0001000100111111011010100;
    rom[35063] = 25'b0001000100110100010111110;
    rom[35064] = 25'b0001000100101001010101001;
    rom[35065] = 25'b0001000100011110010010111;
    rom[35066] = 25'b0001000100010011010000111;
    rom[35067] = 25'b0001000100001000001111010;
    rom[35068] = 25'b0001000011111101001101110;
    rom[35069] = 25'b0001000011110010001100101;
    rom[35070] = 25'b0001000011100111001011110;
    rom[35071] = 25'b0001000011011100001011001;
    rom[35072] = 25'b0001000011010001001010110;
    rom[35073] = 25'b0001000011000110001010111;
    rom[35074] = 25'b0001000010111011001011000;
    rom[35075] = 25'b0001000010110000001011101;
    rom[35076] = 25'b0001000010100101001100011;
    rom[35077] = 25'b0001000010011010001101100;
    rom[35078] = 25'b0001000010001111001110110;
    rom[35079] = 25'b0001000010000100010000011;
    rom[35080] = 25'b0001000001111001010010011;
    rom[35081] = 25'b0001000001101110010100101;
    rom[35082] = 25'b0001000001100011010111001;
    rom[35083] = 25'b0001000001011000011001111;
    rom[35084] = 25'b0001000001001101011101000;
    rom[35085] = 25'b0001000001000010100000011;
    rom[35086] = 25'b0001000000110111100100000;
    rom[35087] = 25'b0001000000101100100111111;
    rom[35088] = 25'b0001000000100001101100001;
    rom[35089] = 25'b0001000000010110110000101;
    rom[35090] = 25'b0001000000001011110101011;
    rom[35091] = 25'b0001000000000000111010100;
    rom[35092] = 25'b0000111111110101111111111;
    rom[35093] = 25'b0000111111101011000101100;
    rom[35094] = 25'b0000111111100000001011100;
    rom[35095] = 25'b0000111111010101010001110;
    rom[35096] = 25'b0000111111001010011000010;
    rom[35097] = 25'b0000111110111111011111001;
    rom[35098] = 25'b0000111110110100100110001;
    rom[35099] = 25'b0000111110101001101101101;
    rom[35100] = 25'b0000111110011110110101010;
    rom[35101] = 25'b0000111110010011111101010;
    rom[35102] = 25'b0000111110001001000101100;
    rom[35103] = 25'b0000111101111110001110001;
    rom[35104] = 25'b0000111101110011010111000;
    rom[35105] = 25'b0000111101101000100000001;
    rom[35106] = 25'b0000111101011101101001101;
    rom[35107] = 25'b0000111101010010110011011;
    rom[35108] = 25'b0000111101000111111101011;
    rom[35109] = 25'b0000111100111101000111110;
    rom[35110] = 25'b0000111100110010010010011;
    rom[35111] = 25'b0000111100100111011101010;
    rom[35112] = 25'b0000111100011100101000100;
    rom[35113] = 25'b0000111100010001110100001;
    rom[35114] = 25'b0000111100000110111111111;
    rom[35115] = 25'b0000111011111100001100000;
    rom[35116] = 25'b0000111011110001011000100;
    rom[35117] = 25'b0000111011100110100101010;
    rom[35118] = 25'b0000111011011011110010001;
    rom[35119] = 25'b0000111011010000111111100;
    rom[35120] = 25'b0000111011000110001101001;
    rom[35121] = 25'b0000111010111011011011001;
    rom[35122] = 25'b0000111010110000101001010;
    rom[35123] = 25'b0000111010100101110111111;
    rom[35124] = 25'b0000111010011011000110101;
    rom[35125] = 25'b0000111010010000010101110;
    rom[35126] = 25'b0000111010000101100101010;
    rom[35127] = 25'b0000111001111010110101000;
    rom[35128] = 25'b0000111001110000000101001;
    rom[35129] = 25'b0000111001100101010101011;
    rom[35130] = 25'b0000111001011010100110000;
    rom[35131] = 25'b0000111001001111110111000;
    rom[35132] = 25'b0000111001000101001000010;
    rom[35133] = 25'b0000111000111010011001111;
    rom[35134] = 25'b0000111000101111101011110;
    rom[35135] = 25'b0000111000100100111101111;
    rom[35136] = 25'b0000111000011010010000011;
    rom[35137] = 25'b0000111000001111100011010;
    rom[35138] = 25'b0000111000000100110110011;
    rom[35139] = 25'b0000110111111010001001110;
    rom[35140] = 25'b0000110111101111011101100;
    rom[35141] = 25'b0000110111100100110001100;
    rom[35142] = 25'b0000110111011010000101111;
    rom[35143] = 25'b0000110111001111011010100;
    rom[35144] = 25'b0000110111000100101111100;
    rom[35145] = 25'b0000110110111010000100110;
    rom[35146] = 25'b0000110110101111011010011;
    rom[35147] = 25'b0000110110100100110000010;
    rom[35148] = 25'b0000110110011010000110011;
    rom[35149] = 25'b0000110110001111011101000;
    rom[35150] = 25'b0000110110000100110011111;
    rom[35151] = 25'b0000110101111010001011000;
    rom[35152] = 25'b0000110101101111100010011;
    rom[35153] = 25'b0000110101100100111010010;
    rom[35154] = 25'b0000110101011010010010011;
    rom[35155] = 25'b0000110101001111101010110;
    rom[35156] = 25'b0000110101000101000011100;
    rom[35157] = 25'b0000110100111010011100100;
    rom[35158] = 25'b0000110100101111110101111;
    rom[35159] = 25'b0000110100100101001111101;
    rom[35160] = 25'b0000110100011010101001101;
    rom[35161] = 25'b0000110100010000000011111;
    rom[35162] = 25'b0000110100000101011110100;
    rom[35163] = 25'b0000110011111010111001100;
    rom[35164] = 25'b0000110011110000010100110;
    rom[35165] = 25'b0000110011100101110000011;
    rom[35166] = 25'b0000110011011011001100010;
    rom[35167] = 25'b0000110011010000101000100;
    rom[35168] = 25'b0000110011000110000101000;
    rom[35169] = 25'b0000110010111011100001111;
    rom[35170] = 25'b0000110010110000111111001;
    rom[35171] = 25'b0000110010100110011100101;
    rom[35172] = 25'b0000110010011011111010100;
    rom[35173] = 25'b0000110010010001011000101;
    rom[35174] = 25'b0000110010000110110111001;
    rom[35175] = 25'b0000110001111100010110000;
    rom[35176] = 25'b0000110001110001110101001;
    rom[35177] = 25'b0000110001100111010100100;
    rom[35178] = 25'b0000110001011100110100011;
    rom[35179] = 25'b0000110001010010010100011;
    rom[35180] = 25'b0000110001000111110100111;
    rom[35181] = 25'b0000110000111101010101101;
    rom[35182] = 25'b0000110000110010110110110;
    rom[35183] = 25'b0000110000101000011000001;
    rom[35184] = 25'b0000110000011101111001111;
    rom[35185] = 25'b0000110000010011011011111;
    rom[35186] = 25'b0000110000001000111110011;
    rom[35187] = 25'b0000101111111110100001000;
    rom[35188] = 25'b0000101111110100000100001;
    rom[35189] = 25'b0000101111101001100111100;
    rom[35190] = 25'b0000101111011111001011001;
    rom[35191] = 25'b0000101111010100101111010;
    rom[35192] = 25'b0000101111001010010011101;
    rom[35193] = 25'b0000101110111111111000010;
    rom[35194] = 25'b0000101110110101011101011;
    rom[35195] = 25'b0000101110101011000010110;
    rom[35196] = 25'b0000101110100000101000011;
    rom[35197] = 25'b0000101110010110001110100;
    rom[35198] = 25'b0000101110001011110100110;
    rom[35199] = 25'b0000101110000001011011100;
    rom[35200] = 25'b0000101101110111000010101;
    rom[35201] = 25'b0000101101101100101010000;
    rom[35202] = 25'b0000101101100010010001101;
    rom[35203] = 25'b0000101101010111111001101;
    rom[35204] = 25'b0000101101001101100010000;
    rom[35205] = 25'b0000101101000011001010110;
    rom[35206] = 25'b0000101100111000110011111;
    rom[35207] = 25'b0000101100101110011101001;
    rom[35208] = 25'b0000101100100100000110111;
    rom[35209] = 25'b0000101100011001110000111;
    rom[35210] = 25'b0000101100001111011011010;
    rom[35211] = 25'b0000101100000101000110000;
    rom[35212] = 25'b0000101011111010110001001;
    rom[35213] = 25'b0000101011110000011100100;
    rom[35214] = 25'b0000101011100110001000010;
    rom[35215] = 25'b0000101011011011110100011;
    rom[35216] = 25'b0000101011010001100000110;
    rom[35217] = 25'b0000101011000111001101100;
    rom[35218] = 25'b0000101010111100111010101;
    rom[35219] = 25'b0000101010110010101000000;
    rom[35220] = 25'b0000101010101000010101111;
    rom[35221] = 25'b0000101010011110000100000;
    rom[35222] = 25'b0000101010010011110010100;
    rom[35223] = 25'b0000101010001001100001011;
    rom[35224] = 25'b0000101001111111010000100;
    rom[35225] = 25'b0000101001110101000000000;
    rom[35226] = 25'b0000101001101010101111110;
    rom[35227] = 25'b0000101001100000100000000;
    rom[35228] = 25'b0000101001010110010000101;
    rom[35229] = 25'b0000101001001100000001011;
    rom[35230] = 25'b0000101001000001110010101;
    rom[35231] = 25'b0000101000110111100100001;
    rom[35232] = 25'b0000101000101101010110001;
    rom[35233] = 25'b0000101000100011001000011;
    rom[35234] = 25'b0000101000011000111011000;
    rom[35235] = 25'b0000101000001110101110000;
    rom[35236] = 25'b0000101000000100100001010;
    rom[35237] = 25'b0000100111111010010100111;
    rom[35238] = 25'b0000100111110000001000111;
    rom[35239] = 25'b0000100111100101111101010;
    rom[35240] = 25'b0000100111011011110010000;
    rom[35241] = 25'b0000100111010001100111000;
    rom[35242] = 25'b0000100111000111011100011;
    rom[35243] = 25'b0000100110111101010010001;
    rom[35244] = 25'b0000100110110011001000010;
    rom[35245] = 25'b0000100110101000111110101;
    rom[35246] = 25'b0000100110011110110101100;
    rom[35247] = 25'b0000100110010100101100101;
    rom[35248] = 25'b0000100110001010100100010;
    rom[35249] = 25'b0000100110000000011100000;
    rom[35250] = 25'b0000100101110110010100010;
    rom[35251] = 25'b0000100101101100001100111;
    rom[35252] = 25'b0000100101100010000101110;
    rom[35253] = 25'b0000100101010111111111000;
    rom[35254] = 25'b0000100101001101111000101;
    rom[35255] = 25'b0000100101000011110010100;
    rom[35256] = 25'b0000100100111001101101000;
    rom[35257] = 25'b0000100100101111100111101;
    rom[35258] = 25'b0000100100100101100010101;
    rom[35259] = 25'b0000100100011011011110001;
    rom[35260] = 25'b0000100100010001011001111;
    rom[35261] = 25'b0000100100000111010110000;
    rom[35262] = 25'b0000100011111101010010100;
    rom[35263] = 25'b0000100011110011001111010;
    rom[35264] = 25'b0000100011101001001100100;
    rom[35265] = 25'b0000100011011111001010000;
    rom[35266] = 25'b0000100011010101000111111;
    rom[35267] = 25'b0000100011001011000110001;
    rom[35268] = 25'b0000100011000001000100111;
    rom[35269] = 25'b0000100010110111000011111;
    rom[35270] = 25'b0000100010101101000011001;
    rom[35271] = 25'b0000100010100011000010111;
    rom[35272] = 25'b0000100010011001000011000;
    rom[35273] = 25'b0000100010001111000011011;
    rom[35274] = 25'b0000100010000101000100001;
    rom[35275] = 25'b0000100001111011000101011;
    rom[35276] = 25'b0000100001110001000110111;
    rom[35277] = 25'b0000100001100111001000110;
    rom[35278] = 25'b0000100001011101001010111;
    rom[35279] = 25'b0000100001010011001101100;
    rom[35280] = 25'b0000100001001001010000101;
    rom[35281] = 25'b0000100000111111010011111;
    rom[35282] = 25'b0000100000110101010111101;
    rom[35283] = 25'b0000100000101011011011101;
    rom[35284] = 25'b0000100000100001100000000;
    rom[35285] = 25'b0000100000010111100100111;
    rom[35286] = 25'b0000100000001101101010001;
    rom[35287] = 25'b0000100000000011101111101;
    rom[35288] = 25'b0000011111111001110101100;
    rom[35289] = 25'b0000011111101111111011110;
    rom[35290] = 25'b0000011111100110000010011;
    rom[35291] = 25'b0000011111011100001001011;
    rom[35292] = 25'b0000011111010010010000110;
    rom[35293] = 25'b0000011111001000011000100;
    rom[35294] = 25'b0000011110111110100000101;
    rom[35295] = 25'b0000011110110100101001001;
    rom[35296] = 25'b0000011110101010110001111;
    rom[35297] = 25'b0000011110100000111011001;
    rom[35298] = 25'b0000011110010111000100110;
    rom[35299] = 25'b0000011110001101001110110;
    rom[35300] = 25'b0000011110000011011001000;
    rom[35301] = 25'b0000011101111001100011101;
    rom[35302] = 25'b0000011101101111101110110;
    rom[35303] = 25'b0000011101100101111010010;
    rom[35304] = 25'b0000011101011100000110000;
    rom[35305] = 25'b0000011101010010010010010;
    rom[35306] = 25'b0000011101001000011110110;
    rom[35307] = 25'b0000011100111110101011110;
    rom[35308] = 25'b0000011100110100111001001;
    rom[35309] = 25'b0000011100101011000110110;
    rom[35310] = 25'b0000011100100001010100110;
    rom[35311] = 25'b0000011100010111100011010;
    rom[35312] = 25'b0000011100001101110010000;
    rom[35313] = 25'b0000011100000100000001010;
    rom[35314] = 25'b0000011011111010010000110;
    rom[35315] = 25'b0000011011110000100000110;
    rom[35316] = 25'b0000011011100110110001000;
    rom[35317] = 25'b0000011011011101000001110;
    rom[35318] = 25'b0000011011010011010010110;
    rom[35319] = 25'b0000011011001001100100010;
    rom[35320] = 25'b0000011010111111110110001;
    rom[35321] = 25'b0000011010110110001000010;
    rom[35322] = 25'b0000011010101100011010111;
    rom[35323] = 25'b0000011010100010101101111;
    rom[35324] = 25'b0000011010011001000001001;
    rom[35325] = 25'b0000011010001111010100111;
    rom[35326] = 25'b0000011010000101101001000;
    rom[35327] = 25'b0000011001111011111101100;
    rom[35328] = 25'b0000011001110010010010011;
    rom[35329] = 25'b0000011001101000100111101;
    rom[35330] = 25'b0000011001011110111101010;
    rom[35331] = 25'b0000011001010101010011010;
    rom[35332] = 25'b0000011001001011101001101;
    rom[35333] = 25'b0000011001000010000000011;
    rom[35334] = 25'b0000011000111000010111101;
    rom[35335] = 25'b0000011000101110101111000;
    rom[35336] = 25'b0000011000100101000111000;
    rom[35337] = 25'b0000011000011011011111011;
    rom[35338] = 25'b0000011000010001111000000;
    rom[35339] = 25'b0000011000001000010001001;
    rom[35340] = 25'b0000010111111110101010101;
    rom[35341] = 25'b0000010111110101000100011;
    rom[35342] = 25'b0000010111101011011110101;
    rom[35343] = 25'b0000010111100001111001010;
    rom[35344] = 25'b0000010111011000010100010;
    rom[35345] = 25'b0000010111001110101111110;
    rom[35346] = 25'b0000010111000101001011100;
    rom[35347] = 25'b0000010110111011100111101;
    rom[35348] = 25'b0000010110110010000100001;
    rom[35349] = 25'b0000010110101000100001001;
    rom[35350] = 25'b0000010110011110111110100;
    rom[35351] = 25'b0000010110010101011100010;
    rom[35352] = 25'b0000010110001011111010010;
    rom[35353] = 25'b0000010110000010011000110;
    rom[35354] = 25'b0000010101111000110111101;
    rom[35355] = 25'b0000010101101111010111000;
    rom[35356] = 25'b0000010101100101110110101;
    rom[35357] = 25'b0000010101011100010110110;
    rom[35358] = 25'b0000010101010010110111001;
    rom[35359] = 25'b0000010101001001010111111;
    rom[35360] = 25'b0000010100111111111001010;
    rom[35361] = 25'b0000010100110110011010111;
    rom[35362] = 25'b0000010100101100111100111;
    rom[35363] = 25'b0000010100100011011111010;
    rom[35364] = 25'b0000010100011010000010001;
    rom[35365] = 25'b0000010100010000100101010;
    rom[35366] = 25'b0000010100000111001000111;
    rom[35367] = 25'b0000010011111101101100110;
    rom[35368] = 25'b0000010011110100010001010;
    rom[35369] = 25'b0000010011101010110110000;
    rom[35370] = 25'b0000010011100001011011001;
    rom[35371] = 25'b0000010011011000000000110;
    rom[35372] = 25'b0000010011001110100110101;
    rom[35373] = 25'b0000010011000101001101000;
    rom[35374] = 25'b0000010010111011110011110;
    rom[35375] = 25'b0000010010110010011011000;
    rom[35376] = 25'b0000010010101001000010100;
    rom[35377] = 25'b0000010010011111101010011;
    rom[35378] = 25'b0000010010010110010010110;
    rom[35379] = 25'b0000010010001100111011100;
    rom[35380] = 25'b0000010010000011100100101;
    rom[35381] = 25'b0000010001111010001110001;
    rom[35382] = 25'b0000010001110000111000001;
    rom[35383] = 25'b0000010001100111100010011;
    rom[35384] = 25'b0000010001011110001101001;
    rom[35385] = 25'b0000010001010100111000010;
    rom[35386] = 25'b0000010001001011100011111;
    rom[35387] = 25'b0000010001000010001111110;
    rom[35388] = 25'b0000010000111000111100001;
    rom[35389] = 25'b0000010000101111101000110;
    rom[35390] = 25'b0000010000100110010101111;
    rom[35391] = 25'b0000010000011101000011100;
    rom[35392] = 25'b0000010000010011110001011;
    rom[35393] = 25'b0000010000001010011111110;
    rom[35394] = 25'b0000010000000001001110100;
    rom[35395] = 25'b0000001111110111111101101;
    rom[35396] = 25'b0000001111101110101101001;
    rom[35397] = 25'b0000001111100101011101001;
    rom[35398] = 25'b0000001111011100001101100;
    rom[35399] = 25'b0000001111010010111110010;
    rom[35400] = 25'b0000001111001001101111011;
    rom[35401] = 25'b0000001111000000100001000;
    rom[35402] = 25'b0000001110110111010011000;
    rom[35403] = 25'b0000001110101110000101010;
    rom[35404] = 25'b0000001110100100111000001;
    rom[35405] = 25'b0000001110011011101011011;
    rom[35406] = 25'b0000001110010010011110111;
    rom[35407] = 25'b0000001110001001010010111;
    rom[35408] = 25'b0000001110000000000111011;
    rom[35409] = 25'b0000001101110110111100001;
    rom[35410] = 25'b0000001101101101110001011;
    rom[35411] = 25'b0000001101100100100111000;
    rom[35412] = 25'b0000001101011011011101000;
    rom[35413] = 25'b0000001101010010010011100;
    rom[35414] = 25'b0000001101001001001010010;
    rom[35415] = 25'b0000001101000000000001101;
    rom[35416] = 25'b0000001100110110111001010;
    rom[35417] = 25'b0000001100101101110001011;
    rom[35418] = 25'b0000001100100100101001111;
    rom[35419] = 25'b0000001100011011100010110;
    rom[35420] = 25'b0000001100010010011100001;
    rom[35421] = 25'b0000001100001001010101111;
    rom[35422] = 25'b0000001100000000001111111;
    rom[35423] = 25'b0000001011110111001010100;
    rom[35424] = 25'b0000001011101110000101100;
    rom[35425] = 25'b0000001011100101000000110;
    rom[35426] = 25'b0000001011011011111100100;
    rom[35427] = 25'b0000001011010010111000110;
    rom[35428] = 25'b0000001011001001110101011;
    rom[35429] = 25'b0000001011000000110010011;
    rom[35430] = 25'b0000001010110111101111111;
    rom[35431] = 25'b0000001010101110101101110;
    rom[35432] = 25'b0000001010100101101100000;
    rom[35433] = 25'b0000001010011100101010101;
    rom[35434] = 25'b0000001010010011101001110;
    rom[35435] = 25'b0000001010001010101001010;
    rom[35436] = 25'b0000001010000001101001010;
    rom[35437] = 25'b0000001001111000101001100;
    rom[35438] = 25'b0000001001101111101010010;
    rom[35439] = 25'b0000001001100110101011011;
    rom[35440] = 25'b0000001001011101101101000;
    rom[35441] = 25'b0000001001010100101111000;
    rom[35442] = 25'b0000001001001011110001100;
    rom[35443] = 25'b0000001001000010110100011;
    rom[35444] = 25'b0000001000111001110111101;
    rom[35445] = 25'b0000001000110000111011010;
    rom[35446] = 25'b0000001000100111111111011;
    rom[35447] = 25'b0000001000011111000011110;
    rom[35448] = 25'b0000001000010110001000110;
    rom[35449] = 25'b0000001000001101001110001;
    rom[35450] = 25'b0000001000000100010011111;
    rom[35451] = 25'b0000000111111011011010000;
    rom[35452] = 25'b0000000111110010100000101;
    rom[35453] = 25'b0000000111101001100111101;
    rom[35454] = 25'b0000000111100000101111001;
    rom[35455] = 25'b0000000111010111110111000;
    rom[35456] = 25'b0000000111001110111111010;
    rom[35457] = 25'b0000000111000110001000000;
    rom[35458] = 25'b0000000110111101010001001;
    rom[35459] = 25'b0000000110110100011010101;
    rom[35460] = 25'b0000000110101011100100101;
    rom[35461] = 25'b0000000110100010101111000;
    rom[35462] = 25'b0000000110011001111001111;
    rom[35463] = 25'b0000000110010001000101001;
    rom[35464] = 25'b0000000110001000010000110;
    rom[35465] = 25'b0000000101111111011100111;
    rom[35466] = 25'b0000000101110110101001011;
    rom[35467] = 25'b0000000101101101110110010;
    rom[35468] = 25'b0000000101100101000011110;
    rom[35469] = 25'b0000000101011100010001100;
    rom[35470] = 25'b0000000101010011011111110;
    rom[35471] = 25'b0000000101001010101110010;
    rom[35472] = 25'b0000000101000001111101011;
    rom[35473] = 25'b0000000100111001001100111;
    rom[35474] = 25'b0000000100110000011100110;
    rom[35475] = 25'b0000000100100111101101001;
    rom[35476] = 25'b0000000100011110111101111;
    rom[35477] = 25'b0000000100010110001111001;
    rom[35478] = 25'b0000000100001101100000110;
    rom[35479] = 25'b0000000100000100110010111;
    rom[35480] = 25'b0000000011111100000101010;
    rom[35481] = 25'b0000000011110011011000001;
    rom[35482] = 25'b0000000011101010101011100;
    rom[35483] = 25'b0000000011100001111111010;
    rom[35484] = 25'b0000000011011001010011011;
    rom[35485] = 25'b0000000011010000101000000;
    rom[35486] = 25'b0000000011000111111101001;
    rom[35487] = 25'b0000000010111111010010101;
    rom[35488] = 25'b0000000010110110101000100;
    rom[35489] = 25'b0000000010101101111110111;
    rom[35490] = 25'b0000000010100101010101101;
    rom[35491] = 25'b0000000010011100101100110;
    rom[35492] = 25'b0000000010010100000100011;
    rom[35493] = 25'b0000000010001011011100100;
    rom[35494] = 25'b0000000010000010110101000;
    rom[35495] = 25'b0000000001111010001110000;
    rom[35496] = 25'b0000000001110001100111010;
    rom[35497] = 25'b0000000001101001000001001;
    rom[35498] = 25'b0000000001100000011011010;
    rom[35499] = 25'b0000000001010111110101111;
    rom[35500] = 25'b0000000001001111010001000;
    rom[35501] = 25'b0000000001000110101100100;
    rom[35502] = 25'b0000000000111110001000100;
    rom[35503] = 25'b0000000000110101100100111;
    rom[35504] = 25'b0000000000101101000001101;
    rom[35505] = 25'b0000000000100100011111000;
    rom[35506] = 25'b0000000000011011111100101;
    rom[35507] = 25'b0000000000010011011010110;
    rom[35508] = 25'b0000000000001010111001011;
    rom[35509] = 25'b0000000000000010011000011;
    rom[35510] = 25'b1111111111111001110111110;
    rom[35511] = 25'b1111111111110001010111110;
    rom[35512] = 25'b1111111111101000111000000;
    rom[35513] = 25'b1111111111100000011000110;
    rom[35514] = 25'b1111111111010111111010000;
    rom[35515] = 25'b1111111111001111011011100;
    rom[35516] = 25'b1111111111000110111101101;
    rom[35517] = 25'b1111111110111110100000001;
    rom[35518] = 25'b1111111110110110000011000;
    rom[35519] = 25'b1111111110101101100110011;
    rom[35520] = 25'b1111111110100101001010001;
    rom[35521] = 25'b1111111110011100101110011;
    rom[35522] = 25'b1111111110010100010011000;
    rom[35523] = 25'b1111111110001011111000010;
    rom[35524] = 25'b1111111110000011011101110;
    rom[35525] = 25'b1111111101111011000011110;
    rom[35526] = 25'b1111111101110010101010010;
    rom[35527] = 25'b1111111101101010010001000;
    rom[35528] = 25'b1111111101100001111000011;
    rom[35529] = 25'b1111111101011001100000001;
    rom[35530] = 25'b1111111101010001001000011;
    rom[35531] = 25'b1111111101001000110001000;
    rom[35532] = 25'b1111111101000000011010000;
    rom[35533] = 25'b1111111100111000000011101;
    rom[35534] = 25'b1111111100101111101101100;
    rom[35535] = 25'b1111111100100111010111111;
    rom[35536] = 25'b1111111100011111000010110;
    rom[35537] = 25'b1111111100010110101110000;
    rom[35538] = 25'b1111111100001110011001110;
    rom[35539] = 25'b1111111100000110000101111;
    rom[35540] = 25'b1111111011111101110010100;
    rom[35541] = 25'b1111111011110101011111101;
    rom[35542] = 25'b1111111011101101001101001;
    rom[35543] = 25'b1111111011100100111011000;
    rom[35544] = 25'b1111111011011100101001100;
    rom[35545] = 25'b1111111011010100011000011;
    rom[35546] = 25'b1111111011001100000111100;
    rom[35547] = 25'b1111111011000011110111010;
    rom[35548] = 25'b1111111010111011100111100;
    rom[35549] = 25'b1111111010110011011000001;
    rom[35550] = 25'b1111111010101011001001001;
    rom[35551] = 25'b1111111010100010111010101;
    rom[35552] = 25'b1111111010011010101100101;
    rom[35553] = 25'b1111111010010010011111000;
    rom[35554] = 25'b1111111010001010010001111;
    rom[35555] = 25'b1111111010000010000101001;
    rom[35556] = 25'b1111111001111001111000111;
    rom[35557] = 25'b1111111001110001101101000;
    rom[35558] = 25'b1111111001101001100001101;
    rom[35559] = 25'b1111111001100001010110110;
    rom[35560] = 25'b1111111001011001001100010;
    rom[35561] = 25'b1111111001010001000010010;
    rom[35562] = 25'b1111111001001000111000110;
    rom[35563] = 25'b1111111001000000101111101;
    rom[35564] = 25'b1111111000111000100110111;
    rom[35565] = 25'b1111111000110000011110110;
    rom[35566] = 25'b1111111000101000010110111;
    rom[35567] = 25'b1111111000100000001111101;
    rom[35568] = 25'b1111111000011000001000101;
    rom[35569] = 25'b1111111000010000000010010;
    rom[35570] = 25'b1111111000000111111100010;
    rom[35571] = 25'b1111110111111111110110110;
    rom[35572] = 25'b1111110111110111110001110;
    rom[35573] = 25'b1111110111101111101101001;
    rom[35574] = 25'b1111110111100111101000111;
    rom[35575] = 25'b1111110111011111100101001;
    rom[35576] = 25'b1111110111010111100001111;
    rom[35577] = 25'b1111110111001111011111000;
    rom[35578] = 25'b1111110111000111011100110;
    rom[35579] = 25'b1111110110111111011010110;
    rom[35580] = 25'b1111110110110111011001010;
    rom[35581] = 25'b1111110110101111011000010;
    rom[35582] = 25'b1111110110100111010111110;
    rom[35583] = 25'b1111110110011111010111101;
    rom[35584] = 25'b1111110110010111011000000;
    rom[35585] = 25'b1111110110001111011000110;
    rom[35586] = 25'b1111110110000111011010000;
    rom[35587] = 25'b1111110101111111011011110;
    rom[35588] = 25'b1111110101110111011101111;
    rom[35589] = 25'b1111110101101111100000100;
    rom[35590] = 25'b1111110101100111100011101;
    rom[35591] = 25'b1111110101011111100111001;
    rom[35592] = 25'b1111110101010111101011001;
    rom[35593] = 25'b1111110101001111101111100;
    rom[35594] = 25'b1111110101000111110100011;
    rom[35595] = 25'b1111110100111111111001110;
    rom[35596] = 25'b1111110100110111111111100;
    rom[35597] = 25'b1111110100110000000101110;
    rom[35598] = 25'b1111110100101000001100100;
    rom[35599] = 25'b1111110100100000010011110;
    rom[35600] = 25'b1111110100011000011011011;
    rom[35601] = 25'b1111110100010000100011011;
    rom[35602] = 25'b1111110100001000101100000;
    rom[35603] = 25'b1111110100000000110101000;
    rom[35604] = 25'b1111110011111000111110100;
    rom[35605] = 25'b1111110011110001001000010;
    rom[35606] = 25'b1111110011101001010010110;
    rom[35607] = 25'b1111110011100001011101100;
    rom[35608] = 25'b1111110011011001101000111;
    rom[35609] = 25'b1111110011010001110100101;
    rom[35610] = 25'b1111110011001010000000110;
    rom[35611] = 25'b1111110011000010001101100;
    rom[35612] = 25'b1111110010111010011010101;
    rom[35613] = 25'b1111110010110010101000001;
    rom[35614] = 25'b1111110010101010110110010;
    rom[35615] = 25'b1111110010100011000100110;
    rom[35616] = 25'b1111110010011011010011110;
    rom[35617] = 25'b1111110010010011100011001;
    rom[35618] = 25'b1111110010001011110011000;
    rom[35619] = 25'b1111110010000100000011011;
    rom[35620] = 25'b1111110001111100010100010;
    rom[35621] = 25'b1111110001110100100101100;
    rom[35622] = 25'b1111110001101100110111001;
    rom[35623] = 25'b1111110001100101001001011;
    rom[35624] = 25'b1111110001011101011100000;
    rom[35625] = 25'b1111110001010101101111001;
    rom[35626] = 25'b1111110001001110000010110;
    rom[35627] = 25'b1111110001000110010110110;
    rom[35628] = 25'b1111110000111110101011010;
    rom[35629] = 25'b1111110000110111000000010;
    rom[35630] = 25'b1111110000101111010101101;
    rom[35631] = 25'b1111110000100111101011101;
    rom[35632] = 25'b1111110000100000000010000;
    rom[35633] = 25'b1111110000011000011000110;
    rom[35634] = 25'b1111110000010000110000001;
    rom[35635] = 25'b1111110000001001000111110;
    rom[35636] = 25'b1111110000000001100000000;
    rom[35637] = 25'b1111101111111001111000110;
    rom[35638] = 25'b1111101111110010010001110;
    rom[35639] = 25'b1111101111101010101011100;
    rom[35640] = 25'b1111101111100011000101100;
    rom[35641] = 25'b1111101111011011100000000;
    rom[35642] = 25'b1111101111010011111011001;
    rom[35643] = 25'b1111101111001100010110100;
    rom[35644] = 25'b1111101111000100110010100;
    rom[35645] = 25'b1111101110111101001110111;
    rom[35646] = 25'b1111101110110101101011110;
    rom[35647] = 25'b1111101110101110001001001;
    rom[35648] = 25'b1111101110100110100110111;
    rom[35649] = 25'b1111101110011111000101001;
    rom[35650] = 25'b1111101110010111100011111;
    rom[35651] = 25'b1111101110010000000011001;
    rom[35652] = 25'b1111101110001000100010110;
    rom[35653] = 25'b1111101110000001000010111;
    rom[35654] = 25'b1111101101111001100011011;
    rom[35655] = 25'b1111101101110010000100100;
    rom[35656] = 25'b1111101101101010100110001;
    rom[35657] = 25'b1111101101100011001000001;
    rom[35658] = 25'b1111101101011011101010101;
    rom[35659] = 25'b1111101101010100001101100;
    rom[35660] = 25'b1111101101001100110000111;
    rom[35661] = 25'b1111101101000101010100111;
    rom[35662] = 25'b1111101100111101111001001;
    rom[35663] = 25'b1111101100110110011110000;
    rom[35664] = 25'b1111101100101111000011010;
    rom[35665] = 25'b1111101100100111101001000;
    rom[35666] = 25'b1111101100100000001111010;
    rom[35667] = 25'b1111101100011000110101111;
    rom[35668] = 25'b1111101100010001011101001;
    rom[35669] = 25'b1111101100001010000100110;
    rom[35670] = 25'b1111101100000010101100111;
    rom[35671] = 25'b1111101011111011010101100;
    rom[35672] = 25'b1111101011110011111110100;
    rom[35673] = 25'b1111101011101100101000000;
    rom[35674] = 25'b1111101011100101010010000;
    rom[35675] = 25'b1111101011011101111100100;
    rom[35676] = 25'b1111101011010110100111100;
    rom[35677] = 25'b1111101011001111010010111;
    rom[35678] = 25'b1111101011000111111110110;
    rom[35679] = 25'b1111101011000000101011001;
    rom[35680] = 25'b1111101010111001010111111;
    rom[35681] = 25'b1111101010110010000101010;
    rom[35682] = 25'b1111101010101010110011000;
    rom[35683] = 25'b1111101010100011100001010;
    rom[35684] = 25'b1111101010011100010000000;
    rom[35685] = 25'b1111101010010100111111001;
    rom[35686] = 25'b1111101010001101101110110;
    rom[35687] = 25'b1111101010000110011110111;
    rom[35688] = 25'b1111101001111111001111100;
    rom[35689] = 25'b1111101001111000000000101;
    rom[35690] = 25'b1111101001110000110010001;
    rom[35691] = 25'b1111101001101001100100001;
    rom[35692] = 25'b1111101001100010010110110;
    rom[35693] = 25'b1111101001011011001001110;
    rom[35694] = 25'b1111101001010011111101010;
    rom[35695] = 25'b1111101001001100110001001;
    rom[35696] = 25'b1111101001000101100101100;
    rom[35697] = 25'b1111101000111110011010011;
    rom[35698] = 25'b1111101000110111001111110;
    rom[35699] = 25'b1111101000110000000101101;
    rom[35700] = 25'b1111101000101000111011111;
    rom[35701] = 25'b1111101000100001110010101;
    rom[35702] = 25'b1111101000011010101001111;
    rom[35703] = 25'b1111101000010011100001110;
    rom[35704] = 25'b1111101000001100011001111;
    rom[35705] = 25'b1111101000000101010010101;
    rom[35706] = 25'b1111100111111110001011110;
    rom[35707] = 25'b1111100111110111000101011;
    rom[35708] = 25'b1111100111101111111111100;
    rom[35709] = 25'b1111100111101000111010001;
    rom[35710] = 25'b1111100111100001110101010;
    rom[35711] = 25'b1111100111011010110000110;
    rom[35712] = 25'b1111100111010011101100110;
    rom[35713] = 25'b1111100111001100101001010;
    rom[35714] = 25'b1111100111000101100110010;
    rom[35715] = 25'b1111100110111110100011110;
    rom[35716] = 25'b1111100110110111100001101;
    rom[35717] = 25'b1111100110110000100000001;
    rom[35718] = 25'b1111100110101001011111000;
    rom[35719] = 25'b1111100110100010011110011;
    rom[35720] = 25'b1111100110011011011110010;
    rom[35721] = 25'b1111100110010100011110101;
    rom[35722] = 25'b1111100110001101011111011;
    rom[35723] = 25'b1111100110000110100000110;
    rom[35724] = 25'b1111100101111111100010100;
    rom[35725] = 25'b1111100101111000100100110;
    rom[35726] = 25'b1111100101110001100111100;
    rom[35727] = 25'b1111100101101010101010101;
    rom[35728] = 25'b1111100101100011101110011;
    rom[35729] = 25'b1111100101011100110010101;
    rom[35730] = 25'b1111100101010101110111001;
    rom[35731] = 25'b1111100101001110111100011;
    rom[35732] = 25'b1111100101001000000010000;
    rom[35733] = 25'b1111100101000001001000000;
    rom[35734] = 25'b1111100100111010001110101;
    rom[35735] = 25'b1111100100110011010101110;
    rom[35736] = 25'b1111100100101100011101010;
    rom[35737] = 25'b1111100100100101100101010;
    rom[35738] = 25'b1111100100011110101101110;
    rom[35739] = 25'b1111100100010111110110110;
    rom[35740] = 25'b1111100100010001000000010;
    rom[35741] = 25'b1111100100001010001010001;
    rom[35742] = 25'b1111100100000011010100101;
    rom[35743] = 25'b1111100011111100011111100;
    rom[35744] = 25'b1111100011110101101010111;
    rom[35745] = 25'b1111100011101110110110110;
    rom[35746] = 25'b1111100011101000000011001;
    rom[35747] = 25'b1111100011100001010000000;
    rom[35748] = 25'b1111100011011010011101011;
    rom[35749] = 25'b1111100011010011101011001;
    rom[35750] = 25'b1111100011001100111001100;
    rom[35751] = 25'b1111100011000110001000010;
    rom[35752] = 25'b1111100010111111010111100;
    rom[35753] = 25'b1111100010111000100111010;
    rom[35754] = 25'b1111100010110001110111100;
    rom[35755] = 25'b1111100010101011001000010;
    rom[35756] = 25'b1111100010100100011001011;
    rom[35757] = 25'b1111100010011101101011001;
    rom[35758] = 25'b1111100010010110111101010;
    rom[35759] = 25'b1111100010010000010000000;
    rom[35760] = 25'b1111100010001001100011000;
    rom[35761] = 25'b1111100010000010110110101;
    rom[35762] = 25'b1111100001111100001010110;
    rom[35763] = 25'b1111100001110101011111011;
    rom[35764] = 25'b1111100001101110110100100;
    rom[35765] = 25'b1111100001101000001010000;
    rom[35766] = 25'b1111100001100001100000000;
    rom[35767] = 25'b1111100001011010110110101;
    rom[35768] = 25'b1111100001010100001101101;
    rom[35769] = 25'b1111100001001101100101001;
    rom[35770] = 25'b1111100001000110111101001;
    rom[35771] = 25'b1111100001000000010101101;
    rom[35772] = 25'b1111100000111001101110101;
    rom[35773] = 25'b1111100000110011001000000;
    rom[35774] = 25'b1111100000101100100010000;
    rom[35775] = 25'b1111100000100101111100011;
    rom[35776] = 25'b1111100000011111010111010;
    rom[35777] = 25'b1111100000011000110010110;
    rom[35778] = 25'b1111100000010010001110101;
    rom[35779] = 25'b1111100000001011101010111;
    rom[35780] = 25'b1111100000000101000111110;
    rom[35781] = 25'b1111011111111110100101001;
    rom[35782] = 25'b1111011111111000000011000;
    rom[35783] = 25'b1111011111110001100001010;
    rom[35784] = 25'b1111011111101011000000001;
    rom[35785] = 25'b1111011111100100011111100;
    rom[35786] = 25'b1111011111011101111111010;
    rom[35787] = 25'b1111011111010111011111100;
    rom[35788] = 25'b1111011111010001000000010;
    rom[35789] = 25'b1111011111001010100001100;
    rom[35790] = 25'b1111011111000100000011010;
    rom[35791] = 25'b1111011110111101100101100;
    rom[35792] = 25'b1111011110110111001000001;
    rom[35793] = 25'b1111011110110000101011011;
    rom[35794] = 25'b1111011110101010001111001;
    rom[35795] = 25'b1111011110100011110011010;
    rom[35796] = 25'b1111011110011101011000000;
    rom[35797] = 25'b1111011110010110111101001;
    rom[35798] = 25'b1111011110010000100010110;
    rom[35799] = 25'b1111011110001010001000111;
    rom[35800] = 25'b1111011110000011101111100;
    rom[35801] = 25'b1111011101111101010110101;
    rom[35802] = 25'b1111011101110110111110010;
    rom[35803] = 25'b1111011101110000100110011;
    rom[35804] = 25'b1111011101101010001110111;
    rom[35805] = 25'b1111011101100011111000000;
    rom[35806] = 25'b1111011101011101100001101;
    rom[35807] = 25'b1111011101010111001011101;
    rom[35808] = 25'b1111011101010000110110010;
    rom[35809] = 25'b1111011101001010100001010;
    rom[35810] = 25'b1111011101000100001100110;
    rom[35811] = 25'b1111011100111101111000110;
    rom[35812] = 25'b1111011100110111100101011;
    rom[35813] = 25'b1111011100110001010010011;
    rom[35814] = 25'b1111011100101010111111111;
    rom[35815] = 25'b1111011100100100101101111;
    rom[35816] = 25'b1111011100011110011100011;
    rom[35817] = 25'b1111011100011000001011010;
    rom[35818] = 25'b1111011100010001111010110;
    rom[35819] = 25'b1111011100001011101010110;
    rom[35820] = 25'b1111011100000101011011010;
    rom[35821] = 25'b1111011011111111001100001;
    rom[35822] = 25'b1111011011111000111101101;
    rom[35823] = 25'b1111011011110010101111100;
    rom[35824] = 25'b1111011011101100100001111;
    rom[35825] = 25'b1111011011100110010100111;
    rom[35826] = 25'b1111011011100000001000010;
    rom[35827] = 25'b1111011011011001111100001;
    rom[35828] = 25'b1111011011010011110000100;
    rom[35829] = 25'b1111011011001101100101011;
    rom[35830] = 25'b1111011011000111011010110;
    rom[35831] = 25'b1111011011000001010000101;
    rom[35832] = 25'b1111011010111011000111000;
    rom[35833] = 25'b1111011010110100111101111;
    rom[35834] = 25'b1111011010101110110101010;
    rom[35835] = 25'b1111011010101000101101000;
    rom[35836] = 25'b1111011010100010100101011;
    rom[35837] = 25'b1111011010011100011110010;
    rom[35838] = 25'b1111011010010110010111100;
    rom[35839] = 25'b1111011010010000010001011;
    rom[35840] = 25'b1111011010001010001011101;
    rom[35841] = 25'b1111011010000100000110100;
    rom[35842] = 25'b1111011001111110000001110;
    rom[35843] = 25'b1111011001110111111101100;
    rom[35844] = 25'b1111011001110001111001111;
    rom[35845] = 25'b1111011001101011110110101;
    rom[35846] = 25'b1111011001100101110011111;
    rom[35847] = 25'b1111011001011111110001101;
    rom[35848] = 25'b1111011001011001101111111;
    rom[35849] = 25'b1111011001010011101110110;
    rom[35850] = 25'b1111011001001101101110000;
    rom[35851] = 25'b1111011001000111101101101;
    rom[35852] = 25'b1111011001000001101110000;
    rom[35853] = 25'b1111011000111011101110101;
    rom[35854] = 25'b1111011000110101101111111;
    rom[35855] = 25'b1111011000101111110001101;
    rom[35856] = 25'b1111011000101001110011110;
    rom[35857] = 25'b1111011000100011110110101;
    rom[35858] = 25'b1111011000011101111001110;
    rom[35859] = 25'b1111011000010111111101100;
    rom[35860] = 25'b1111011000010010000001101;
    rom[35861] = 25'b1111011000001100000110011;
    rom[35862] = 25'b1111011000000110001011101;
    rom[35863] = 25'b1111011000000000010001010;
    rom[35864] = 25'b1111010111111010010111100;
    rom[35865] = 25'b1111010111110100011110001;
    rom[35866] = 25'b1111010111101110100101010;
    rom[35867] = 25'b1111010111101000101101000;
    rom[35868] = 25'b1111010111100010110101001;
    rom[35869] = 25'b1111010111011100111101111;
    rom[35870] = 25'b1111010111010111000111000;
    rom[35871] = 25'b1111010111010001010000110;
    rom[35872] = 25'b1111010111001011011010111;
    rom[35873] = 25'b1111010111000101100101100;
    rom[35874] = 25'b1111010110111111110000110;
    rom[35875] = 25'b1111010110111001111100011;
    rom[35876] = 25'b1111010110110100001000100;
    rom[35877] = 25'b1111010110101110010101001;
    rom[35878] = 25'b1111010110101000100010010;
    rom[35879] = 25'b1111010110100010101111111;
    rom[35880] = 25'b1111010110011100111110001;
    rom[35881] = 25'b1111010110010111001100101;
    rom[35882] = 25'b1111010110010001011011111;
    rom[35883] = 25'b1111010110001011101011100;
    rom[35884] = 25'b1111010110000101111011101;
    rom[35885] = 25'b1111010110000000001100010;
    rom[35886] = 25'b1111010101111010011101010;
    rom[35887] = 25'b1111010101110100101110111;
    rom[35888] = 25'b1111010101101111000001000;
    rom[35889] = 25'b1111010101101001010011110;
    rom[35890] = 25'b1111010101100011100110110;
    rom[35891] = 25'b1111010101011101111010011;
    rom[35892] = 25'b1111010101011000001110100;
    rom[35893] = 25'b1111010101010010100011001;
    rom[35894] = 25'b1111010101001100111000010;
    rom[35895] = 25'b1111010101000111001101111;
    rom[35896] = 25'b1111010101000001100100000;
    rom[35897] = 25'b1111010100111011111010100;
    rom[35898] = 25'b1111010100110110010001101;
    rom[35899] = 25'b1111010100110000101001010;
    rom[35900] = 25'b1111010100101011000001010;
    rom[35901] = 25'b1111010100100101011010000;
    rom[35902] = 25'b1111010100011111110011000;
    rom[35903] = 25'b1111010100011010001100101;
    rom[35904] = 25'b1111010100010100100110110;
    rom[35905] = 25'b1111010100001111000001010;
    rom[35906] = 25'b1111010100001001011100011;
    rom[35907] = 25'b1111010100000011111000000;
    rom[35908] = 25'b1111010011111110010100001;
    rom[35909] = 25'b1111010011111000110000101;
    rom[35910] = 25'b1111010011110011001101110;
    rom[35911] = 25'b1111010011101101101011010;
    rom[35912] = 25'b1111010011101000001001100;
    rom[35913] = 25'b1111010011100010101000000;
    rom[35914] = 25'b1111010011011101000111001;
    rom[35915] = 25'b1111010011010111100110110;
    rom[35916] = 25'b1111010011010010000110110;
    rom[35917] = 25'b1111010011001100100111011;
    rom[35918] = 25'b1111010011000111001000100;
    rom[35919] = 25'b1111010011000001101010000;
    rom[35920] = 25'b1111010010111100001100001;
    rom[35921] = 25'b1111010010110110101110110;
    rom[35922] = 25'b1111010010110001010001111;
    rom[35923] = 25'b1111010010101011110101011;
    rom[35924] = 25'b1111010010100110011001100;
    rom[35925] = 25'b1111010010100000111110000;
    rom[35926] = 25'b1111010010011011100011001;
    rom[35927] = 25'b1111010010010110001000110;
    rom[35928] = 25'b1111010010010000101110111;
    rom[35929] = 25'b1111010010001011010101011;
    rom[35930] = 25'b1111010010000101111100100;
    rom[35931] = 25'b1111010010000000100100001;
    rom[35932] = 25'b1111010001111011001100001;
    rom[35933] = 25'b1111010001110101110100110;
    rom[35934] = 25'b1111010001110000011101111;
    rom[35935] = 25'b1111010001101011000111011;
    rom[35936] = 25'b1111010001100101110001100;
    rom[35937] = 25'b1111010001100000011100001;
    rom[35938] = 25'b1111010001011011000111010;
    rom[35939] = 25'b1111010001010101110010110;
    rom[35940] = 25'b1111010001010000011110111;
    rom[35941] = 25'b1111010001001011001011100;
    rom[35942] = 25'b1111010001000101111000100;
    rom[35943] = 25'b1111010001000000100110010;
    rom[35944] = 25'b1111010000111011010100010;
    rom[35945] = 25'b1111010000110110000010111;
    rom[35946] = 25'b1111010000110000110010000;
    rom[35947] = 25'b1111010000101011100001101;
    rom[35948] = 25'b1111010000100110010001110;
    rom[35949] = 25'b1111010000100001000010010;
    rom[35950] = 25'b1111010000011011110011011;
    rom[35951] = 25'b1111010000010110100101000;
    rom[35952] = 25'b1111010000010001010111001;
    rom[35953] = 25'b1111010000001100001001110;
    rom[35954] = 25'b1111010000000110111100110;
    rom[35955] = 25'b1111010000000001110000011;
    rom[35956] = 25'b1111001111111100100100100;
    rom[35957] = 25'b1111001111110111011001001;
    rom[35958] = 25'b1111001111110010001110010;
    rom[35959] = 25'b1111001111101101000011111;
    rom[35960] = 25'b1111001111100111111010000;
    rom[35961] = 25'b1111001111100010110000101;
    rom[35962] = 25'b1111001111011101100111110;
    rom[35963] = 25'b1111001111011000011111011;
    rom[35964] = 25'b1111001111010011010111100;
    rom[35965] = 25'b1111001111001110010000001;
    rom[35966] = 25'b1111001111001001001001010;
    rom[35967] = 25'b1111001111000100000010111;
    rom[35968] = 25'b1111001110111110111101000;
    rom[35969] = 25'b1111001110111001110111110;
    rom[35970] = 25'b1111001110110100110010110;
    rom[35971] = 25'b1111001110101111101110100;
    rom[35972] = 25'b1111001110101010101010101;
    rom[35973] = 25'b1111001110100101100111010;
    rom[35974] = 25'b1111001110100000100100011;
    rom[35975] = 25'b1111001110011011100010000;
    rom[35976] = 25'b1111001110010110100000001;
    rom[35977] = 25'b1111001110010001011110111;
    rom[35978] = 25'b1111001110001100011110000;
    rom[35979] = 25'b1111001110000111011101101;
    rom[35980] = 25'b1111001110000010011101110;
    rom[35981] = 25'b1111001101111101011110100;
    rom[35982] = 25'b1111001101111000011111101;
    rom[35983] = 25'b1111001101110011100001011;
    rom[35984] = 25'b1111001101101110100011011;
    rom[35985] = 25'b1111001101101001100110001;
    rom[35986] = 25'b1111001101100100101001011;
    rom[35987] = 25'b1111001101011111101101000;
    rom[35988] = 25'b1111001101011010110001010;
    rom[35989] = 25'b1111001101010101110101111;
    rom[35990] = 25'b1111001101010000111011000;
    rom[35991] = 25'b1111001101001100000000101;
    rom[35992] = 25'b1111001101000111000110111;
    rom[35993] = 25'b1111001101000010001101101;
    rom[35994] = 25'b1111001100111101010100111;
    rom[35995] = 25'b1111001100111000011100100;
    rom[35996] = 25'b1111001100110011100100110;
    rom[35997] = 25'b1111001100101110101101011;
    rom[35998] = 25'b1111001100101001110110101;
    rom[35999] = 25'b1111001100100101000000011;
    rom[36000] = 25'b1111001100100000001010100;
    rom[36001] = 25'b1111001100011011010101010;
    rom[36002] = 25'b1111001100010110100000100;
    rom[36003] = 25'b1111001100010001101100001;
    rom[36004] = 25'b1111001100001100111000011;
    rom[36005] = 25'b1111001100001000000101001;
    rom[36006] = 25'b1111001100000011010010011;
    rom[36007] = 25'b1111001011111110100000000;
    rom[36008] = 25'b1111001011111001101110010;
    rom[36009] = 25'b1111001011110100111101000;
    rom[36010] = 25'b1111001011110000001100010;
    rom[36011] = 25'b1111001011101011011100000;
    rom[36012] = 25'b1111001011100110101100010;
    rom[36013] = 25'b1111001011100001111101000;
    rom[36014] = 25'b1111001011011101001110010;
    rom[36015] = 25'b1111001011011000100000000;
    rom[36016] = 25'b1111001011010011110010010;
    rom[36017] = 25'b1111001011001111000101001;
    rom[36018] = 25'b1111001011001010011000010;
    rom[36019] = 25'b1111001011000101101100000;
    rom[36020] = 25'b1111001011000001000000011;
    rom[36021] = 25'b1111001010111100010101000;
    rom[36022] = 25'b1111001010110111101010011;
    rom[36023] = 25'b1111001010110011000000001;
    rom[36024] = 25'b1111001010101110010110011;
    rom[36025] = 25'b1111001010101001101101010;
    rom[36026] = 25'b1111001010100101000100100;
    rom[36027] = 25'b1111001010100000011100010;
    rom[36028] = 25'b1111001010011011110100101;
    rom[36029] = 25'b1111001010010111001101011;
    rom[36030] = 25'b1111001010010010100110101;
    rom[36031] = 25'b1111001010001110000000100;
    rom[36032] = 25'b1111001010001001011010110;
    rom[36033] = 25'b1111001010000100110101100;
    rom[36034] = 25'b1111001010000000010000111;
    rom[36035] = 25'b1111001001111011101100101;
    rom[36036] = 25'b1111001001110111001001000;
    rom[36037] = 25'b1111001001110010100101111;
    rom[36038] = 25'b1111001001101110000011001;
    rom[36039] = 25'b1111001001101001100001000;
    rom[36040] = 25'b1111001001100100111111010;
    rom[36041] = 25'b1111001001100000011110001;
    rom[36042] = 25'b1111001001011011111101100;
    rom[36043] = 25'b1111001001010111011101010;
    rom[36044] = 25'b1111001001010010111101101;
    rom[36045] = 25'b1111001001001110011110100;
    rom[36046] = 25'b1111001001001001111111110;
    rom[36047] = 25'b1111001001000101100001101;
    rom[36048] = 25'b1111001001000001000100000;
    rom[36049] = 25'b1111001000111100100110111;
    rom[36050] = 25'b1111001000111000001010010;
    rom[36051] = 25'b1111001000110011101110000;
    rom[36052] = 25'b1111001000101111010010100;
    rom[36053] = 25'b1111001000101010110111010;
    rom[36054] = 25'b1111001000100110011100101;
    rom[36055] = 25'b1111001000100010000010100;
    rom[36056] = 25'b1111001000011101101000111;
    rom[36057] = 25'b1111001000011001001111110;
    rom[36058] = 25'b1111001000010100110111001;
    rom[36059] = 25'b1111001000010000011111000;
    rom[36060] = 25'b1111001000001100000111100;
    rom[36061] = 25'b1111001000000111110000010;
    rom[36062] = 25'b1111001000000011011001101;
    rom[36063] = 25'b1111000111111111000011100;
    rom[36064] = 25'b1111000111111010101110000;
    rom[36065] = 25'b1111000111110110011000111;
    rom[36066] = 25'b1111000111110010000100010;
    rom[36067] = 25'b1111000111101101110000001;
    rom[36068] = 25'b1111000111101001011100101;
    rom[36069] = 25'b1111000111100101001001100;
    rom[36070] = 25'b1111000111100000110110111;
    rom[36071] = 25'b1111000111011100100100110;
    rom[36072] = 25'b1111000111011000010011001;
    rom[36073] = 25'b1111000111010100000010001;
    rom[36074] = 25'b1111000111001111110001100;
    rom[36075] = 25'b1111000111001011100001100;
    rom[36076] = 25'b1111000111000111010001111;
    rom[36077] = 25'b1111000111000011000010110;
    rom[36078] = 25'b1111000110111110110100010;
    rom[36079] = 25'b1111000110111010100110010;
    rom[36080] = 25'b1111000110110110011000101;
    rom[36081] = 25'b1111000110110010001011100;
    rom[36082] = 25'b1111000110101101111111000;
    rom[36083] = 25'b1111000110101001110010111;
    rom[36084] = 25'b1111000110100101100111011;
    rom[36085] = 25'b1111000110100001011100011;
    rom[36086] = 25'b1111000110011101010001110;
    rom[36087] = 25'b1111000110011001000111110;
    rom[36088] = 25'b1111000110010100111110010;
    rom[36089] = 25'b1111000110010000110101001;
    rom[36090] = 25'b1111000110001100101100101;
    rom[36091] = 25'b1111000110001000100100101;
    rom[36092] = 25'b1111000110000100011101001;
    rom[36093] = 25'b1111000110000000010110000;
    rom[36094] = 25'b1111000101111100001111100;
    rom[36095] = 25'b1111000101111000001001100;
    rom[36096] = 25'b1111000101110100000011111;
    rom[36097] = 25'b1111000101101111111110111;
    rom[36098] = 25'b1111000101101011111010011;
    rom[36099] = 25'b1111000101100111110110010;
    rom[36100] = 25'b1111000101100011110010110;
    rom[36101] = 25'b1111000101011111101111111;
    rom[36102] = 25'b1111000101011011101101010;
    rom[36103] = 25'b1111000101010111101011010;
    rom[36104] = 25'b1111000101010011101001110;
    rom[36105] = 25'b1111000101001111101000110;
    rom[36106] = 25'b1111000101001011101000010;
    rom[36107] = 25'b1111000101000111101000010;
    rom[36108] = 25'b1111000101000011101000110;
    rom[36109] = 25'b1111000100111111101001101;
    rom[36110] = 25'b1111000100111011101011010;
    rom[36111] = 25'b1111000100110111101101001;
    rom[36112] = 25'b1111000100110011101111101;
    rom[36113] = 25'b1111000100101111110010101;
    rom[36114] = 25'b1111000100101011110110001;
    rom[36115] = 25'b1111000100100111111010001;
    rom[36116] = 25'b1111000100100011111110110;
    rom[36117] = 25'b1111000100100000000011101;
    rom[36118] = 25'b1111000100011100001001010;
    rom[36119] = 25'b1111000100011000001111010;
    rom[36120] = 25'b1111000100010100010101101;
    rom[36121] = 25'b1111000100010000011100110;
    rom[36122] = 25'b1111000100001100100100010;
    rom[36123] = 25'b1111000100001000101100001;
    rom[36124] = 25'b1111000100000100110100110;
    rom[36125] = 25'b1111000100000000111101110;
    rom[36126] = 25'b1111000011111101000111010;
    rom[36127] = 25'b1111000011111001010001010;
    rom[36128] = 25'b1111000011110101011011110;
    rom[36129] = 25'b1111000011110001100110110;
    rom[36130] = 25'b1111000011101101110010010;
    rom[36131] = 25'b1111000011101001111110010;
    rom[36132] = 25'b1111000011100110001010111;
    rom[36133] = 25'b1111000011100010010111111;
    rom[36134] = 25'b1111000011011110100101011;
    rom[36135] = 25'b1111000011011010110011011;
    rom[36136] = 25'b1111000011010111000001111;
    rom[36137] = 25'b1111000011010011010000111;
    rom[36138] = 25'b1111000011001111100000011;
    rom[36139] = 25'b1111000011001011110000100;
    rom[36140] = 25'b1111000011001000000001000;
    rom[36141] = 25'b1111000011000100010010000;
    rom[36142] = 25'b1111000011000000100011100;
    rom[36143] = 25'b1111000010111100110101100;
    rom[36144] = 25'b1111000010111001001000000;
    rom[36145] = 25'b1111000010110101011011001;
    rom[36146] = 25'b1111000010110001101110101;
    rom[36147] = 25'b1111000010101110000010101;
    rom[36148] = 25'b1111000010101010010111001;
    rom[36149] = 25'b1111000010100110101100010;
    rom[36150] = 25'b1111000010100011000001110;
    rom[36151] = 25'b1111000010011111010111101;
    rom[36152] = 25'b1111000010011011101110010;
    rom[36153] = 25'b1111000010011000000101010;
    rom[36154] = 25'b1111000010010100011100110;
    rom[36155] = 25'b1111000010010000110100110;
    rom[36156] = 25'b1111000010001101001101010;
    rom[36157] = 25'b1111000010001001100110010;
    rom[36158] = 25'b1111000010000101111111110;
    rom[36159] = 25'b1111000010000010011001111;
    rom[36160] = 25'b1111000001111110110100010;
    rom[36161] = 25'b1111000001111011001111011;
    rom[36162] = 25'b1111000001110111101010111;
    rom[36163] = 25'b1111000001110100000110111;
    rom[36164] = 25'b1111000001110000100011011;
    rom[36165] = 25'b1111000001101101000000011;
    rom[36166] = 25'b1111000001101001011101111;
    rom[36167] = 25'b1111000001100101111011111;
    rom[36168] = 25'b1111000001100010011010011;
    rom[36169] = 25'b1111000001011110111001011;
    rom[36170] = 25'b1111000001011011011000111;
    rom[36171] = 25'b1111000001010111111000111;
    rom[36172] = 25'b1111000001010100011001011;
    rom[36173] = 25'b1111000001010000111010011;
    rom[36174] = 25'b1111000001001101011011111;
    rom[36175] = 25'b1111000001001001111101111;
    rom[36176] = 25'b1111000001000110100000011;
    rom[36177] = 25'b1111000001000011000011011;
    rom[36178] = 25'b1111000000111111100110110;
    rom[36179] = 25'b1111000000111100001010110;
    rom[36180] = 25'b1111000000111000101111010;
    rom[36181] = 25'b1111000000110101010100010;
    rom[36182] = 25'b1111000000110001111001110;
    rom[36183] = 25'b1111000000101110011111110;
    rom[36184] = 25'b1111000000101011000110001;
    rom[36185] = 25'b1111000000100111101101001;
    rom[36186] = 25'b1111000000100100010100101;
    rom[36187] = 25'b1111000000100000111100100;
    rom[36188] = 25'b1111000000011101100101000;
    rom[36189] = 25'b1111000000011010001101111;
    rom[36190] = 25'b1111000000010110110111011;
    rom[36191] = 25'b1111000000010011100001011;
    rom[36192] = 25'b1111000000010000001011110;
    rom[36193] = 25'b1111000000001100110110110;
    rom[36194] = 25'b1111000000001001100010010;
    rom[36195] = 25'b1111000000000110001110001;
    rom[36196] = 25'b1111000000000010111010100;
    rom[36197] = 25'b1110111111111111100111100;
    rom[36198] = 25'b1110111111111100010100111;
    rom[36199] = 25'b1110111111111001000010111;
    rom[36200] = 25'b1110111111110101110001010;
    rom[36201] = 25'b1110111111110010100000010;
    rom[36202] = 25'b1110111111101111001111101;
    rom[36203] = 25'b1110111111101011111111100;
    rom[36204] = 25'b1110111111101000101111111;
    rom[36205] = 25'b1110111111100101100000110;
    rom[36206] = 25'b1110111111100010010010010;
    rom[36207] = 25'b1110111111011111000100001;
    rom[36208] = 25'b1110111111011011110110100;
    rom[36209] = 25'b1110111111011000101001011;
    rom[36210] = 25'b1110111111010101011100110;
    rom[36211] = 25'b1110111111010010010000101;
    rom[36212] = 25'b1110111111001111000101000;
    rom[36213] = 25'b1110111111001011111001111;
    rom[36214] = 25'b1110111111001000101111010;
    rom[36215] = 25'b1110111111000101100101000;
    rom[36216] = 25'b1110111111000010011011011;
    rom[36217] = 25'b1110111110111111010010010;
    rom[36218] = 25'b1110111110111100001001100;
    rom[36219] = 25'b1110111110111001000001011;
    rom[36220] = 25'b1110111110110101111001110;
    rom[36221] = 25'b1110111110110010110010100;
    rom[36222] = 25'b1110111110101111101011111;
    rom[36223] = 25'b1110111110101100100101101;
    rom[36224] = 25'b1110111110101001100000000;
    rom[36225] = 25'b1110111110100110011010111;
    rom[36226] = 25'b1110111110100011010110000;
    rom[36227] = 25'b1110111110100000010001111;
    rom[36228] = 25'b1110111110011101001110010;
    rom[36229] = 25'b1110111110011010001010111;
    rom[36230] = 25'b1110111110010111001000010;
    rom[36231] = 25'b1110111110010100000110000;
    rom[36232] = 25'b1110111110010001000100010;
    rom[36233] = 25'b1110111110001110000011000;
    rom[36234] = 25'b1110111110001011000010010;
    rom[36235] = 25'b1110111110001000000010000;
    rom[36236] = 25'b1110111110000101000010001;
    rom[36237] = 25'b1110111110000010000010111;
    rom[36238] = 25'b1110111101111111000100001;
    rom[36239] = 25'b1110111101111100000101111;
    rom[36240] = 25'b1110111101111001001000000;
    rom[36241] = 25'b1110111101110110001010110;
    rom[36242] = 25'b1110111101110011001101111;
    rom[36243] = 25'b1110111101110000010001101;
    rom[36244] = 25'b1110111101101101010101110;
    rom[36245] = 25'b1110111101101010011010011;
    rom[36246] = 25'b1110111101100111011111101;
    rom[36247] = 25'b1110111101100100100101010;
    rom[36248] = 25'b1110111101100001101011011;
    rom[36249] = 25'b1110111101011110110010000;
    rom[36250] = 25'b1110111101011011111001001;
    rom[36251] = 25'b1110111101011001000000110;
    rom[36252] = 25'b1110111101010110001000111;
    rom[36253] = 25'b1110111101010011010001100;
    rom[36254] = 25'b1110111101010000011010100;
    rom[36255] = 25'b1110111101001101100100001;
    rom[36256] = 25'b1110111101001010101110010;
    rom[36257] = 25'b1110111101000111111000110;
    rom[36258] = 25'b1110111101000101000011110;
    rom[36259] = 25'b1110111101000010001111011;
    rom[36260] = 25'b1110111100111111011011011;
    rom[36261] = 25'b1110111100111100100111111;
    rom[36262] = 25'b1110111100111001110100111;
    rom[36263] = 25'b1110111100110111000010011;
    rom[36264] = 25'b1110111100110100010000011;
    rom[36265] = 25'b1110111100110001011110111;
    rom[36266] = 25'b1110111100101110101101111;
    rom[36267] = 25'b1110111100101011111101011;
    rom[36268] = 25'b1110111100101001001101010;
    rom[36269] = 25'b1110111100100110011101110;
    rom[36270] = 25'b1110111100100011101110101;
    rom[36271] = 25'b1110111100100001000000001;
    rom[36272] = 25'b1110111100011110010010000;
    rom[36273] = 25'b1110111100011011100100011;
    rom[36274] = 25'b1110111100011000110111010;
    rom[36275] = 25'b1110111100010110001010101;
    rom[36276] = 25'b1110111100010011011110101;
    rom[36277] = 25'b1110111100010000110010111;
    rom[36278] = 25'b1110111100001110000111110;
    rom[36279] = 25'b1110111100001011011101001;
    rom[36280] = 25'b1110111100001000110010111;
    rom[36281] = 25'b1110111100000110001001010;
    rom[36282] = 25'b1110111100000011100000001;
    rom[36283] = 25'b1110111100000000110111011;
    rom[36284] = 25'b1110111011111110001111001;
    rom[36285] = 25'b1110111011111011100111011;
    rom[36286] = 25'b1110111011111001000000001;
    rom[36287] = 25'b1110111011110110011001011;
    rom[36288] = 25'b1110111011110011110011001;
    rom[36289] = 25'b1110111011110001001101010;
    rom[36290] = 25'b1110111011101110101000000;
    rom[36291] = 25'b1110111011101100000011010;
    rom[36292] = 25'b1110111011101001011110111;
    rom[36293] = 25'b1110111011100110111011001;
    rom[36294] = 25'b1110111011100100010111101;
    rom[36295] = 25'b1110111011100001110100111;
    rom[36296] = 25'b1110111011011111010010100;
    rom[36297] = 25'b1110111011011100110000100;
    rom[36298] = 25'b1110111011011010001111001;
    rom[36299] = 25'b1110111011010111101110010;
    rom[36300] = 25'b1110111011010101001101111;
    rom[36301] = 25'b1110111011010010101101111;
    rom[36302] = 25'b1110111011010000001110100;
    rom[36303] = 25'b1110111011001101101111100;
    rom[36304] = 25'b1110111011001011010001000;
    rom[36305] = 25'b1110111011001000110011000;
    rom[36306] = 25'b1110111011000110010101100;
    rom[36307] = 25'b1110111011000011111000011;
    rom[36308] = 25'b1110111011000001011011111;
    rom[36309] = 25'b1110111010111110111111111;
    rom[36310] = 25'b1110111010111100100100010;
    rom[36311] = 25'b1110111010111010001001001;
    rom[36312] = 25'b1110111010110111101110101;
    rom[36313] = 25'b1110111010110101010100100;
    rom[36314] = 25'b1110111010110010111010110;
    rom[36315] = 25'b1110111010110000100001110;
    rom[36316] = 25'b1110111010101110001001000;
    rom[36317] = 25'b1110111010101011110000110;
    rom[36318] = 25'b1110111010101001011001001;
    rom[36319] = 25'b1110111010100111000001111;
    rom[36320] = 25'b1110111010100100101011001;
    rom[36321] = 25'b1110111010100010010101000;
    rom[36322] = 25'b1110111010011111111111001;
    rom[36323] = 25'b1110111010011101101001111;
    rom[36324] = 25'b1110111010011011010101001;
    rom[36325] = 25'b1110111010011001000000110;
    rom[36326] = 25'b1110111010010110101101000;
    rom[36327] = 25'b1110111010010100011001101;
    rom[36328] = 25'b1110111010010010000110101;
    rom[36329] = 25'b1110111010001111110100011;
    rom[36330] = 25'b1110111010001101100010011;
    rom[36331] = 25'b1110111010001011010001000;
    rom[36332] = 25'b1110111010001001000000000;
    rom[36333] = 25'b1110111010000110101111101;
    rom[36334] = 25'b1110111010000100011111101;
    rom[36335] = 25'b1110111010000010010000001;
    rom[36336] = 25'b1110111010000000000001001;
    rom[36337] = 25'b1110111001111101110010100;
    rom[36338] = 25'b1110111001111011100100100;
    rom[36339] = 25'b1110111001111001010110111;
    rom[36340] = 25'b1110111001110111001001111;
    rom[36341] = 25'b1110111001110100111101010;
    rom[36342] = 25'b1110111001110010110001001;
    rom[36343] = 25'b1110111001110000100101100;
    rom[36344] = 25'b1110111001101110011010011;
    rom[36345] = 25'b1110111001101100001111101;
    rom[36346] = 25'b1110111001101010000101100;
    rom[36347] = 25'b1110111001100111111011110;
    rom[36348] = 25'b1110111001100101110010011;
    rom[36349] = 25'b1110111001100011101001110;
    rom[36350] = 25'b1110111001100001100001100;
    rom[36351] = 25'b1110111001011111011001101;
    rom[36352] = 25'b1110111001011101010010010;
    rom[36353] = 25'b1110111001011011001011011;
    rom[36354] = 25'b1110111001011001000101000;
    rom[36355] = 25'b1110111001010110111111010;
    rom[36356] = 25'b1110111001010100111001110;
    rom[36357] = 25'b1110111001010010110100110;
    rom[36358] = 25'b1110111001010000110000011;
    rom[36359] = 25'b1110111001001110101100011;
    rom[36360] = 25'b1110111001001100101000111;
    rom[36361] = 25'b1110111001001010100101111;
    rom[36362] = 25'b1110111001001000100011011;
    rom[36363] = 25'b1110111001000110100001010;
    rom[36364] = 25'b1110111001000100011111101;
    rom[36365] = 25'b1110111001000010011110100;
    rom[36366] = 25'b1110111001000000011101111;
    rom[36367] = 25'b1110111000111110011101110;
    rom[36368] = 25'b1110111000111100011110001;
    rom[36369] = 25'b1110111000111010011110111;
    rom[36370] = 25'b1110111000111000100000001;
    rom[36371] = 25'b1110111000110110100001111;
    rom[36372] = 25'b1110111000110100100100001;
    rom[36373] = 25'b1110111000110010100110110;
    rom[36374] = 25'b1110111000110000101001111;
    rom[36375] = 25'b1110111000101110101101101;
    rom[36376] = 25'b1110111000101100110001110;
    rom[36377] = 25'b1110111000101010110110011;
    rom[36378] = 25'b1110111000101000111011100;
    rom[36379] = 25'b1110111000100111000001000;
    rom[36380] = 25'b1110111000100101000111000;
    rom[36381] = 25'b1110111000100011001101100;
    rom[36382] = 25'b1110111000100001010100100;
    rom[36383] = 25'b1110111000011111011100000;
    rom[36384] = 25'b1110111000011101100011111;
    rom[36385] = 25'b1110111000011011101100010;
    rom[36386] = 25'b1110111000011001110101001;
    rom[36387] = 25'b1110111000010111111110100;
    rom[36388] = 25'b1110111000010110001000011;
    rom[36389] = 25'b1110111000010100010010101;
    rom[36390] = 25'b1110111000010010011101011;
    rom[36391] = 25'b1110111000010000101000101;
    rom[36392] = 25'b1110111000001110110100010;
    rom[36393] = 25'b1110111000001101000000100;
    rom[36394] = 25'b1110111000001011001101001;
    rom[36395] = 25'b1110111000001001011010010;
    rom[36396] = 25'b1110111000000111100111111;
    rom[36397] = 25'b1110111000000101110110000;
    rom[36398] = 25'b1110111000000100000100100;
    rom[36399] = 25'b1110111000000010010011101;
    rom[36400] = 25'b1110111000000000100011000;
    rom[36401] = 25'b1110110111111110110011000;
    rom[36402] = 25'b1110110111111101000011100;
    rom[36403] = 25'b1110110111111011010100011;
    rom[36404] = 25'b1110110111111001100101101;
    rom[36405] = 25'b1110110111110111110111101;
    rom[36406] = 25'b1110110111110110001001111;
    rom[36407] = 25'b1110110111110100011100101;
    rom[36408] = 25'b1110110111110010110000000;
    rom[36409] = 25'b1110110111110001000011101;
    rom[36410] = 25'b1110110111101111010111111;
    rom[36411] = 25'b1110110111101101101100101;
    rom[36412] = 25'b1110110111101100000001101;
    rom[36413] = 25'b1110110111101010010111010;
    rom[36414] = 25'b1110110111101000101101011;
    rom[36415] = 25'b1110110111100111000100000;
    rom[36416] = 25'b1110110111100101011010111;
    rom[36417] = 25'b1110110111100011110010011;
    rom[36418] = 25'b1110110111100010001010011;
    rom[36419] = 25'b1110110111100000100010110;
    rom[36420] = 25'b1110110111011110111011110;
    rom[36421] = 25'b1110110111011101010101000;
    rom[36422] = 25'b1110110111011011101110111;
    rom[36423] = 25'b1110110111011010001001010;
    rom[36424] = 25'b1110110111011000100100000;
    rom[36425] = 25'b1110110111010110111111010;
    rom[36426] = 25'b1110110111010101011010111;
    rom[36427] = 25'b1110110111010011110111000;
    rom[36428] = 25'b1110110111010010010011101;
    rom[36429] = 25'b1110110111010000110000110;
    rom[36430] = 25'b1110110111001111001110010;
    rom[36431] = 25'b1110110111001101101100011;
    rom[36432] = 25'b1110110111001100001010111;
    rom[36433] = 25'b1110110111001010101001110;
    rom[36434] = 25'b1110110111001001001001010;
    rom[36435] = 25'b1110110111000111101001001;
    rom[36436] = 25'b1110110111000110001001100;
    rom[36437] = 25'b1110110111000100101010011;
    rom[36438] = 25'b1110110111000011001011101;
    rom[36439] = 25'b1110110111000001101101011;
    rom[36440] = 25'b1110110111000000001111101;
    rom[36441] = 25'b1110110110111110110010010;
    rom[36442] = 25'b1110110110111101010101100;
    rom[36443] = 25'b1110110110111011111001000;
    rom[36444] = 25'b1110110110111010011101001;
    rom[36445] = 25'b1110110110111001000001101;
    rom[36446] = 25'b1110110110110111100110101;
    rom[36447] = 25'b1110110110110110001100001;
    rom[36448] = 25'b1110110110110100110010001;
    rom[36449] = 25'b1110110110110011011000100;
    rom[36450] = 25'b1110110110110001111111011;
    rom[36451] = 25'b1110110110110000100110101;
    rom[36452] = 25'b1110110110101111001110011;
    rom[36453] = 25'b1110110110101101110110110;
    rom[36454] = 25'b1110110110101100011111011;
    rom[36455] = 25'b1110110110101011001000100;
    rom[36456] = 25'b1110110110101001110010001;
    rom[36457] = 25'b1110110110101000011100010;
    rom[36458] = 25'b1110110110100111000110111;
    rom[36459] = 25'b1110110110100101110001111;
    rom[36460] = 25'b1110110110100100011101010;
    rom[36461] = 25'b1110110110100011001001010;
    rom[36462] = 25'b1110110110100001110101101;
    rom[36463] = 25'b1110110110100000100010100;
    rom[36464] = 25'b1110110110011111001111111;
    rom[36465] = 25'b1110110110011101111101101;
    rom[36466] = 25'b1110110110011100101011111;
    rom[36467] = 25'b1110110110011011011010101;
    rom[36468] = 25'b1110110110011010001001110;
    rom[36469] = 25'b1110110110011000111001011;
    rom[36470] = 25'b1110110110010111101001100;
    rom[36471] = 25'b1110110110010110011010000;
    rom[36472] = 25'b1110110110010101001011000;
    rom[36473] = 25'b1110110110010011111100100;
    rom[36474] = 25'b1110110110010010101110011;
    rom[36475] = 25'b1110110110010001100000110;
    rom[36476] = 25'b1110110110010000010011100;
    rom[36477] = 25'b1110110110001111000110111;
    rom[36478] = 25'b1110110110001101111010101;
    rom[36479] = 25'b1110110110001100101110111;
    rom[36480] = 25'b1110110110001011100011100;
    rom[36481] = 25'b1110110110001010011000101;
    rom[36482] = 25'b1110110110001001001110001;
    rom[36483] = 25'b1110110110001000000100001;
    rom[36484] = 25'b1110110110000110111010101;
    rom[36485] = 25'b1110110110000101110001101;
    rom[36486] = 25'b1110110110000100101001000;
    rom[36487] = 25'b1110110110000011100000111;
    rom[36488] = 25'b1110110110000010011001001;
    rom[36489] = 25'b1110110110000001010001111;
    rom[36490] = 25'b1110110110000000001011001;
    rom[36491] = 25'b1110110101111111000100111;
    rom[36492] = 25'b1110110101111101111111000;
    rom[36493] = 25'b1110110101111100111001101;
    rom[36494] = 25'b1110110101111011110100101;
    rom[36495] = 25'b1110110101111010110000001;
    rom[36496] = 25'b1110110101111001101100000;
    rom[36497] = 25'b1110110101111000101000011;
    rom[36498] = 25'b1110110101110111100101010;
    rom[36499] = 25'b1110110101110110100010101;
    rom[36500] = 25'b1110110101110101100000011;
    rom[36501] = 25'b1110110101110100011110101;
    rom[36502] = 25'b1110110101110011011101010;
    rom[36503] = 25'b1110110101110010011100011;
    rom[36504] = 25'b1110110101110001011011111;
    rom[36505] = 25'b1110110101110000011100000;
    rom[36506] = 25'b1110110101101111011100100;
    rom[36507] = 25'b1110110101101110011101011;
    rom[36508] = 25'b1110110101101101011110110;
    rom[36509] = 25'b1110110101101100100000101;
    rom[36510] = 25'b1110110101101011100010111;
    rom[36511] = 25'b1110110101101010100101101;
    rom[36512] = 25'b1110110101101001101000111;
    rom[36513] = 25'b1110110101101000101100100;
    rom[36514] = 25'b1110110101100111110000101;
    rom[36515] = 25'b1110110101100110110101001;
    rom[36516] = 25'b1110110101100101111010001;
    rom[36517] = 25'b1110110101100100111111100;
    rom[36518] = 25'b1110110101100100000101100;
    rom[36519] = 25'b1110110101100011001011110;
    rom[36520] = 25'b1110110101100010010010101;
    rom[36521] = 25'b1110110101100001011001110;
    rom[36522] = 25'b1110110101100000100001100;
    rom[36523] = 25'b1110110101011111101001100;
    rom[36524] = 25'b1110110101011110110010001;
    rom[36525] = 25'b1110110101011101111011001;
    rom[36526] = 25'b1110110101011101000100101;
    rom[36527] = 25'b1110110101011100001110100;
    rom[36528] = 25'b1110110101011011011001000;
    rom[36529] = 25'b1110110101011010100011110;
    rom[36530] = 25'b1110110101011001101111000;
    rom[36531] = 25'b1110110101011000111010110;
    rom[36532] = 25'b1110110101011000000110111;
    rom[36533] = 25'b1110110101010111010011100;
    rom[36534] = 25'b1110110101010110100000101;
    rom[36535] = 25'b1110110101010101101110000;
    rom[36536] = 25'b1110110101010100111100000;
    rom[36537] = 25'b1110110101010100001010011;
    rom[36538] = 25'b1110110101010011011001001;
    rom[36539] = 25'b1110110101010010101000100;
    rom[36540] = 25'b1110110101010001111000010;
    rom[36541] = 25'b1110110101010001001000011;
    rom[36542] = 25'b1110110101010000011001000;
    rom[36543] = 25'b1110110101001111101010000;
    rom[36544] = 25'b1110110101001110111011100;
    rom[36545] = 25'b1110110101001110001101100;
    rom[36546] = 25'b1110110101001101011111111;
    rom[36547] = 25'b1110110101001100110010110;
    rom[36548] = 25'b1110110101001100000110000;
    rom[36549] = 25'b1110110101001011011001110;
    rom[36550] = 25'b1110110101001010101101111;
    rom[36551] = 25'b1110110101001010000010100;
    rom[36552] = 25'b1110110101001001010111100;
    rom[36553] = 25'b1110110101001000101101000;
    rom[36554] = 25'b1110110101001000000010111;
    rom[36555] = 25'b1110110101000111011001010;
    rom[36556] = 25'b1110110101000110110000001;
    rom[36557] = 25'b1110110101000110000111011;
    rom[36558] = 25'b1110110101000101011111000;
    rom[36559] = 25'b1110110101000100110111001;
    rom[36560] = 25'b1110110101000100001111110;
    rom[36561] = 25'b1110110101000011101000110;
    rom[36562] = 25'b1110110101000011000010010;
    rom[36563] = 25'b1110110101000010011100001;
    rom[36564] = 25'b1110110101000001110110011;
    rom[36565] = 25'b1110110101000001010001010;
    rom[36566] = 25'b1110110101000000101100011;
    rom[36567] = 25'b1110110101000000001000001;
    rom[36568] = 25'b1110110100111111100100001;
    rom[36569] = 25'b1110110100111111000000101;
    rom[36570] = 25'b1110110100111110011101101;
    rom[36571] = 25'b1110110100111101111011001;
    rom[36572] = 25'b1110110100111101011000111;
    rom[36573] = 25'b1110110100111100110111010;
    rom[36574] = 25'b1110110100111100010101111;
    rom[36575] = 25'b1110110100111011110101000;
    rom[36576] = 25'b1110110100111011010100101;
    rom[36577] = 25'b1110110100111010110100101;
    rom[36578] = 25'b1110110100111010010101001;
    rom[36579] = 25'b1110110100111001110110000;
    rom[36580] = 25'b1110110100111001010111011;
    rom[36581] = 25'b1110110100111000111001001;
    rom[36582] = 25'b1110110100111000011011010;
    rom[36583] = 25'b1110110100110111111110000;
    rom[36584] = 25'b1110110100110111100001000;
    rom[36585] = 25'b1110110100110111000100100;
    rom[36586] = 25'b1110110100110110101000011;
    rom[36587] = 25'b1110110100110110001100110;
    rom[36588] = 25'b1110110100110101110001101;
    rom[36589] = 25'b1110110100110101010110111;
    rom[36590] = 25'b1110110100110100111100101;
    rom[36591] = 25'b1110110100110100100010110;
    rom[36592] = 25'b1110110100110100001001010;
    rom[36593] = 25'b1110110100110011110000001;
    rom[36594] = 25'b1110110100110011010111101;
    rom[36595] = 25'b1110110100110010111111011;
    rom[36596] = 25'b1110110100110010100111110;
    rom[36597] = 25'b1110110100110010010000100;
    rom[36598] = 25'b1110110100110001111001101;
    rom[36599] = 25'b1110110100110001100011001;
    rom[36600] = 25'b1110110100110001001101001;
    rom[36601] = 25'b1110110100110000110111100;
    rom[36602] = 25'b1110110100110000100010100;
    rom[36603] = 25'b1110110100110000001101110;
    rom[36604] = 25'b1110110100101111111001100;
    rom[36605] = 25'b1110110100101111100101100;
    rom[36606] = 25'b1110110100101111010010001;
    rom[36607] = 25'b1110110100101110111111001;
    rom[36608] = 25'b1110110100101110101100101;
    rom[36609] = 25'b1110110100101110011010100;
    rom[36610] = 25'b1110110100101110001000110;
    rom[36611] = 25'b1110110100101101110111100;
    rom[36612] = 25'b1110110100101101100110101;
    rom[36613] = 25'b1110110100101101010110010;
    rom[36614] = 25'b1110110100101101000110010;
    rom[36615] = 25'b1110110100101100110110101;
    rom[36616] = 25'b1110110100101100100111100;
    rom[36617] = 25'b1110110100101100011000110;
    rom[36618] = 25'b1110110100101100001010101;
    rom[36619] = 25'b1110110100101011111100101;
    rom[36620] = 25'b1110110100101011101111010;
    rom[36621] = 25'b1110110100101011100010010;
    rom[36622] = 25'b1110110100101011010101101;
    rom[36623] = 25'b1110110100101011001001100;
    rom[36624] = 25'b1110110100101010111101110;
    rom[36625] = 25'b1110110100101010110010100;
    rom[36626] = 25'b1110110100101010100111101;
    rom[36627] = 25'b1110110100101010011101001;
    rom[36628] = 25'b1110110100101010010011001;
    rom[36629] = 25'b1110110100101010001001100;
    rom[36630] = 25'b1110110100101010000000011;
    rom[36631] = 25'b1110110100101001110111101;
    rom[36632] = 25'b1110110100101001101111001;
    rom[36633] = 25'b1110110100101001100111011;
    rom[36634] = 25'b1110110100101001011111111;
    rom[36635] = 25'b1110110100101001011000110;
    rom[36636] = 25'b1110110100101001010010001;
    rom[36637] = 25'b1110110100101001001011111;
    rom[36638] = 25'b1110110100101001000110001;
    rom[36639] = 25'b1110110100101001000000101;
    rom[36640] = 25'b1110110100101000111011110;
    rom[36641] = 25'b1110110100101000110111010;
    rom[36642] = 25'b1110110100101000110011001;
    rom[36643] = 25'b1110110100101000101111011;
    rom[36644] = 25'b1110110100101000101100001;
    rom[36645] = 25'b1110110100101000101001010;
    rom[36646] = 25'b1110110100101000100110110;
    rom[36647] = 25'b1110110100101000100100111;
    rom[36648] = 25'b1110110100101000100011001;
    rom[36649] = 25'b1110110100101000100010000;
    rom[36650] = 25'b1110110100101000100001010;
    rom[36651] = 25'b1110110100101000100000111;
    rom[36652] = 25'b1110110100101000100001000;
    rom[36653] = 25'b1110110100101000100001100;
    rom[36654] = 25'b1110110100101000100010011;
    rom[36655] = 25'b1110110100101000100011110;
    rom[36656] = 25'b1110110100101000100101100;
    rom[36657] = 25'b1110110100101000100111101;
    rom[36658] = 25'b1110110100101000101010010;
    rom[36659] = 25'b1110110100101000101101010;
    rom[36660] = 25'b1110110100101000110000101;
    rom[36661] = 25'b1110110100101000110100011;
    rom[36662] = 25'b1110110100101000111000110;
    rom[36663] = 25'b1110110100101000111101010;
    rom[36664] = 25'b1110110100101001000010100;
    rom[36665] = 25'b1110110100101001001000000;
    rom[36666] = 25'b1110110100101001001101111;
    rom[36667] = 25'b1110110100101001010100001;
    rom[36668] = 25'b1110110100101001011010111;
    rom[36669] = 25'b1110110100101001100010000;
    rom[36670] = 25'b1110110100101001101001101;
    rom[36671] = 25'b1110110100101001110001100;
    rom[36672] = 25'b1110110100101001111001111;
    rom[36673] = 25'b1110110100101010000010110;
    rom[36674] = 25'b1110110100101010001011111;
    rom[36675] = 25'b1110110100101010010101100;
    rom[36676] = 25'b1110110100101010011111100;
    rom[36677] = 25'b1110110100101010101010000;
    rom[36678] = 25'b1110110100101010110100111;
    rom[36679] = 25'b1110110100101011000000001;
    rom[36680] = 25'b1110110100101011001011110;
    rom[36681] = 25'b1110110100101011011000000;
    rom[36682] = 25'b1110110100101011100100100;
    rom[36683] = 25'b1110110100101011110001011;
    rom[36684] = 25'b1110110100101011111110101;
    rom[36685] = 25'b1110110100101100001100011;
    rom[36686] = 25'b1110110100101100011010100;
    rom[36687] = 25'b1110110100101100101001001;
    rom[36688] = 25'b1110110100101100111000000;
    rom[36689] = 25'b1110110100101101000111011;
    rom[36690] = 25'b1110110100101101010111001;
    rom[36691] = 25'b1110110100101101100111010;
    rom[36692] = 25'b1110110100101101110111111;
    rom[36693] = 25'b1110110100101110001000111;
    rom[36694] = 25'b1110110100101110011010010;
    rom[36695] = 25'b1110110100101110101100001;
    rom[36696] = 25'b1110110100101110111110011;
    rom[36697] = 25'b1110110100101111010001000;
    rom[36698] = 25'b1110110100101111100100000;
    rom[36699] = 25'b1110110100101111110111100;
    rom[36700] = 25'b1110110100110000001011010;
    rom[36701] = 25'b1110110100110000011111100;
    rom[36702] = 25'b1110110100110000110100010;
    rom[36703] = 25'b1110110100110001001001010;
    rom[36704] = 25'b1110110100110001011110101;
    rom[36705] = 25'b1110110100110001110100100;
    rom[36706] = 25'b1110110100110010001010111;
    rom[36707] = 25'b1110110100110010100001100;
    rom[36708] = 25'b1110110100110010111000101;
    rom[36709] = 25'b1110110100110011010000000;
    rom[36710] = 25'b1110110100110011101000000;
    rom[36711] = 25'b1110110100110100000000010;
    rom[36712] = 25'b1110110100110100011000111;
    rom[36713] = 25'b1110110100110100110010000;
    rom[36714] = 25'b1110110100110101001011100;
    rom[36715] = 25'b1110110100110101100101011;
    rom[36716] = 25'b1110110100110101111111101;
    rom[36717] = 25'b1110110100110110011010011;
    rom[36718] = 25'b1110110100110110110101011;
    rom[36719] = 25'b1110110100110111010001000;
    rom[36720] = 25'b1110110100110111101100110;
    rom[36721] = 25'b1110110100111000001001001;
    rom[36722] = 25'b1110110100111000100101111;
    rom[36723] = 25'b1110110100111001000010111;
    rom[36724] = 25'b1110110100111001100000011;
    rom[36725] = 25'b1110110100111001111110010;
    rom[36726] = 25'b1110110100111010011100100;
    rom[36727] = 25'b1110110100111010111011010;
    rom[36728] = 25'b1110110100111011011010011;
    rom[36729] = 25'b1110110100111011111001111;
    rom[36730] = 25'b1110110100111100011001101;
    rom[36731] = 25'b1110110100111100111010000;
    rom[36732] = 25'b1110110100111101011010101;
    rom[36733] = 25'b1110110100111101111011110;
    rom[36734] = 25'b1110110100111110011101001;
    rom[36735] = 25'b1110110100111110111111001;
    rom[36736] = 25'b1110110100111111100001010;
    rom[36737] = 25'b1110110101000000000011111;
    rom[36738] = 25'b1110110101000000100111000;
    rom[36739] = 25'b1110110101000001001010011;
    rom[36740] = 25'b1110110101000001101110010;
    rom[36741] = 25'b1110110101000010010010100;
    rom[36742] = 25'b1110110101000010110111001;
    rom[36743] = 25'b1110110101000011011100001;
    rom[36744] = 25'b1110110101000100000001100;
    rom[36745] = 25'b1110110101000100100111011;
    rom[36746] = 25'b1110110101000101001101100;
    rom[36747] = 25'b1110110101000101110100001;
    rom[36748] = 25'b1110110101000110011011001;
    rom[36749] = 25'b1110110101000111000010100;
    rom[36750] = 25'b1110110101000111101010010;
    rom[36751] = 25'b1110110101001000010010011;
    rom[36752] = 25'b1110110101001000111011000;
    rom[36753] = 25'b1110110101001001100011111;
    rom[36754] = 25'b1110110101001010001101010;
    rom[36755] = 25'b1110110101001010110110111;
    rom[36756] = 25'b1110110101001011100001000;
    rom[36757] = 25'b1110110101001100001011100;
    rom[36758] = 25'b1110110101001100110110011;
    rom[36759] = 25'b1110110101001101100001101;
    rom[36760] = 25'b1110110101001110001101011;
    rom[36761] = 25'b1110110101001110111001011;
    rom[36762] = 25'b1110110101001111100101111;
    rom[36763] = 25'b1110110101010000010010101;
    rom[36764] = 25'b1110110101010000111111111;
    rom[36765] = 25'b1110110101010001101101100;
    rom[36766] = 25'b1110110101010010011011100;
    rom[36767] = 25'b1110110101010011001001111;
    rom[36768] = 25'b1110110101010011111000100;
    rom[36769] = 25'b1110110101010100100111110;
    rom[36770] = 25'b1110110101010101010111010;
    rom[36771] = 25'b1110110101010110000111001;
    rom[36772] = 25'b1110110101010110110111100;
    rom[36773] = 25'b1110110101010111101000010;
    rom[36774] = 25'b1110110101011000011001010;
    rom[36775] = 25'b1110110101011001001010110;
    rom[36776] = 25'b1110110101011001111100101;
    rom[36777] = 25'b1110110101011010101110111;
    rom[36778] = 25'b1110110101011011100001100;
    rom[36779] = 25'b1110110101011100010100011;
    rom[36780] = 25'b1110110101011101000111110;
    rom[36781] = 25'b1110110101011101111011100;
    rom[36782] = 25'b1110110101011110101111101;
    rom[36783] = 25'b1110110101011111100100010;
    rom[36784] = 25'b1110110101100000011001001;
    rom[36785] = 25'b1110110101100001001110011;
    rom[36786] = 25'b1110110101100010000100000;
    rom[36787] = 25'b1110110101100010111010001;
    rom[36788] = 25'b1110110101100011110000100;
    rom[36789] = 25'b1110110101100100100111011;
    rom[36790] = 25'b1110110101100101011110100;
    rom[36791] = 25'b1110110101100110010110001;
    rom[36792] = 25'b1110110101100111001110000;
    rom[36793] = 25'b1110110101101000000110011;
    rom[36794] = 25'b1110110101101000111111000;
    rom[36795] = 25'b1110110101101001111000001;
    rom[36796] = 25'b1110110101101010110001101;
    rom[36797] = 25'b1110110101101011101011011;
    rom[36798] = 25'b1110110101101100100101110;
    rom[36799] = 25'b1110110101101101100000010;
    rom[36800] = 25'b1110110101101110011011001;
    rom[36801] = 25'b1110110101101111010110101;
    rom[36802] = 25'b1110110101110000010010010;
    rom[36803] = 25'b1110110101110001001110011;
    rom[36804] = 25'b1110110101110010001010111;
    rom[36805] = 25'b1110110101110011000111110;
    rom[36806] = 25'b1110110101110100000101000;
    rom[36807] = 25'b1110110101110101000010100;
    rom[36808] = 25'b1110110101110110000000100;
    rom[36809] = 25'b1110110101110110111110111;
    rom[36810] = 25'b1110110101110111111101100;
    rom[36811] = 25'b1110110101111000111100101;
    rom[36812] = 25'b1110110101111001111100010;
    rom[36813] = 25'b1110110101111010111100000;
    rom[36814] = 25'b1110110101111011111100010;
    rom[36815] = 25'b1110110101111100111100111;
    rom[36816] = 25'b1110110101111101111101110;
    rom[36817] = 25'b1110110101111110111111001;
    rom[36818] = 25'b1110110110000000000000110;
    rom[36819] = 25'b1110110110000001000010111;
    rom[36820] = 25'b1110110110000010000101010;
    rom[36821] = 25'b1110110110000011001000001;
    rom[36822] = 25'b1110110110000100001011010;
    rom[36823] = 25'b1110110110000101001110111;
    rom[36824] = 25'b1110110110000110010010110;
    rom[36825] = 25'b1110110110000111010111001;
    rom[36826] = 25'b1110110110001000011011110;
    rom[36827] = 25'b1110110110001001100000111;
    rom[36828] = 25'b1110110110001010100110010;
    rom[36829] = 25'b1110110110001011101100000;
    rom[36830] = 25'b1110110110001100110010001;
    rom[36831] = 25'b1110110110001101111000101;
    rom[36832] = 25'b1110110110001110111111100;
    rom[36833] = 25'b1110110110010000000110110;
    rom[36834] = 25'b1110110110010001001110011;
    rom[36835] = 25'b1110110110010010010110010;
    rom[36836] = 25'b1110110110010011011110101;
    rom[36837] = 25'b1110110110010100100111011;
    rom[36838] = 25'b1110110110010101110000011;
    rom[36839] = 25'b1110110110010110111001111;
    rom[36840] = 25'b1110110110011000000011110;
    rom[36841] = 25'b1110110110011001001101111;
    rom[36842] = 25'b1110110110011010011000011;
    rom[36843] = 25'b1110110110011011100011010;
    rom[36844] = 25'b1110110110011100101110100;
    rom[36845] = 25'b1110110110011101111010001;
    rom[36846] = 25'b1110110110011111000110001;
    rom[36847] = 25'b1110110110100000010010011;
    rom[36848] = 25'b1110110110100001011111001;
    rom[36849] = 25'b1110110110100010101100010;
    rom[36850] = 25'b1110110110100011111001101;
    rom[36851] = 25'b1110110110100101000111011;
    rom[36852] = 25'b1110110110100110010101101;
    rom[36853] = 25'b1110110110100111100100001;
    rom[36854] = 25'b1110110110101000110011000;
    rom[36855] = 25'b1110110110101010000010010;
    rom[36856] = 25'b1110110110101011010001110;
    rom[36857] = 25'b1110110110101100100001110;
    rom[36858] = 25'b1110110110101101110010000;
    rom[36859] = 25'b1110110110101111000010110;
    rom[36860] = 25'b1110110110110000010011110;
    rom[36861] = 25'b1110110110110001100101001;
    rom[36862] = 25'b1110110110110010110110111;
    rom[36863] = 25'b1110110110110100001001000;
    rom[36864] = 25'b1110110110110101011011100;
    rom[36865] = 25'b1110110110110110101110010;
    rom[36866] = 25'b1110110110111000000001011;
    rom[36867] = 25'b1110110110111001010100111;
    rom[36868] = 25'b1110110110111010101000111;
    rom[36869] = 25'b1110110110111011111101001;
    rom[36870] = 25'b1110110110111101010001110;
    rom[36871] = 25'b1110110110111110100110101;
    rom[36872] = 25'b1110110110111111111100000;
    rom[36873] = 25'b1110110111000001010001101;
    rom[36874] = 25'b1110110111000010100111101;
    rom[36875] = 25'b1110110111000011111110000;
    rom[36876] = 25'b1110110111000101010100110;
    rom[36877] = 25'b1110110111000110101011110;
    rom[36878] = 25'b1110110111001000000011010;
    rom[36879] = 25'b1110110111001001011011000;
    rom[36880] = 25'b1110110111001010110011001;
    rom[36881] = 25'b1110110111001100001011101;
    rom[36882] = 25'b1110110111001101100100100;
    rom[36883] = 25'b1110110111001110111101101;
    rom[36884] = 25'b1110110111010000010111001;
    rom[36885] = 25'b1110110111010001110001000;
    rom[36886] = 25'b1110110111010011001011010;
    rom[36887] = 25'b1110110111010100100101111;
    rom[36888] = 25'b1110110111010110000000111;
    rom[36889] = 25'b1110110111010111011100001;
    rom[36890] = 25'b1110110111011000110111110;
    rom[36891] = 25'b1110110111011010010011110;
    rom[36892] = 25'b1110110111011011110000001;
    rom[36893] = 25'b1110110111011101001100110;
    rom[36894] = 25'b1110110111011110101001110;
    rom[36895] = 25'b1110110111100000000111001;
    rom[36896] = 25'b1110110111100001100100111;
    rom[36897] = 25'b1110110111100011000011000;
    rom[36898] = 25'b1110110111100100100001011;
    rom[36899] = 25'b1110110111100110000000001;
    rom[36900] = 25'b1110110111100111011111010;
    rom[36901] = 25'b1110110111101000111110101;
    rom[36902] = 25'b1110110111101010011110100;
    rom[36903] = 25'b1110110111101011111110101;
    rom[36904] = 25'b1110110111101101011111001;
    rom[36905] = 25'b1110110111101111000000000;
    rom[36906] = 25'b1110110111110000100001001;
    rom[36907] = 25'b1110110111110010000010101;
    rom[36908] = 25'b1110110111110011100100100;
    rom[36909] = 25'b1110110111110101000110110;
    rom[36910] = 25'b1110110111110110101001010;
    rom[36911] = 25'b1110110111111000001100001;
    rom[36912] = 25'b1110110111111001101111011;
    rom[36913] = 25'b1110110111111011010011000;
    rom[36914] = 25'b1110110111111100110110111;
    rom[36915] = 25'b1110110111111110011011001;
    rom[36916] = 25'b1110110111111111111111110;
    rom[36917] = 25'b1110111000000001100100101;
    rom[36918] = 25'b1110111000000011001001111;
    rom[36919] = 25'b1110111000000100101111100;
    rom[36920] = 25'b1110111000000110010101100;
    rom[36921] = 25'b1110111000000111111011110;
    rom[36922] = 25'b1110111000001001100010011;
    rom[36923] = 25'b1110111000001011001001011;
    rom[36924] = 25'b1110111000001100110000110;
    rom[36925] = 25'b1110111000001110011000011;
    rom[36926] = 25'b1110111000010000000000010;
    rom[36927] = 25'b1110111000010001101000101;
    rom[36928] = 25'b1110111000010011010001010;
    rom[36929] = 25'b1110111000010100111010010;
    rom[36930] = 25'b1110111000010110100011101;
    rom[36931] = 25'b1110111000011000001101011;
    rom[36932] = 25'b1110111000011001110111011;
    rom[36933] = 25'b1110111000011011100001101;
    rom[36934] = 25'b1110111000011101001100011;
    rom[36935] = 25'b1110111000011110110111010;
    rom[36936] = 25'b1110111000100000100010101;
    rom[36937] = 25'b1110111000100010001110011;
    rom[36938] = 25'b1110111000100011111010010;
    rom[36939] = 25'b1110111000100101100110101;
    rom[36940] = 25'b1110111000100111010011011;
    rom[36941] = 25'b1110111000101001000000010;
    rom[36942] = 25'b1110111000101010101101101;
    rom[36943] = 25'b1110111000101100011011010;
    rom[36944] = 25'b1110111000101110001001010;
    rom[36945] = 25'b1110111000101111110111101;
    rom[36946] = 25'b1110111000110001100110011;
    rom[36947] = 25'b1110111000110011010101010;
    rom[36948] = 25'b1110111000110101000100101;
    rom[36949] = 25'b1110111000110110110100010;
    rom[36950] = 25'b1110111000111000100100010;
    rom[36951] = 25'b1110111000111010010100100;
    rom[36952] = 25'b1110111000111100000101001;
    rom[36953] = 25'b1110111000111101110110001;
    rom[36954] = 25'b1110111000111111100111011;
    rom[36955] = 25'b1110111001000001011001001;
    rom[36956] = 25'b1110111001000011001011000;
    rom[36957] = 25'b1110111001000100111101010;
    rom[36958] = 25'b1110111001000110101111111;
    rom[36959] = 25'b1110111001001000100010111;
    rom[36960] = 25'b1110111001001010010110001;
    rom[36961] = 25'b1110111001001100001001101;
    rom[36962] = 25'b1110111001001101111101100;
    rom[36963] = 25'b1110111001001111110001110;
    rom[36964] = 25'b1110111001010001100110011;
    rom[36965] = 25'b1110111001010011011011010;
    rom[36966] = 25'b1110111001010101010000100;
    rom[36967] = 25'b1110111001010111000101111;
    rom[36968] = 25'b1110111001011000111011110;
    rom[36969] = 25'b1110111001011010110001111;
    rom[36970] = 25'b1110111001011100101000011;
    rom[36971] = 25'b1110111001011110011111010;
    rom[36972] = 25'b1110111001100000010110011;
    rom[36973] = 25'b1110111001100010001101111;
    rom[36974] = 25'b1110111001100100000101101;
    rom[36975] = 25'b1110111001100101111101110;
    rom[36976] = 25'b1110111001100111110110010;
    rom[36977] = 25'b1110111001101001101111000;
    rom[36978] = 25'b1110111001101011101000000;
    rom[36979] = 25'b1110111001101101100001011;
    rom[36980] = 25'b1110111001101111011011000;
    rom[36981] = 25'b1110111001110001010101000;
    rom[36982] = 25'b1110111001110011001111011;
    rom[36983] = 25'b1110111001110101001010001;
    rom[36984] = 25'b1110111001110111000101000;
    rom[36985] = 25'b1110111001111001000000011;
    rom[36986] = 25'b1110111001111010111100000;
    rom[36987] = 25'b1110111001111100110111111;
    rom[36988] = 25'b1110111001111110110100001;
    rom[36989] = 25'b1110111010000000110000101;
    rom[36990] = 25'b1110111010000010101101100;
    rom[36991] = 25'b1110111010000100101010101;
    rom[36992] = 25'b1110111010000110101000010;
    rom[36993] = 25'b1110111010001000100110001;
    rom[36994] = 25'b1110111010001010100100001;
    rom[36995] = 25'b1110111010001100100010101;
    rom[36996] = 25'b1110111010001110100001011;
    rom[36997] = 25'b1110111010010000100000011;
    rom[36998] = 25'b1110111010010010011111111;
    rom[36999] = 25'b1110111010010100011111100;
    rom[37000] = 25'b1110111010010110011111101;
    rom[37001] = 25'b1110111010011000011111111;
    rom[37002] = 25'b1110111010011010100000100;
    rom[37003] = 25'b1110111010011100100001100;
    rom[37004] = 25'b1110111010011110100010110;
    rom[37005] = 25'b1110111010100000100100011;
    rom[37006] = 25'b1110111010100010100110001;
    rom[37007] = 25'b1110111010100100101000011;
    rom[37008] = 25'b1110111010100110101010111;
    rom[37009] = 25'b1110111010101000101101110;
    rom[37010] = 25'b1110111010101010110000111;
    rom[37011] = 25'b1110111010101100110100010;
    rom[37012] = 25'b1110111010101110111000000;
    rom[37013] = 25'b1110111010110000111100000;
    rom[37014] = 25'b1110111010110011000000011;
    rom[37015] = 25'b1110111010110101000101000;
    rom[37016] = 25'b1110111010110111001010000;
    rom[37017] = 25'b1110111010111001001111010;
    rom[37018] = 25'b1110111010111011010100111;
    rom[37019] = 25'b1110111010111101011010110;
    rom[37020] = 25'b1110111010111111100000111;
    rom[37021] = 25'b1110111011000001100111011;
    rom[37022] = 25'b1110111011000011101110010;
    rom[37023] = 25'b1110111011000101110101010;
    rom[37024] = 25'b1110111011000111111100101;
    rom[37025] = 25'b1110111011001010000100100;
    rom[37026] = 25'b1110111011001100001100011;
    rom[37027] = 25'b1110111011001110010100110;
    rom[37028] = 25'b1110111011010000011101011;
    rom[37029] = 25'b1110111011010010100110010;
    rom[37030] = 25'b1110111011010100101111100;
    rom[37031] = 25'b1110111011010110111001000;
    rom[37032] = 25'b1110111011011001000010111;
    rom[37033] = 25'b1110111011011011001101000;
    rom[37034] = 25'b1110111011011101010111011;
    rom[37035] = 25'b1110111011011111100010001;
    rom[37036] = 25'b1110111011100001101101001;
    rom[37037] = 25'b1110111011100011111000100;
    rom[37038] = 25'b1110111011100110000100001;
    rom[37039] = 25'b1110111011101000010000001;
    rom[37040] = 25'b1110111011101010011100010;
    rom[37041] = 25'b1110111011101100101000110;
    rom[37042] = 25'b1110111011101110110101101;
    rom[37043] = 25'b1110111011110001000010110;
    rom[37044] = 25'b1110111011110011010000001;
    rom[37045] = 25'b1110111011110101011101111;
    rom[37046] = 25'b1110111011110111101011111;
    rom[37047] = 25'b1110111011111001111010001;
    rom[37048] = 25'b1110111011111100001000110;
    rom[37049] = 25'b1110111011111110010111101;
    rom[37050] = 25'b1110111100000000100110111;
    rom[37051] = 25'b1110111100000010110110011;
    rom[37052] = 25'b1110111100000101000110001;
    rom[37053] = 25'b1110111100000111010110001;
    rom[37054] = 25'b1110111100001001100110100;
    rom[37055] = 25'b1110111100001011110111001;
    rom[37056] = 25'b1110111100001110001000001;
    rom[37057] = 25'b1110111100010000011001011;
    rom[37058] = 25'b1110111100010010101010111;
    rom[37059] = 25'b1110111100010100111100110;
    rom[37060] = 25'b1110111100010111001110111;
    rom[37061] = 25'b1110111100011001100001010;
    rom[37062] = 25'b1110111100011011110100000;
    rom[37063] = 25'b1110111100011110000111000;
    rom[37064] = 25'b1110111100100000011010010;
    rom[37065] = 25'b1110111100100010101101110;
    rom[37066] = 25'b1110111100100101000001110;
    rom[37067] = 25'b1110111100100111010101111;
    rom[37068] = 25'b1110111100101001101010011;
    rom[37069] = 25'b1110111100101011111111000;
    rom[37070] = 25'b1110111100101110010100000;
    rom[37071] = 25'b1110111100110000101001011;
    rom[37072] = 25'b1110111100110010111111000;
    rom[37073] = 25'b1110111100110101010100110;
    rom[37074] = 25'b1110111100110111101010111;
    rom[37075] = 25'b1110111100111010000001011;
    rom[37076] = 25'b1110111100111100011000010;
    rom[37077] = 25'b1110111100111110101111010;
    rom[37078] = 25'b1110111101000001000110100;
    rom[37079] = 25'b1110111101000011011110000;
    rom[37080] = 25'b1110111101000101110101111;
    rom[37081] = 25'b1110111101001000001110001;
    rom[37082] = 25'b1110111101001010100110100;
    rom[37083] = 25'b1110111101001100111111011;
    rom[37084] = 25'b1110111101001111011000010;
    rom[37085] = 25'b1110111101010001110001100;
    rom[37086] = 25'b1110111101010100001011001;
    rom[37087] = 25'b1110111101010110100101000;
    rom[37088] = 25'b1110111101011000111111001;
    rom[37089] = 25'b1110111101011011011001100;
    rom[37090] = 25'b1110111101011101110100010;
    rom[37091] = 25'b1110111101100000001111010;
    rom[37092] = 25'b1110111101100010101010100;
    rom[37093] = 25'b1110111101100101000110001;
    rom[37094] = 25'b1110111101100111100001111;
    rom[37095] = 25'b1110111101101001111110000;
    rom[37096] = 25'b1110111101101100011010011;
    rom[37097] = 25'b1110111101101110110111000;
    rom[37098] = 25'b1110111101110001010011111;
    rom[37099] = 25'b1110111101110011110001001;
    rom[37100] = 25'b1110111101110110001110101;
    rom[37101] = 25'b1110111101111000101100011;
    rom[37102] = 25'b1110111101111011001010100;
    rom[37103] = 25'b1110111101111101101000110;
    rom[37104] = 25'b1110111110000000000111011;
    rom[37105] = 25'b1110111110000010100110001;
    rom[37106] = 25'b1110111110000101000101010;
    rom[37107] = 25'b1110111110000111100100110;
    rom[37108] = 25'b1110111110001010000100011;
    rom[37109] = 25'b1110111110001100100100011;
    rom[37110] = 25'b1110111110001111000100101;
    rom[37111] = 25'b1110111110010001100101001;
    rom[37112] = 25'b1110111110010100000110000;
    rom[37113] = 25'b1110111110010110100111000;
    rom[37114] = 25'b1110111110011001001000011;
    rom[37115] = 25'b1110111110011011101001111;
    rom[37116] = 25'b1110111110011110001011111;
    rom[37117] = 25'b1110111110100000101110000;
    rom[37118] = 25'b1110111110100011010000011;
    rom[37119] = 25'b1110111110100101110011000;
    rom[37120] = 25'b1110111110101000010110000;
    rom[37121] = 25'b1110111110101010111001010;
    rom[37122] = 25'b1110111110101101011100110;
    rom[37123] = 25'b1110111110110000000000100;
    rom[37124] = 25'b1110111110110010100100100;
    rom[37125] = 25'b1110111110110101001000111;
    rom[37126] = 25'b1110111110110111101101011;
    rom[37127] = 25'b1110111110111010010010010;
    rom[37128] = 25'b1110111110111100110111010;
    rom[37129] = 25'b1110111110111111011100110;
    rom[37130] = 25'b1110111111000010000010011;
    rom[37131] = 25'b1110111111000100101000010;
    rom[37132] = 25'b1110111111000111001110100;
    rom[37133] = 25'b1110111111001001110100111;
    rom[37134] = 25'b1110111111001100011011100;
    rom[37135] = 25'b1110111111001111000010100;
    rom[37136] = 25'b1110111111010001101001110;
    rom[37137] = 25'b1110111111010100010001010;
    rom[37138] = 25'b1110111111010110111001000;
    rom[37139] = 25'b1110111111011001100001000;
    rom[37140] = 25'b1110111111011100001001010;
    rom[37141] = 25'b1110111111011110110001110;
    rom[37142] = 25'b1110111111100001011010101;
    rom[37143] = 25'b1110111111100100000011101;
    rom[37144] = 25'b1110111111100110101101000;
    rom[37145] = 25'b1110111111101001010110101;
    rom[37146] = 25'b1110111111101100000000100;
    rom[37147] = 25'b1110111111101110101010100;
    rom[37148] = 25'b1110111111110001010101000;
    rom[37149] = 25'b1110111111110011111111100;
    rom[37150] = 25'b1110111111110110101010100;
    rom[37151] = 25'b1110111111111001010101100;
    rom[37152] = 25'b1110111111111100000001000;
    rom[37153] = 25'b1110111111111110101100101;
    rom[37154] = 25'b1111000000000001011000101;
    rom[37155] = 25'b1111000000000100000100110;
    rom[37156] = 25'b1111000000000110110001001;
    rom[37157] = 25'b1111000000001001011101111;
    rom[37158] = 25'b1111000000001100001010110;
    rom[37159] = 25'b1111000000001110111000000;
    rom[37160] = 25'b1111000000010001100101100;
    rom[37161] = 25'b1111000000010100010011001;
    rom[37162] = 25'b1111000000010111000001001;
    rom[37163] = 25'b1111000000011001101111011;
    rom[37164] = 25'b1111000000011100011101111;
    rom[37165] = 25'b1111000000011111001100100;
    rom[37166] = 25'b1111000000100001111011101;
    rom[37167] = 25'b1111000000100100101010110;
    rom[37168] = 25'b1111000000100111011010011;
    rom[37169] = 25'b1111000000101010001010000;
    rom[37170] = 25'b1111000000101100111010000;
    rom[37171] = 25'b1111000000101111101010010;
    rom[37172] = 25'b1111000000110010011010110;
    rom[37173] = 25'b1111000000110101001011100;
    rom[37174] = 25'b1111000000110111111100100;
    rom[37175] = 25'b1111000000111010101101110;
    rom[37176] = 25'b1111000000111101011111010;
    rom[37177] = 25'b1111000001000000010001000;
    rom[37178] = 25'b1111000001000011000011000;
    rom[37179] = 25'b1111000001000101110101010;
    rom[37180] = 25'b1111000001001000100111110;
    rom[37181] = 25'b1111000001001011011010100;
    rom[37182] = 25'b1111000001001110001101100;
    rom[37183] = 25'b1111000001010001000000110;
    rom[37184] = 25'b1111000001010011110100010;
    rom[37185] = 25'b1111000001010110100111111;
    rom[37186] = 25'b1111000001011001011011111;
    rom[37187] = 25'b1111000001011100010000000;
    rom[37188] = 25'b1111000001011111000100101;
    rom[37189] = 25'b1111000001100001111001010;
    rom[37190] = 25'b1111000001100100101110001;
    rom[37191] = 25'b1111000001100111100011011;
    rom[37192] = 25'b1111000001101010011000110;
    rom[37193] = 25'b1111000001101101001110100;
    rom[37194] = 25'b1111000001110000000100100;
    rom[37195] = 25'b1111000001110010111010101;
    rom[37196] = 25'b1111000001110101110001000;
    rom[37197] = 25'b1111000001111000100111110;
    rom[37198] = 25'b1111000001111011011110100;
    rom[37199] = 25'b1111000001111110010101101;
    rom[37200] = 25'b1111000010000001001101001;
    rom[37201] = 25'b1111000010000100000100101;
    rom[37202] = 25'b1111000010000110111100101;
    rom[37203] = 25'b1111000010001001110100101;
    rom[37204] = 25'b1111000010001100101101000;
    rom[37205] = 25'b1111000010001111100101100;
    rom[37206] = 25'b1111000010010010011110011;
    rom[37207] = 25'b1111000010010101010111011;
    rom[37208] = 25'b1111000010011000010000110;
    rom[37209] = 25'b1111000010011011001010010;
    rom[37210] = 25'b1111000010011110000100000;
    rom[37211] = 25'b1111000010100000111101111;
    rom[37212] = 25'b1111000010100011111000010;
    rom[37213] = 25'b1111000010100110110010101;
    rom[37214] = 25'b1111000010101001101101011;
    rom[37215] = 25'b1111000010101100101000010;
    rom[37216] = 25'b1111000010101111100011100;
    rom[37217] = 25'b1111000010110010011111000;
    rom[37218] = 25'b1111000010110101011010101;
    rom[37219] = 25'b1111000010111000010110100;
    rom[37220] = 25'b1111000010111011010010100;
    rom[37221] = 25'b1111000010111110001110111;
    rom[37222] = 25'b1111000011000001001011100;
    rom[37223] = 25'b1111000011000100001000010;
    rom[37224] = 25'b1111000011000111000101010;
    rom[37225] = 25'b1111000011001010000010101;
    rom[37226] = 25'b1111000011001101000000001;
    rom[37227] = 25'b1111000011001111111101111;
    rom[37228] = 25'b1111000011010010111011110;
    rom[37229] = 25'b1111000011010101111010000;
    rom[37230] = 25'b1111000011011000111000011;
    rom[37231] = 25'b1111000011011011110111000;
    rom[37232] = 25'b1111000011011110110101111;
    rom[37233] = 25'b1111000011100001110101001;
    rom[37234] = 25'b1111000011100100110100011;
    rom[37235] = 25'b1111000011100111110100000;
    rom[37236] = 25'b1111000011101010110011110;
    rom[37237] = 25'b1111000011101101110011110;
    rom[37238] = 25'b1111000011110000110100001;
    rom[37239] = 25'b1111000011110011110100100;
    rom[37240] = 25'b1111000011110110110101010;
    rom[37241] = 25'b1111000011111001110110001;
    rom[37242] = 25'b1111000011111100110111010;
    rom[37243] = 25'b1111000011111111111000101;
    rom[37244] = 25'b1111000100000010111010010;
    rom[37245] = 25'b1111000100000101111100001;
    rom[37246] = 25'b1111000100001000111110001;
    rom[37247] = 25'b1111000100001100000000011;
    rom[37248] = 25'b1111000100001111000010111;
    rom[37249] = 25'b1111000100010010000101101;
    rom[37250] = 25'b1111000100010101001000101;
    rom[37251] = 25'b1111000100011000001011110;
    rom[37252] = 25'b1111000100011011001111001;
    rom[37253] = 25'b1111000100011110010010101;
    rom[37254] = 25'b1111000100100001010110100;
    rom[37255] = 25'b1111000100100100011010101;
    rom[37256] = 25'b1111000100100111011110111;
    rom[37257] = 25'b1111000100101010100011010;
    rom[37258] = 25'b1111000100101101101000000;
    rom[37259] = 25'b1111000100110000101100111;
    rom[37260] = 25'b1111000100110011110010001;
    rom[37261] = 25'b1111000100110110110111011;
    rom[37262] = 25'b1111000100111001111101000;
    rom[37263] = 25'b1111000100111101000010110;
    rom[37264] = 25'b1111000101000000001000110;
    rom[37265] = 25'b1111000101000011001111000;
    rom[37266] = 25'b1111000101000110010101100;
    rom[37267] = 25'b1111000101001001011100001;
    rom[37268] = 25'b1111000101001100100011000;
    rom[37269] = 25'b1111000101001111101010001;
    rom[37270] = 25'b1111000101010010110001011;
    rom[37271] = 25'b1111000101010101111000111;
    rom[37272] = 25'b1111000101011001000000101;
    rom[37273] = 25'b1111000101011100001000101;
    rom[37274] = 25'b1111000101011111010000110;
    rom[37275] = 25'b1111000101100010011001001;
    rom[37276] = 25'b1111000101100101100001110;
    rom[37277] = 25'b1111000101101000101010100;
    rom[37278] = 25'b1111000101101011110011100;
    rom[37279] = 25'b1111000101101110111100110;
    rom[37280] = 25'b1111000101110010000110001;
    rom[37281] = 25'b1111000101110101001111110;
    rom[37282] = 25'b1111000101111000011001101;
    rom[37283] = 25'b1111000101111011100011101;
    rom[37284] = 25'b1111000101111110101110000;
    rom[37285] = 25'b1111000110000001111000011;
    rom[37286] = 25'b1111000110000101000011001;
    rom[37287] = 25'b1111000110001000001110000;
    rom[37288] = 25'b1111000110001011011001001;
    rom[37289] = 25'b1111000110001110100100011;
    rom[37290] = 25'b1111000110010001101111111;
    rom[37291] = 25'b1111000110010100111011101;
    rom[37292] = 25'b1111000110011000000111100;
    rom[37293] = 25'b1111000110011011010011110;
    rom[37294] = 25'b1111000110011110100000000;
    rom[37295] = 25'b1111000110100001101100101;
    rom[37296] = 25'b1111000110100100111001011;
    rom[37297] = 25'b1111000110101000000110011;
    rom[37298] = 25'b1111000110101011010011100;
    rom[37299] = 25'b1111000110101110100000111;
    rom[37300] = 25'b1111000110110001101110011;
    rom[37301] = 25'b1111000110110100111100001;
    rom[37302] = 25'b1111000110111000001010001;
    rom[37303] = 25'b1111000110111011011000011;
    rom[37304] = 25'b1111000110111110100110110;
    rom[37305] = 25'b1111000111000001110101010;
    rom[37306] = 25'b1111000111000101000100000;
    rom[37307] = 25'b1111000111001000010011000;
    rom[37308] = 25'b1111000111001011100010010;
    rom[37309] = 25'b1111000111001110110001100;
    rom[37310] = 25'b1111000111010010000001001;
    rom[37311] = 25'b1111000111010101010000111;
    rom[37312] = 25'b1111000111011000100000111;
    rom[37313] = 25'b1111000111011011110001001;
    rom[37314] = 25'b1111000111011111000001100;
    rom[37315] = 25'b1111000111100010010010000;
    rom[37316] = 25'b1111000111100101100010111;
    rom[37317] = 25'b1111000111101000110011110;
    rom[37318] = 25'b1111000111101100000101000;
    rom[37319] = 25'b1111000111101111010110011;
    rom[37320] = 25'b1111000111110010100111111;
    rom[37321] = 25'b1111000111110101111001101;
    rom[37322] = 25'b1111000111111001001011100;
    rom[37323] = 25'b1111000111111100011101101;
    rom[37324] = 25'b1111000111111111110000000;
    rom[37325] = 25'b1111001000000011000010101;
    rom[37326] = 25'b1111001000000110010101010;
    rom[37327] = 25'b1111001000001001101000010;
    rom[37328] = 25'b1111001000001100111011010;
    rom[37329] = 25'b1111001000010000001110101;
    rom[37330] = 25'b1111001000010011100010001;
    rom[37331] = 25'b1111001000010110110101110;
    rom[37332] = 25'b1111001000011010001001101;
    rom[37333] = 25'b1111001000011101011101110;
    rom[37334] = 25'b1111001000100000110010000;
    rom[37335] = 25'b1111001000100100000110100;
    rom[37336] = 25'b1111001000100111011011001;
    rom[37337] = 25'b1111001000101010101111111;
    rom[37338] = 25'b1111001000101110000100111;
    rom[37339] = 25'b1111001000110001011010001;
    rom[37340] = 25'b1111001000110100101111100;
    rom[37341] = 25'b1111001000111000000101001;
    rom[37342] = 25'b1111001000111011011010111;
    rom[37343] = 25'b1111001000111110110000110;
    rom[37344] = 25'b1111001001000010000111000;
    rom[37345] = 25'b1111001001000101011101010;
    rom[37346] = 25'b1111001001001000110011110;
    rom[37347] = 25'b1111001001001100001010100;
    rom[37348] = 25'b1111001001001111100001011;
    rom[37349] = 25'b1111001001010010111000011;
    rom[37350] = 25'b1111001001010110001111110;
    rom[37351] = 25'b1111001001011001100111001;
    rom[37352] = 25'b1111001001011100111110110;
    rom[37353] = 25'b1111001001100000010110101;
    rom[37354] = 25'b1111001001100011101110100;
    rom[37355] = 25'b1111001001100111000110101;
    rom[37356] = 25'b1111001001101010011111000;
    rom[37357] = 25'b1111001001101101110111100;
    rom[37358] = 25'b1111001001110001010000010;
    rom[37359] = 25'b1111001001110100101001010;
    rom[37360] = 25'b1111001001111000000010010;
    rom[37361] = 25'b1111001001111011011011101;
    rom[37362] = 25'b1111001001111110110101000;
    rom[37363] = 25'b1111001010000010001110100;
    rom[37364] = 25'b1111001010000101101000011;
    rom[37365] = 25'b1111001010001001000010010;
    rom[37366] = 25'b1111001010001100011100100;
    rom[37367] = 25'b1111001010001111110110110;
    rom[37368] = 25'b1111001010010011010001011;
    rom[37369] = 25'b1111001010010110101100000;
    rom[37370] = 25'b1111001010011010000110111;
    rom[37371] = 25'b1111001010011101100001111;
    rom[37372] = 25'b1111001010100000111101001;
    rom[37373] = 25'b1111001010100100011000101;
    rom[37374] = 25'b1111001010100111110100001;
    rom[37375] = 25'b1111001010101011001111111;
    rom[37376] = 25'b1111001010101110101011110;
    rom[37377] = 25'b1111001010110010000111111;
    rom[37378] = 25'b1111001010110101100100001;
    rom[37379] = 25'b1111001010111001000000101;
    rom[37380] = 25'b1111001010111100011101001;
    rom[37381] = 25'b1111001010111111111001111;
    rom[37382] = 25'b1111001011000011010110111;
    rom[37383] = 25'b1111001011000110110100000;
    rom[37384] = 25'b1111001011001010010001011;
    rom[37385] = 25'b1111001011001101101110110;
    rom[37386] = 25'b1111001011010001001100100;
    rom[37387] = 25'b1111001011010100101010010;
    rom[37388] = 25'b1111001011011000001000010;
    rom[37389] = 25'b1111001011011011100110011;
    rom[37390] = 25'b1111001011011111000100101;
    rom[37391] = 25'b1111001011100010100011010;
    rom[37392] = 25'b1111001011100110000001111;
    rom[37393] = 25'b1111001011101001100000101;
    rom[37394] = 25'b1111001011101100111111110;
    rom[37395] = 25'b1111001011110000011110111;
    rom[37396] = 25'b1111001011110011111110001;
    rom[37397] = 25'b1111001011110111011101101;
    rom[37398] = 25'b1111001011111010111101010;
    rom[37399] = 25'b1111001011111110011101001;
    rom[37400] = 25'b1111001100000001111101010;
    rom[37401] = 25'b1111001100000101011101011;
    rom[37402] = 25'b1111001100001000111101101;
    rom[37403] = 25'b1111001100001100011110001;
    rom[37404] = 25'b1111001100001111111110111;
    rom[37405] = 25'b1111001100010011011111101;
    rom[37406] = 25'b1111001100010111000000101;
    rom[37407] = 25'b1111001100011010100001110;
    rom[37408] = 25'b1111001100011110000011000;
    rom[37409] = 25'b1111001100100001100100100;
    rom[37410] = 25'b1111001100100101000110001;
    rom[37411] = 25'b1111001100101000101000000;
    rom[37412] = 25'b1111001100101100001001111;
    rom[37413] = 25'b1111001100101111101100000;
    rom[37414] = 25'b1111001100110011001110010;
    rom[37415] = 25'b1111001100110110110000101;
    rom[37416] = 25'b1111001100111010010011010;
    rom[37417] = 25'b1111001100111101110110000;
    rom[37418] = 25'b1111001101000001011000111;
    rom[37419] = 25'b1111001101000100111100000;
    rom[37420] = 25'b1111001101001000011111010;
    rom[37421] = 25'b1111001101001100000010101;
    rom[37422] = 25'b1111001101001111100110001;
    rom[37423] = 25'b1111001101010011001001110;
    rom[37424] = 25'b1111001101010110101101101;
    rom[37425] = 25'b1111001101011010010001110;
    rom[37426] = 25'b1111001101011101110101111;
    rom[37427] = 25'b1111001101100001011010010;
    rom[37428] = 25'b1111001101100100111110101;
    rom[37429] = 25'b1111001101101000100011011;
    rom[37430] = 25'b1111001101101100001000000;
    rom[37431] = 25'b1111001101101111101101000;
    rom[37432] = 25'b1111001101110011010010001;
    rom[37433] = 25'b1111001101110110110111011;
    rom[37434] = 25'b1111001101111010011100110;
    rom[37435] = 25'b1111001101111110000010010;
    rom[37436] = 25'b1111001110000001101000000;
    rom[37437] = 25'b1111001110000101001101111;
    rom[37438] = 25'b1111001110001000110011111;
    rom[37439] = 25'b1111001110001100011010000;
    rom[37440] = 25'b1111001110010000000000011;
    rom[37441] = 25'b1111001110010011100110110;
    rom[37442] = 25'b1111001110010111001101011;
    rom[37443] = 25'b1111001110011010110100001;
    rom[37444] = 25'b1111001110011110011011000;
    rom[37445] = 25'b1111001110100010000010000;
    rom[37446] = 25'b1111001110100101101001010;
    rom[37447] = 25'b1111001110101001010000101;
    rom[37448] = 25'b1111001110101100111000001;
    rom[37449] = 25'b1111001110110000011111110;
    rom[37450] = 25'b1111001110110100000111100;
    rom[37451] = 25'b1111001110110111101111100;
    rom[37452] = 25'b1111001110111011010111100;
    rom[37453] = 25'b1111001110111110111111110;
    rom[37454] = 25'b1111001111000010101000001;
    rom[37455] = 25'b1111001111000110010000101;
    rom[37456] = 25'b1111001111001001111001010;
    rom[37457] = 25'b1111001111001101100010001;
    rom[37458] = 25'b1111001111010001001011001;
    rom[37459] = 25'b1111001111010100110100001;
    rom[37460] = 25'b1111001111011000011101011;
    rom[37461] = 25'b1111001111011100000110110;
    rom[37462] = 25'b1111001111011111110000010;
    rom[37463] = 25'b1111001111100011011010000;
    rom[37464] = 25'b1111001111100111000011110;
    rom[37465] = 25'b1111001111101010101101101;
    rom[37466] = 25'b1111001111101110010111110;
    rom[37467] = 25'b1111001111110010000010000;
    rom[37468] = 25'b1111001111110101101100010;
    rom[37469] = 25'b1111001111111001010110111;
    rom[37470] = 25'b1111001111111101000001100;
    rom[37471] = 25'b1111010000000000101100010;
    rom[37472] = 25'b1111010000000100010111010;
    rom[37473] = 25'b1111010000001000000010010;
    rom[37474] = 25'b1111010000001011101101011;
    rom[37475] = 25'b1111010000001111011000110;
    rom[37476] = 25'b1111010000010011000100001;
    rom[37477] = 25'b1111010000010110101111110;
    rom[37478] = 25'b1111010000011010011011100;
    rom[37479] = 25'b1111010000011110000111011;
    rom[37480] = 25'b1111010000100001110011011;
    rom[37481] = 25'b1111010000100101011111100;
    rom[37482] = 25'b1111010000101001001011111;
    rom[37483] = 25'b1111010000101100111000010;
    rom[37484] = 25'b1111010000110000100100111;
    rom[37485] = 25'b1111010000110100010001100;
    rom[37486] = 25'b1111010000110111111110010;
    rom[37487] = 25'b1111010000111011101011010;
    rom[37488] = 25'b1111010000111111011000011;
    rom[37489] = 25'b1111010001000011000101100;
    rom[37490] = 25'b1111010001000110110010111;
    rom[37491] = 25'b1111010001001010100000010;
    rom[37492] = 25'b1111010001001110001101111;
    rom[37493] = 25'b1111010001010001111011101;
    rom[37494] = 25'b1111010001010101101001100;
    rom[37495] = 25'b1111010001011001010111100;
    rom[37496] = 25'b1111010001011101000101101;
    rom[37497] = 25'b1111010001100000110011111;
    rom[37498] = 25'b1111010001100100100010010;
    rom[37499] = 25'b1111010001101000010000110;
    rom[37500] = 25'b1111010001101011111111011;
    rom[37501] = 25'b1111010001101111101110001;
    rom[37502] = 25'b1111010001110011011101000;
    rom[37503] = 25'b1111010001110111001100000;
    rom[37504] = 25'b1111010001111010111011001;
    rom[37505] = 25'b1111010001111110101010011;
    rom[37506] = 25'b1111010010000010011001111;
    rom[37507] = 25'b1111010010000110001001011;
    rom[37508] = 25'b1111010010001001111001000;
    rom[37509] = 25'b1111010010001101101000110;
    rom[37510] = 25'b1111010010010001011000101;
    rom[37511] = 25'b1111010010010101001000101;
    rom[37512] = 25'b1111010010011000111000110;
    rom[37513] = 25'b1111010010011100101001001;
    rom[37514] = 25'b1111010010100000011001100;
    rom[37515] = 25'b1111010010100100001001111;
    rom[37516] = 25'b1111010010100111111010101;
    rom[37517] = 25'b1111010010101011101011011;
    rom[37518] = 25'b1111010010101111011100001;
    rom[37519] = 25'b1111010010110011001101010;
    rom[37520] = 25'b1111010010110110111110010;
    rom[37521] = 25'b1111010010111010101111100;
    rom[37522] = 25'b1111010010111110100000111;
    rom[37523] = 25'b1111010011000010010010011;
    rom[37524] = 25'b1111010011000110000011111;
    rom[37525] = 25'b1111010011001001110101101;
    rom[37526] = 25'b1111010011001101100111011;
    rom[37527] = 25'b1111010011010001011001011;
    rom[37528] = 25'b1111010011010101001011011;
    rom[37529] = 25'b1111010011011000111101101;
    rom[37530] = 25'b1111010011011100101111111;
    rom[37531] = 25'b1111010011100000100010010;
    rom[37532] = 25'b1111010011100100010100110;
    rom[37533] = 25'b1111010011101000000111011;
    rom[37534] = 25'b1111010011101011111010010;
    rom[37535] = 25'b1111010011101111101101000;
    rom[37536] = 25'b1111010011110011100000000;
    rom[37537] = 25'b1111010011110111010011001;
    rom[37538] = 25'b1111010011111011000110010;
    rom[37539] = 25'b1111010011111110111001101;
    rom[37540] = 25'b1111010100000010101101001;
    rom[37541] = 25'b1111010100000110100000101;
    rom[37542] = 25'b1111010100001010010100010;
    rom[37543] = 25'b1111010100001110001000000;
    rom[37544] = 25'b1111010100010001111011111;
    rom[37545] = 25'b1111010100010101101111111;
    rom[37546] = 25'b1111010100011001100100000;
    rom[37547] = 25'b1111010100011101011000010;
    rom[37548] = 25'b1111010100100001001100100;
    rom[37549] = 25'b1111010100100101000000111;
    rom[37550] = 25'b1111010100101000110101100;
    rom[37551] = 25'b1111010100101100101010001;
    rom[37552] = 25'b1111010100110000011110111;
    rom[37553] = 25'b1111010100110100010011110;
    rom[37554] = 25'b1111010100111000001000101;
    rom[37555] = 25'b1111010100111011111101110;
    rom[37556] = 25'b1111010100111111110011000;
    rom[37557] = 25'b1111010101000011101000010;
    rom[37558] = 25'b1111010101000111011101110;
    rom[37559] = 25'b1111010101001011010011001;
    rom[37560] = 25'b1111010101001111001000110;
    rom[37561] = 25'b1111010101010010111110011;
    rom[37562] = 25'b1111010101010110110100011;
    rom[37563] = 25'b1111010101011010101010010;
    rom[37564] = 25'b1111010101011110100000001;
    rom[37565] = 25'b1111010101100010010110011;
    rom[37566] = 25'b1111010101100110001100100;
    rom[37567] = 25'b1111010101101010000010111;
    rom[37568] = 25'b1111010101101101111001011;
    rom[37569] = 25'b1111010101110001101111111;
    rom[37570] = 25'b1111010101110101100110100;
    rom[37571] = 25'b1111010101111001011101010;
    rom[37572] = 25'b1111010101111101010100000;
    rom[37573] = 25'b1111010110000001001011000;
    rom[37574] = 25'b1111010110000101000010001;
    rom[37575] = 25'b1111010110001000111001001;
    rom[37576] = 25'b1111010110001100110000011;
    rom[37577] = 25'b1111010110010000100111110;
    rom[37578] = 25'b1111010110010100011111001;
    rom[37579] = 25'b1111010110011000010110110;
    rom[37580] = 25'b1111010110011100001110011;
    rom[37581] = 25'b1111010110100000000110000;
    rom[37582] = 25'b1111010110100011111101111;
    rom[37583] = 25'b1111010110100111110101111;
    rom[37584] = 25'b1111010110101011101101111;
    rom[37585] = 25'b1111010110101111100101111;
    rom[37586] = 25'b1111010110110011011110001;
    rom[37587] = 25'b1111010110110111010110011;
    rom[37588] = 25'b1111010110111011001110111;
    rom[37589] = 25'b1111010110111111000111011;
    rom[37590] = 25'b1111010111000010111111111;
    rom[37591] = 25'b1111010111000110111000100;
    rom[37592] = 25'b1111010111001010110001010;
    rom[37593] = 25'b1111010111001110101010010;
    rom[37594] = 25'b1111010111010010100011001;
    rom[37595] = 25'b1111010111010110011100010;
    rom[37596] = 25'b1111010111011010010101011;
    rom[37597] = 25'b1111010111011110001110100;
    rom[37598] = 25'b1111010111100010000111111;
    rom[37599] = 25'b1111010111100110000001011;
    rom[37600] = 25'b1111010111101001111010111;
    rom[37601] = 25'b1111010111101101110100011;
    rom[37602] = 25'b1111010111110001101110001;
    rom[37603] = 25'b1111010111110101100111111;
    rom[37604] = 25'b1111010111111001100001110;
    rom[37605] = 25'b1111010111111101011011110;
    rom[37606] = 25'b1111011000000001010101110;
    rom[37607] = 25'b1111011000000101001111110;
    rom[37608] = 25'b1111011000001001001010001;
    rom[37609] = 25'b1111011000001101000100011;
    rom[37610] = 25'b1111011000010000111110110;
    rom[37611] = 25'b1111011000010100111001001;
    rom[37612] = 25'b1111011000011000110011110;
    rom[37613] = 25'b1111011000011100101110011;
    rom[37614] = 25'b1111011000100000101001001;
    rom[37615] = 25'b1111011000100100100011111;
    rom[37616] = 25'b1111011000101000011110111;
    rom[37617] = 25'b1111011000101100011001111;
    rom[37618] = 25'b1111011000110000010100111;
    rom[37619] = 25'b1111011000110100010000000;
    rom[37620] = 25'b1111011000111000001011010;
    rom[37621] = 25'b1111011000111100000110100;
    rom[37622] = 25'b1111011001000000000001111;
    rom[37623] = 25'b1111011001000011111101011;
    rom[37624] = 25'b1111011001000111111001000;
    rom[37625] = 25'b1111011001001011110100101;
    rom[37626] = 25'b1111011001001111110000011;
    rom[37627] = 25'b1111011001010011101100001;
    rom[37628] = 25'b1111011001010111101000000;
    rom[37629] = 25'b1111011001011011100011111;
    rom[37630] = 25'b1111011001011111100000000;
    rom[37631] = 25'b1111011001100011011100001;
    rom[37632] = 25'b1111011001100111011000010;
    rom[37633] = 25'b1111011001101011010100101;
    rom[37634] = 25'b1111011001101111010000111;
    rom[37635] = 25'b1111011001110011001101011;
    rom[37636] = 25'b1111011001110111001001111;
    rom[37637] = 25'b1111011001111011000110011;
    rom[37638] = 25'b1111011001111111000011001;
    rom[37639] = 25'b1111011010000010111111110;
    rom[37640] = 25'b1111011010000110111100101;
    rom[37641] = 25'b1111011010001010111001100;
    rom[37642] = 25'b1111011010001110110110100;
    rom[37643] = 25'b1111011010010010110011100;
    rom[37644] = 25'b1111011010010110110000100;
    rom[37645] = 25'b1111011010011010101101110;
    rom[37646] = 25'b1111011010011110101011000;
    rom[37647] = 25'b1111011010100010101000011;
    rom[37648] = 25'b1111011010100110100101110;
    rom[37649] = 25'b1111011010101010100011010;
    rom[37650] = 25'b1111011010101110100000110;
    rom[37651] = 25'b1111011010110010011110011;
    rom[37652] = 25'b1111011010110110011100001;
    rom[37653] = 25'b1111011010111010011001110;
    rom[37654] = 25'b1111011010111110010111101;
    rom[37655] = 25'b1111011011000010010101100;
    rom[37656] = 25'b1111011011000110010011100;
    rom[37657] = 25'b1111011011001010010001100;
    rom[37658] = 25'b1111011011001110001111101;
    rom[37659] = 25'b1111011011010010001101110;
    rom[37660] = 25'b1111011011010110001100000;
    rom[37661] = 25'b1111011011011010001010010;
    rom[37662] = 25'b1111011011011110001000101;
    rom[37663] = 25'b1111011011100010000111001;
    rom[37664] = 25'b1111011011100110000101101;
    rom[37665] = 25'b1111011011101010000100010;
    rom[37666] = 25'b1111011011101110000010111;
    rom[37667] = 25'b1111011011110010000001100;
    rom[37668] = 25'b1111011011110110000000010;
    rom[37669] = 25'b1111011011111001111111001;
    rom[37670] = 25'b1111011011111101111110001;
    rom[37671] = 25'b1111011100000001111101000;
    rom[37672] = 25'b1111011100000101111100001;
    rom[37673] = 25'b1111011100001001111011001;
    rom[37674] = 25'b1111011100001101111010010;
    rom[37675] = 25'b1111011100010001111001100;
    rom[37676] = 25'b1111011100010101111000110;
    rom[37677] = 25'b1111011100011001111000001;
    rom[37678] = 25'b1111011100011101110111100;
    rom[37679] = 25'b1111011100100001110110111;
    rom[37680] = 25'b1111011100100101110110100;
    rom[37681] = 25'b1111011100101001110110000;
    rom[37682] = 25'b1111011100101101110101110;
    rom[37683] = 25'b1111011100110001110101011;
    rom[37684] = 25'b1111011100110101110101001;
    rom[37685] = 25'b1111011100111001110101000;
    rom[37686] = 25'b1111011100111101110100111;
    rom[37687] = 25'b1111011101000001110100110;
    rom[37688] = 25'b1111011101000101110100111;
    rom[37689] = 25'b1111011101001001110100110;
    rom[37690] = 25'b1111011101001101110101000;
    rom[37691] = 25'b1111011101010001110101001;
    rom[37692] = 25'b1111011101010101110101011;
    rom[37693] = 25'b1111011101011001110101101;
    rom[37694] = 25'b1111011101011101110110000;
    rom[37695] = 25'b1111011101100001110110011;
    rom[37696] = 25'b1111011101100101110110110;
    rom[37697] = 25'b1111011101101001110111010;
    rom[37698] = 25'b1111011101101101110111111;
    rom[37699] = 25'b1111011101110001111000100;
    rom[37700] = 25'b1111011101110101111001001;
    rom[37701] = 25'b1111011101111001111001111;
    rom[37702] = 25'b1111011101111101111010101;
    rom[37703] = 25'b1111011110000001111011100;
    rom[37704] = 25'b1111011110000101111100010;
    rom[37705] = 25'b1111011110001001111101001;
    rom[37706] = 25'b1111011110001101111110001;
    rom[37707] = 25'b1111011110010001111111001;
    rom[37708] = 25'b1111011110010110000000010;
    rom[37709] = 25'b1111011110011010000001100;
    rom[37710] = 25'b1111011110011110000010100;
    rom[37711] = 25'b1111011110100010000011111;
    rom[37712] = 25'b1111011110100110000101001;
    rom[37713] = 25'b1111011110101010000110011;
    rom[37714] = 25'b1111011110101110000111110;
    rom[37715] = 25'b1111011110110010001001010;
    rom[37716] = 25'b1111011110110110001010110;
    rom[37717] = 25'b1111011110111010001100001;
    rom[37718] = 25'b1111011110111110001101110;
    rom[37719] = 25'b1111011111000010001111011;
    rom[37720] = 25'b1111011111000110010001000;
    rom[37721] = 25'b1111011111001010010010110;
    rom[37722] = 25'b1111011111001110010100100;
    rom[37723] = 25'b1111011111010010010110010;
    rom[37724] = 25'b1111011111010110011000001;
    rom[37725] = 25'b1111011111011010011010000;
    rom[37726] = 25'b1111011111011110011011111;
    rom[37727] = 25'b1111011111100010011101111;
    rom[37728] = 25'b1111011111100110011111111;
    rom[37729] = 25'b1111011111101010100001111;
    rom[37730] = 25'b1111011111101110100100000;
    rom[37731] = 25'b1111011111110010100110001;
    rom[37732] = 25'b1111011111110110101000011;
    rom[37733] = 25'b1111011111111010101010101;
    rom[37734] = 25'b1111011111111110101100111;
    rom[37735] = 25'b1111100000000010101111001;
    rom[37736] = 25'b1111100000000110110001100;
    rom[37737] = 25'b1111100000001010110011111;
    rom[37738] = 25'b1111100000001110110110010;
    rom[37739] = 25'b1111100000010010111000110;
    rom[37740] = 25'b1111100000010110111011010;
    rom[37741] = 25'b1111100000011010111101110;
    rom[37742] = 25'b1111100000011111000000011;
    rom[37743] = 25'b1111100000100011000011000;
    rom[37744] = 25'b1111100000100111000101101;
    rom[37745] = 25'b1111100000101011001000011;
    rom[37746] = 25'b1111100000101111001011001;
    rom[37747] = 25'b1111100000110011001101111;
    rom[37748] = 25'b1111100000110111010000101;
    rom[37749] = 25'b1111100000111011010011100;
    rom[37750] = 25'b1111100000111111010110011;
    rom[37751] = 25'b1111100001000011011001011;
    rom[37752] = 25'b1111100001000111011100010;
    rom[37753] = 25'b1111100001001011011111010;
    rom[37754] = 25'b1111100001001111100010010;
    rom[37755] = 25'b1111100001010011100101010;
    rom[37756] = 25'b1111100001010111101000100;
    rom[37757] = 25'b1111100001011011101011100;
    rom[37758] = 25'b1111100001011111101110101;
    rom[37759] = 25'b1111100001100011110001111;
    rom[37760] = 25'b1111100001100111110101000;
    rom[37761] = 25'b1111100001101011111000010;
    rom[37762] = 25'b1111100001101111111011101;
    rom[37763] = 25'b1111100001110011111110111;
    rom[37764] = 25'b1111100001111000000010010;
    rom[37765] = 25'b1111100001111100000101101;
    rom[37766] = 25'b1111100010000000001001000;
    rom[37767] = 25'b1111100010000100001100011;
    rom[37768] = 25'b1111100010001000001111111;
    rom[37769] = 25'b1111100010001100010011011;
    rom[37770] = 25'b1111100010010000010110111;
    rom[37771] = 25'b1111100010010100011010011;
    rom[37772] = 25'b1111100010011000011110000;
    rom[37773] = 25'b1111100010011100100001101;
    rom[37774] = 25'b1111100010100000100101010;
    rom[37775] = 25'b1111100010100100101000111;
    rom[37776] = 25'b1111100010101000101100100;
    rom[37777] = 25'b1111100010101100110000010;
    rom[37778] = 25'b1111100010110000110100000;
    rom[37779] = 25'b1111100010110100110111101;
    rom[37780] = 25'b1111100010111000111011100;
    rom[37781] = 25'b1111100010111100111111010;
    rom[37782] = 25'b1111100011000001000011001;
    rom[37783] = 25'b1111100011000101000111000;
    rom[37784] = 25'b1111100011001001001010111;
    rom[37785] = 25'b1111100011001101001110110;
    rom[37786] = 25'b1111100011010001010010101;
    rom[37787] = 25'b1111100011010101010110101;
    rom[37788] = 25'b1111100011011001011010100;
    rom[37789] = 25'b1111100011011101011110100;
    rom[37790] = 25'b1111100011100001100010101;
    rom[37791] = 25'b1111100011100101100110101;
    rom[37792] = 25'b1111100011101001101010110;
    rom[37793] = 25'b1111100011101101101110110;
    rom[37794] = 25'b1111100011110001110010111;
    rom[37795] = 25'b1111100011110101110111000;
    rom[37796] = 25'b1111100011111001111011001;
    rom[37797] = 25'b1111100011111101111111010;
    rom[37798] = 25'b1111100100000010000011011;
    rom[37799] = 25'b1111100100000110000111101;
    rom[37800] = 25'b1111100100001010001011111;
    rom[37801] = 25'b1111100100001110010000000;
    rom[37802] = 25'b1111100100010010010100010;
    rom[37803] = 25'b1111100100010110011000100;
    rom[37804] = 25'b1111100100011010011100111;
    rom[37805] = 25'b1111100100011110100001001;
    rom[37806] = 25'b1111100100100010100101011;
    rom[37807] = 25'b1111100100100110101001110;
    rom[37808] = 25'b1111100100101010101110001;
    rom[37809] = 25'b1111100100101110110010100;
    rom[37810] = 25'b1111100100110010110110110;
    rom[37811] = 25'b1111100100110110111011001;
    rom[37812] = 25'b1111100100111010111111100;
    rom[37813] = 25'b1111100100111111000100000;
    rom[37814] = 25'b1111100101000011001000011;
    rom[37815] = 25'b1111100101000111001100111;
    rom[37816] = 25'b1111100101001011010001010;
    rom[37817] = 25'b1111100101001111010101110;
    rom[37818] = 25'b1111100101010011011010001;
    rom[37819] = 25'b1111100101010111011110101;
    rom[37820] = 25'b1111100101011011100011010;
    rom[37821] = 25'b1111100101011111100111101;
    rom[37822] = 25'b1111100101100011101100010;
    rom[37823] = 25'b1111100101100111110000110;
    rom[37824] = 25'b1111100101101011110101010;
    rom[37825] = 25'b1111100101101111111001110;
    rom[37826] = 25'b1111100101110011111110010;
    rom[37827] = 25'b1111100101111000000010111;
    rom[37828] = 25'b1111100101111100000111100;
    rom[37829] = 25'b1111100110000000001100000;
    rom[37830] = 25'b1111100110000100010000101;
    rom[37831] = 25'b1111100110001000010101010;
    rom[37832] = 25'b1111100110001100011001110;
    rom[37833] = 25'b1111100110010000011110011;
    rom[37834] = 25'b1111100110010100100011001;
    rom[37835] = 25'b1111100110011000100111101;
    rom[37836] = 25'b1111100110011100101100010;
    rom[37837] = 25'b1111100110100000110000111;
    rom[37838] = 25'b1111100110100100110101100;
    rom[37839] = 25'b1111100110101000111010010;
    rom[37840] = 25'b1111100110101100111110111;
    rom[37841] = 25'b1111100110110001000011100;
    rom[37842] = 25'b1111100110110101001000001;
    rom[37843] = 25'b1111100110111001001100110;
    rom[37844] = 25'b1111100110111101010001011;
    rom[37845] = 25'b1111100111000001010110000;
    rom[37846] = 25'b1111100111000101011010110;
    rom[37847] = 25'b1111100111001001011111011;
    rom[37848] = 25'b1111100111001101100100001;
    rom[37849] = 25'b1111100111010001101000110;
    rom[37850] = 25'b1111100111010101101101011;
    rom[37851] = 25'b1111100111011001110010000;
    rom[37852] = 25'b1111100111011101110110110;
    rom[37853] = 25'b1111100111100001111011011;
    rom[37854] = 25'b1111100111100110000000000;
    rom[37855] = 25'b1111100111101010000100101;
    rom[37856] = 25'b1111100111101110001001011;
    rom[37857] = 25'b1111100111110010001110000;
    rom[37858] = 25'b1111100111110110010010110;
    rom[37859] = 25'b1111100111111010010111011;
    rom[37860] = 25'b1111100111111110011100000;
    rom[37861] = 25'b1111101000000010100000101;
    rom[37862] = 25'b1111101000000110100101010;
    rom[37863] = 25'b1111101000001010101001111;
    rom[37864] = 25'b1111101000001110101110100;
    rom[37865] = 25'b1111101000010010110011010;
    rom[37866] = 25'b1111101000010110110111111;
    rom[37867] = 25'b1111101000011010111100100;
    rom[37868] = 25'b1111101000011111000001000;
    rom[37869] = 25'b1111101000100011000101101;
    rom[37870] = 25'b1111101000100111001010011;
    rom[37871] = 25'b1111101000101011001110111;
    rom[37872] = 25'b1111101000101111010011100;
    rom[37873] = 25'b1111101000110011011000000;
    rom[37874] = 25'b1111101000110111011100110;
    rom[37875] = 25'b1111101000111011100001010;
    rom[37876] = 25'b1111101000111111100101110;
    rom[37877] = 25'b1111101001000011101010011;
    rom[37878] = 25'b1111101001000111101110111;
    rom[37879] = 25'b1111101001001011110011100;
    rom[37880] = 25'b1111101001001111111000000;
    rom[37881] = 25'b1111101001010011111100100;
    rom[37882] = 25'b1111101001011000000001000;
    rom[37883] = 25'b1111101001011100000101100;
    rom[37884] = 25'b1111101001100000001010000;
    rom[37885] = 25'b1111101001100100001110100;
    rom[37886] = 25'b1111101001101000010010111;
    rom[37887] = 25'b1111101001101100010111011;
    rom[37888] = 25'b1111101001110000011011111;
    rom[37889] = 25'b1111101001110100100000010;
    rom[37890] = 25'b1111101001111000100100101;
    rom[37891] = 25'b1111101001111100101001001;
    rom[37892] = 25'b1111101010000000101101100;
    rom[37893] = 25'b1111101010000100110001111;
    rom[37894] = 25'b1111101010001000110110010;
    rom[37895] = 25'b1111101010001100111010101;
    rom[37896] = 25'b1111101010010000111110111;
    rom[37897] = 25'b1111101010010101000011010;
    rom[37898] = 25'b1111101010011001000111101;
    rom[37899] = 25'b1111101010011101001011111;
    rom[37900] = 25'b1111101010100001010000001;
    rom[37901] = 25'b1111101010100101010100011;
    rom[37902] = 25'b1111101010101001011000100;
    rom[37903] = 25'b1111101010101101011100111;
    rom[37904] = 25'b1111101010110001100001000;
    rom[37905] = 25'b1111101010110101100101001;
    rom[37906] = 25'b1111101010111001101001011;
    rom[37907] = 25'b1111101010111101101101100;
    rom[37908] = 25'b1111101011000001110001110;
    rom[37909] = 25'b1111101011000101110101110;
    rom[37910] = 25'b1111101011001001111001111;
    rom[37911] = 25'b1111101011001101111110000;
    rom[37912] = 25'b1111101011010010000010000;
    rom[37913] = 25'b1111101011010110000110000;
    rom[37914] = 25'b1111101011011010001010000;
    rom[37915] = 25'b1111101011011110001110000;
    rom[37916] = 25'b1111101011100010010010000;
    rom[37917] = 25'b1111101011100110010110000;
    rom[37918] = 25'b1111101011101010011001111;
    rom[37919] = 25'b1111101011101110011101110;
    rom[37920] = 25'b1111101011110010100001101;
    rom[37921] = 25'b1111101011110110100101101;
    rom[37922] = 25'b1111101011111010101001011;
    rom[37923] = 25'b1111101011111110101101001;
    rom[37924] = 25'b1111101100000010110001000;
    rom[37925] = 25'b1111101100000110110100110;
    rom[37926] = 25'b1111101100001010111000100;
    rom[37927] = 25'b1111101100001110111100010;
    rom[37928] = 25'b1111101100010010111111111;
    rom[37929] = 25'b1111101100010111000011100;
    rom[37930] = 25'b1111101100011011000111001;
    rom[37931] = 25'b1111101100011111001010110;
    rom[37932] = 25'b1111101100100011001110011;
    rom[37933] = 25'b1111101100100111010001111;
    rom[37934] = 25'b1111101100101011010101100;
    rom[37935] = 25'b1111101100101111011000111;
    rom[37936] = 25'b1111101100110011011100100;
    rom[37937] = 25'b1111101100110111011111111;
    rom[37938] = 25'b1111101100111011100011011;
    rom[37939] = 25'b1111101100111111100110110;
    rom[37940] = 25'b1111101101000011101010001;
    rom[37941] = 25'b1111101101000111101101011;
    rom[37942] = 25'b1111101101001011110000101;
    rom[37943] = 25'b1111101101001111110100000;
    rom[37944] = 25'b1111101101010011110111010;
    rom[37945] = 25'b1111101101010111111010011;
    rom[37946] = 25'b1111101101011011111101101;
    rom[37947] = 25'b1111101101100000000000110;
    rom[37948] = 25'b1111101101100100000011111;
    rom[37949] = 25'b1111101101101000000111000;
    rom[37950] = 25'b1111101101101100001010000;
    rom[37951] = 25'b1111101101110000001101000;
    rom[37952] = 25'b1111101101110100010000000;
    rom[37953] = 25'b1111101101111000010011000;
    rom[37954] = 25'b1111101101111100010101111;
    rom[37955] = 25'b1111101110000000011000110;
    rom[37956] = 25'b1111101110000100011011101;
    rom[37957] = 25'b1111101110001000011110011;
    rom[37958] = 25'b1111101110001100100001010;
    rom[37959] = 25'b1111101110010000100100000;
    rom[37960] = 25'b1111101110010100100110110;
    rom[37961] = 25'b1111101110011000101001011;
    rom[37962] = 25'b1111101110011100101100000;
    rom[37963] = 25'b1111101110100000101110101;
    rom[37964] = 25'b1111101110100100110001001;
    rom[37965] = 25'b1111101110101000110011101;
    rom[37966] = 25'b1111101110101100110110001;
    rom[37967] = 25'b1111101110110000111000101;
    rom[37968] = 25'b1111101110110100111011000;
    rom[37969] = 25'b1111101110111000111101100;
    rom[37970] = 25'b1111101110111100111111110;
    rom[37971] = 25'b1111101111000001000010001;
    rom[37972] = 25'b1111101111000101000100010;
    rom[37973] = 25'b1111101111001001000110100;
    rom[37974] = 25'b1111101111001101001000110;
    rom[37975] = 25'b1111101111010001001010111;
    rom[37976] = 25'b1111101111010101001101000;
    rom[37977] = 25'b1111101111011001001111000;
    rom[37978] = 25'b1111101111011101010001000;
    rom[37979] = 25'b1111101111100001010011000;
    rom[37980] = 25'b1111101111100101010101000;
    rom[37981] = 25'b1111101111101001010110111;
    rom[37982] = 25'b1111101111101101011000101;
    rom[37983] = 25'b1111101111110001011010100;
    rom[37984] = 25'b1111101111110101011100010;
    rom[37985] = 25'b1111101111111001011110000;
    rom[37986] = 25'b1111101111111101011111101;
    rom[37987] = 25'b1111110000000001100001011;
    rom[37988] = 25'b1111110000000101100010111;
    rom[37989] = 25'b1111110000001001100100100;
    rom[37990] = 25'b1111110000001101100101111;
    rom[37991] = 25'b1111110000010001100111011;
    rom[37992] = 25'b1111110000010101101000110;
    rom[37993] = 25'b1111110000011001101010001;
    rom[37994] = 25'b1111110000011101101011011;
    rom[37995] = 25'b1111110000100001101100110;
    rom[37996] = 25'b1111110000100101101110000;
    rom[37997] = 25'b1111110000101001101111001;
    rom[37998] = 25'b1111110000101101110000010;
    rom[37999] = 25'b1111110000110001110001010;
    rom[38000] = 25'b1111110000110101110010011;
    rom[38001] = 25'b1111110000111001110011011;
    rom[38002] = 25'b1111110000111101110100010;
    rom[38003] = 25'b1111110001000001110101001;
    rom[38004] = 25'b1111110001000101110110000;
    rom[38005] = 25'b1111110001001001110110110;
    rom[38006] = 25'b1111110001001101110111100;
    rom[38007] = 25'b1111110001010001111000001;
    rom[38008] = 25'b1111110001010101111000110;
    rom[38009] = 25'b1111110001011001111001011;
    rom[38010] = 25'b1111110001011101111001111;
    rom[38011] = 25'b1111110001100001111010011;
    rom[38012] = 25'b1111110001100101111010111;
    rom[38013] = 25'b1111110001101001111011001;
    rom[38014] = 25'b1111110001101101111011100;
    rom[38015] = 25'b1111110001110001111011110;
    rom[38016] = 25'b1111110001110101111100000;
    rom[38017] = 25'b1111110001111001111100001;
    rom[38018] = 25'b1111110001111101111100010;
    rom[38019] = 25'b1111110010000001111100010;
    rom[38020] = 25'b1111110010000101111100010;
    rom[38021] = 25'b1111110010001001111100010;
    rom[38022] = 25'b1111110010001101111100001;
    rom[38023] = 25'b1111110010010001111100000;
    rom[38024] = 25'b1111110010010101111011110;
    rom[38025] = 25'b1111110010011001111011100;
    rom[38026] = 25'b1111110010011101111011001;
    rom[38027] = 25'b1111110010100001111010110;
    rom[38028] = 25'b1111110010100101111010010;
    rom[38029] = 25'b1111110010101001111001110;
    rom[38030] = 25'b1111110010101101111001010;
    rom[38031] = 25'b1111110010110001111000101;
    rom[38032] = 25'b1111110010110101111000000;
    rom[38033] = 25'b1111110010111001110111001;
    rom[38034] = 25'b1111110010111101110110011;
    rom[38035] = 25'b1111110011000001110101100;
    rom[38036] = 25'b1111110011000101110100101;
    rom[38037] = 25'b1111110011001001110011110;
    rom[38038] = 25'b1111110011001101110010101;
    rom[38039] = 25'b1111110011010001110001100;
    rom[38040] = 25'b1111110011010101110000011;
    rom[38041] = 25'b1111110011011001101111010;
    rom[38042] = 25'b1111110011011101101101111;
    rom[38043] = 25'b1111110011100001101100100;
    rom[38044] = 25'b1111110011100101101011010;
    rom[38045] = 25'b1111110011101001101001110;
    rom[38046] = 25'b1111110011101101101000001;
    rom[38047] = 25'b1111110011110001100110101;
    rom[38048] = 25'b1111110011110101100101000;
    rom[38049] = 25'b1111110011111001100011010;
    rom[38050] = 25'b1111110011111101100001100;
    rom[38051] = 25'b1111110100000001011111101;
    rom[38052] = 25'b1111110100000101011101110;
    rom[38053] = 25'b1111110100001001011011110;
    rom[38054] = 25'b1111110100001101011001110;
    rom[38055] = 25'b1111110100010001010111110;
    rom[38056] = 25'b1111110100010101010101100;
    rom[38057] = 25'b1111110100011001010011010;
    rom[38058] = 25'b1111110100011101010001000;
    rom[38059] = 25'b1111110100100001001110101;
    rom[38060] = 25'b1111110100100101001100001;
    rom[38061] = 25'b1111110100101001001001110;
    rom[38062] = 25'b1111110100101101000111001;
    rom[38063] = 25'b1111110100110001000100100;
    rom[38064] = 25'b1111110100110101000001110;
    rom[38065] = 25'b1111110100111000111111000;
    rom[38066] = 25'b1111110100111100111100010;
    rom[38067] = 25'b1111110101000000111001010;
    rom[38068] = 25'b1111110101000100110110011;
    rom[38069] = 25'b1111110101001000110011011;
    rom[38070] = 25'b1111110101001100110000010;
    rom[38071] = 25'b1111110101010000101101001;
    rom[38072] = 25'b1111110101010100101001110;
    rom[38073] = 25'b1111110101011000100110100;
    rom[38074] = 25'b1111110101011100100011001;
    rom[38075] = 25'b1111110101100000011111101;
    rom[38076] = 25'b1111110101100100011100001;
    rom[38077] = 25'b1111110101101000011000100;
    rom[38078] = 25'b1111110101101100010100111;
    rom[38079] = 25'b1111110101110000010001001;
    rom[38080] = 25'b1111110101110100001101010;
    rom[38081] = 25'b1111110101111000001001011;
    rom[38082] = 25'b1111110101111100000101100;
    rom[38083] = 25'b1111110110000000000001011;
    rom[38084] = 25'b1111110110000011111101010;
    rom[38085] = 25'b1111110110000111111001001;
    rom[38086] = 25'b1111110110001011110100111;
    rom[38087] = 25'b1111110110001111110000100;
    rom[38088] = 25'b1111110110010011101100001;
    rom[38089] = 25'b1111110110010111100111101;
    rom[38090] = 25'b1111110110011011100011001;
    rom[38091] = 25'b1111110110011111011110100;
    rom[38092] = 25'b1111110110100011011001110;
    rom[38093] = 25'b1111110110100111010101000;
    rom[38094] = 25'b1111110110101011010000001;
    rom[38095] = 25'b1111110110101111001011001;
    rom[38096] = 25'b1111110110110011000110001;
    rom[38097] = 25'b1111110110110111000001001;
    rom[38098] = 25'b1111110110111010111011111;
    rom[38099] = 25'b1111110110111110110110101;
    rom[38100] = 25'b1111110111000010110001011;
    rom[38101] = 25'b1111110111000110101011111;
    rom[38102] = 25'b1111110111001010100110011;
    rom[38103] = 25'b1111110111001110100000110;
    rom[38104] = 25'b1111110111010010011011001;
    rom[38105] = 25'b1111110111010110010101100;
    rom[38106] = 25'b1111110111011010001111110;
    rom[38107] = 25'b1111110111011110001001111;
    rom[38108] = 25'b1111110111100010000011110;
    rom[38109] = 25'b1111110111100101111101110;
    rom[38110] = 25'b1111110111101001110111101;
    rom[38111] = 25'b1111110111101101110001011;
    rom[38112] = 25'b1111110111110001101011001;
    rom[38113] = 25'b1111110111110101100100110;
    rom[38114] = 25'b1111110111111001011110011;
    rom[38115] = 25'b1111110111111101010111111;
    rom[38116] = 25'b1111111000000001010001001;
    rom[38117] = 25'b1111111000000101001010100;
    rom[38118] = 25'b1111111000001001000011101;
    rom[38119] = 25'b1111111000001100111100111;
    rom[38120] = 25'b1111111000010000110101111;
    rom[38121] = 25'b1111111000010100101110111;
    rom[38122] = 25'b1111111000011000100111110;
    rom[38123] = 25'b1111111000011100100000100;
    rom[38124] = 25'b1111111000100000011001010;
    rom[38125] = 25'b1111111000100100010001111;
    rom[38126] = 25'b1111111000101000001010011;
    rom[38127] = 25'b1111111000101100000010111;
    rom[38128] = 25'b1111111000101111111011010;
    rom[38129] = 25'b1111111000110011110011100;
    rom[38130] = 25'b1111111000110111101011101;
    rom[38131] = 25'b1111111000111011100011110;
    rom[38132] = 25'b1111111000111111011011111;
    rom[38133] = 25'b1111111001000011010011110;
    rom[38134] = 25'b1111111001000111001011101;
    rom[38135] = 25'b1111111001001011000011011;
    rom[38136] = 25'b1111111001001110111011000;
    rom[38137] = 25'b1111111001010010110010101;
    rom[38138] = 25'b1111111001010110101010001;
    rom[38139] = 25'b1111111001011010100001100;
    rom[38140] = 25'b1111111001011110011000111;
    rom[38141] = 25'b1111111001100010010000000;
    rom[38142] = 25'b1111111001100110000111001;
    rom[38143] = 25'b1111111001101001111110001;
    rom[38144] = 25'b1111111001101101110101001;
    rom[38145] = 25'b1111111001110001101100000;
    rom[38146] = 25'b1111111001110101100010110;
    rom[38147] = 25'b1111111001111001011001100;
    rom[38148] = 25'b1111111001111101010000001;
    rom[38149] = 25'b1111111010000001000110100;
    rom[38150] = 25'b1111111010000100111100111;
    rom[38151] = 25'b1111111010001000110011010;
    rom[38152] = 25'b1111111010001100101001011;
    rom[38153] = 25'b1111111010010000011111101;
    rom[38154] = 25'b1111111010010100010101100;
    rom[38155] = 25'b1111111010011000001011100;
    rom[38156] = 25'b1111111010011100000001011;
    rom[38157] = 25'b1111111010011111110111001;
    rom[38158] = 25'b1111111010100011101100110;
    rom[38159] = 25'b1111111010100111100010011;
    rom[38160] = 25'b1111111010101011010111110;
    rom[38161] = 25'b1111111010101111001101001;
    rom[38162] = 25'b1111111010110011000010011;
    rom[38163] = 25'b1111111010110110110111100;
    rom[38164] = 25'b1111111010111010101100110;
    rom[38165] = 25'b1111111010111110100001101;
    rom[38166] = 25'b1111111011000010010110100;
    rom[38167] = 25'b1111111011000110001011010;
    rom[38168] = 25'b1111111011001010000000000;
    rom[38169] = 25'b1111111011001101110100101;
    rom[38170] = 25'b1111111011010001101001001;
    rom[38171] = 25'b1111111011010101011101100;
    rom[38172] = 25'b1111111011011001010001111;
    rom[38173] = 25'b1111111011011101000110000;
    rom[38174] = 25'b1111111011100000111010001;
    rom[38175] = 25'b1111111011100100101110000;
    rom[38176] = 25'b1111111011101000100010000;
    rom[38177] = 25'b1111111011101100010101111;
    rom[38178] = 25'b1111111011110000001001100;
    rom[38179] = 25'b1111111011110011111101001;
    rom[38180] = 25'b1111111011110111110000101;
    rom[38181] = 25'b1111111011111011100100000;
    rom[38182] = 25'b1111111011111111010111010;
    rom[38183] = 25'b1111111100000011001010100;
    rom[38184] = 25'b1111111100000110111101101;
    rom[38185] = 25'b1111111100001010110000101;
    rom[38186] = 25'b1111111100001110100011100;
    rom[38187] = 25'b1111111100010010010110010;
    rom[38188] = 25'b1111111100010110001001000;
    rom[38189] = 25'b1111111100011001111011100;
    rom[38190] = 25'b1111111100011101101110000;
    rom[38191] = 25'b1111111100100001100000011;
    rom[38192] = 25'b1111111100100101010010110;
    rom[38193] = 25'b1111111100101001000100111;
    rom[38194] = 25'b1111111100101100110110111;
    rom[38195] = 25'b1111111100110000101000111;
    rom[38196] = 25'b1111111100110100011010110;
    rom[38197] = 25'b1111111100111000001100100;
    rom[38198] = 25'b1111111100111011111110001;
    rom[38199] = 25'b1111111100111111101111101;
    rom[38200] = 25'b1111111101000011100001001;
    rom[38201] = 25'b1111111101000111010010100;
    rom[38202] = 25'b1111111101001011000011101;
    rom[38203] = 25'b1111111101001110110100110;
    rom[38204] = 25'b1111111101010010100101110;
    rom[38205] = 25'b1111111101010110010110101;
    rom[38206] = 25'b1111111101011010000111011;
    rom[38207] = 25'b1111111101011101111000001;
    rom[38208] = 25'b1111111101100001101000110;
    rom[38209] = 25'b1111111101100101011001010;
    rom[38210] = 25'b1111111101101001001001101;
    rom[38211] = 25'b1111111101101100111001110;
    rom[38212] = 25'b1111111101110000101010000;
    rom[38213] = 25'b1111111101110100011010000;
    rom[38214] = 25'b1111111101111000001001111;
    rom[38215] = 25'b1111111101111011111001110;
    rom[38216] = 25'b1111111101111111101001011;
    rom[38217] = 25'b1111111110000011011001000;
    rom[38218] = 25'b1111111110000111001000100;
    rom[38219] = 25'b1111111110001010110111111;
    rom[38220] = 25'b1111111110001110100111001;
    rom[38221] = 25'b1111111110010010010110010;
    rom[38222] = 25'b1111111110010110000101011;
    rom[38223] = 25'b1111111110011001110100010;
    rom[38224] = 25'b1111111110011101100011001;
    rom[38225] = 25'b1111111110100001010001111;
    rom[38226] = 25'b1111111110100101000000011;
    rom[38227] = 25'b1111111110101000101110111;
    rom[38228] = 25'b1111111110101100011101010;
    rom[38229] = 25'b1111111110110000001011100;
    rom[38230] = 25'b1111111110110011111001101;
    rom[38231] = 25'b1111111110110111100111101;
    rom[38232] = 25'b1111111110111011010101100;
    rom[38233] = 25'b1111111110111111000011010;
    rom[38234] = 25'b1111111111000010110001000;
    rom[38235] = 25'b1111111111000110011110100;
    rom[38236] = 25'b1111111111001010001100000;
    rom[38237] = 25'b1111111111001101111001010;
    rom[38238] = 25'b1111111111010001100110101;
    rom[38239] = 25'b1111111111010101010011110;
    rom[38240] = 25'b1111111111011001000000101;
    rom[38241] = 25'b1111111111011100101101100;
    rom[38242] = 25'b1111111111100000011010010;
    rom[38243] = 25'b1111111111100100000111000;
    rom[38244] = 25'b1111111111100111110011011;
    rom[38245] = 25'b1111111111101011011111111;
    rom[38246] = 25'b1111111111101111001100001;
    rom[38247] = 25'b1111111111110010111000010;
    rom[38248] = 25'b1111111111110110100100011;
    rom[38249] = 25'b1111111111111010010000010;
    rom[38250] = 25'b1111111111111101111100001;
    rom[38251] = 25'b0000000000000001100111110;
    rom[38252] = 25'b0000000000000101010011010;
    rom[38253] = 25'b0000000000001000111110110;
    rom[38254] = 25'b0000000000001100101010001;
    rom[38255] = 25'b0000000000010000010101010;
    rom[38256] = 25'b0000000000010100000000011;
    rom[38257] = 25'b0000000000010111101011011;
    rom[38258] = 25'b0000000000011011010110010;
    rom[38259] = 25'b0000000000011111000000111;
    rom[38260] = 25'b0000000000100010101011100;
    rom[38261] = 25'b0000000000100110010110000;
    rom[38262] = 25'b0000000000101010000000011;
    rom[38263] = 25'b0000000000101101101010101;
    rom[38264] = 25'b0000000000110001010100110;
    rom[38265] = 25'b0000000000110100111110110;
    rom[38266] = 25'b0000000000111000101000101;
    rom[38267] = 25'b0000000000111100010010011;
    rom[38268] = 25'b0000000000111111111100000;
    rom[38269] = 25'b0000000001000011100101011;
    rom[38270] = 25'b0000000001000111001110111;
    rom[38271] = 25'b0000000001001010111000001;
    rom[38272] = 25'b0000000001001110100001010;
    rom[38273] = 25'b0000000001010010001010010;
    rom[38274] = 25'b0000000001010101110011010;
    rom[38275] = 25'b0000000001011001011011111;
    rom[38276] = 25'b0000000001011101000100100;
    rom[38277] = 25'b0000000001100000101101001;
    rom[38278] = 25'b0000000001100100010101011;
    rom[38279] = 25'b0000000001100111111101101;
    rom[38280] = 25'b0000000001101011100101111;
    rom[38281] = 25'b0000000001101111001101111;
    rom[38282] = 25'b0000000001110010110101110;
    rom[38283] = 25'b0000000001110110011101100;
    rom[38284] = 25'b0000000001111010000101001;
    rom[38285] = 25'b0000000001111101101100101;
    rom[38286] = 25'b0000000010000001010100000;
    rom[38287] = 25'b0000000010000100111011010;
    rom[38288] = 25'b0000000010001000100010011;
    rom[38289] = 25'b0000000010001100001001010;
    rom[38290] = 25'b0000000010001111110000001;
    rom[38291] = 25'b0000000010010011010110111;
    rom[38292] = 25'b0000000010010110111101100;
    rom[38293] = 25'b0000000010011010100100000;
    rom[38294] = 25'b0000000010011110001010011;
    rom[38295] = 25'b0000000010100001110000100;
    rom[38296] = 25'b0000000010100101010110101;
    rom[38297] = 25'b0000000010101000111100101;
    rom[38298] = 25'b0000000010101100100010011;
    rom[38299] = 25'b0000000010110000001000001;
    rom[38300] = 25'b0000000010110011101101101;
    rom[38301] = 25'b0000000010110111010011001;
    rom[38302] = 25'b0000000010111010111000011;
    rom[38303] = 25'b0000000010111110011101100;
    rom[38304] = 25'b0000000011000010000010100;
    rom[38305] = 25'b0000000011000101100111100;
    rom[38306] = 25'b0000000011001001001100010;
    rom[38307] = 25'b0000000011001100110001000;
    rom[38308] = 25'b0000000011010000010101011;
    rom[38309] = 25'b0000000011010011111001110;
    rom[38310] = 25'b0000000011010111011110000;
    rom[38311] = 25'b0000000011011011000010001;
    rom[38312] = 25'b0000000011011110100110001;
    rom[38313] = 25'b0000000011100010001001111;
    rom[38314] = 25'b0000000011100101101101101;
    rom[38315] = 25'b0000000011101001010001001;
    rom[38316] = 25'b0000000011101100110100101;
    rom[38317] = 25'b0000000011110000011000000;
    rom[38318] = 25'b0000000011110011111011001;
    rom[38319] = 25'b0000000011110111011110001;
    rom[38320] = 25'b0000000011111011000001000;
    rom[38321] = 25'b0000000011111110100011110;
    rom[38322] = 25'b0000000100000010000110011;
    rom[38323] = 25'b0000000100000101101000111;
    rom[38324] = 25'b0000000100001001001011010;
    rom[38325] = 25'b0000000100001100101101011;
    rom[38326] = 25'b0000000100010000001111100;
    rom[38327] = 25'b0000000100010011110001011;
    rom[38328] = 25'b0000000100010111010011010;
    rom[38329] = 25'b0000000100011010110101000;
    rom[38330] = 25'b0000000100011110010110100;
    rom[38331] = 25'b0000000100100001110111111;
    rom[38332] = 25'b0000000100100101011001001;
    rom[38333] = 25'b0000000100101000111010010;
    rom[38334] = 25'b0000000100101100011011010;
    rom[38335] = 25'b0000000100101111111100000;
    rom[38336] = 25'b0000000100110011011100101;
    rom[38337] = 25'b0000000100110110111101010;
    rom[38338] = 25'b0000000100111010011101101;
    rom[38339] = 25'b0000000100111101111101111;
    rom[38340] = 25'b0000000101000001011110000;
    rom[38341] = 25'b0000000101000100111110001;
    rom[38342] = 25'b0000000101001000011101111;
    rom[38343] = 25'b0000000101001011111101101;
    rom[38344] = 25'b0000000101001111011101010;
    rom[38345] = 25'b0000000101010010111100101;
    rom[38346] = 25'b0000000101010110011011111;
    rom[38347] = 25'b0000000101011001111011001;
    rom[38348] = 25'b0000000101011101011010001;
    rom[38349] = 25'b0000000101100000111000111;
    rom[38350] = 25'b0000000101100100010111101;
    rom[38351] = 25'b0000000101100111110110010;
    rom[38352] = 25'b0000000101101011010100101;
    rom[38353] = 25'b0000000101101110110010111;
    rom[38354] = 25'b0000000101110010010001001;
    rom[38355] = 25'b0000000101110101101111001;
    rom[38356] = 25'b0000000101111001001101000;
    rom[38357] = 25'b0000000101111100101010101;
    rom[38358] = 25'b0000000110000000001000010;
    rom[38359] = 25'b0000000110000011100101101;
    rom[38360] = 25'b0000000110000111000011000;
    rom[38361] = 25'b0000000110001010100000001;
    rom[38362] = 25'b0000000110001101111101001;
    rom[38363] = 25'b0000000110010001011010000;
    rom[38364] = 25'b0000000110010100110110101;
    rom[38365] = 25'b0000000110011000010011010;
    rom[38366] = 25'b0000000110011011101111101;
    rom[38367] = 25'b0000000110011111001011111;
    rom[38368] = 25'b0000000110100010101000000;
    rom[38369] = 25'b0000000110100110000100000;
    rom[38370] = 25'b0000000110101001011111110;
    rom[38371] = 25'b0000000110101100111011100;
    rom[38372] = 25'b0000000110110000010111001;
    rom[38373] = 25'b0000000110110011110010100;
    rom[38374] = 25'b0000000110110111001101101;
    rom[38375] = 25'b0000000110111010101000110;
    rom[38376] = 25'b0000000110111110000011110;
    rom[38377] = 25'b0000000111000001011110100;
    rom[38378] = 25'b0000000111000100111001001;
    rom[38379] = 25'b0000000111001000010011101;
    rom[38380] = 25'b0000000111001011101110000;
    rom[38381] = 25'b0000000111001111001000001;
    rom[38382] = 25'b0000000111010010100010010;
    rom[38383] = 25'b0000000111010101111100001;
    rom[38384] = 25'b0000000111011001010101111;
    rom[38385] = 25'b0000000111011100101111100;
    rom[38386] = 25'b0000000111100000001000111;
    rom[38387] = 25'b0000000111100011100010010;
    rom[38388] = 25'b0000000111100110111011011;
    rom[38389] = 25'b0000000111101010010100010;
    rom[38390] = 25'b0000000111101101101101001;
    rom[38391] = 25'b0000000111110001000101111;
    rom[38392] = 25'b0000000111110100011110100;
    rom[38393] = 25'b0000000111110111110110111;
    rom[38394] = 25'b0000000111111011001111000;
    rom[38395] = 25'b0000000111111110100111001;
    rom[38396] = 25'b0000001000000001111111000;
    rom[38397] = 25'b0000001000000101010110111;
    rom[38398] = 25'b0000001000001000101110100;
    rom[38399] = 25'b0000001000001100000110000;
    rom[38400] = 25'b0000001000001111011101010;
    rom[38401] = 25'b0000001000010010110100100;
    rom[38402] = 25'b0000001000010110001011100;
    rom[38403] = 25'b0000001000011001100010011;
    rom[38404] = 25'b0000001000011100111001001;
    rom[38405] = 25'b0000001000100000001111101;
    rom[38406] = 25'b0000001000100011100110000;
    rom[38407] = 25'b0000001000100110111100010;
    rom[38408] = 25'b0000001000101010010010011;
    rom[38409] = 25'b0000001000101101101000011;
    rom[38410] = 25'b0000001000110000111110001;
    rom[38411] = 25'b0000001000110100010011101;
    rom[38412] = 25'b0000001000110111101001001;
    rom[38413] = 25'b0000001000111010111110100;
    rom[38414] = 25'b0000001000111110010011101;
    rom[38415] = 25'b0000001001000001101000101;
    rom[38416] = 25'b0000001001000100111101100;
    rom[38417] = 25'b0000001001001000010010001;
    rom[38418] = 25'b0000001001001011100110110;
    rom[38419] = 25'b0000001001001110111011001;
    rom[38420] = 25'b0000001001010010001111011;
    rom[38421] = 25'b0000001001010101100011011;
    rom[38422] = 25'b0000001001011000110111010;
    rom[38423] = 25'b0000001001011100001011000;
    rom[38424] = 25'b0000001001011111011110101;
    rom[38425] = 25'b0000001001100010110010001;
    rom[38426] = 25'b0000001001100110000101010;
    rom[38427] = 25'b0000001001101001011000100;
    rom[38428] = 25'b0000001001101100101011011;
    rom[38429] = 25'b0000001001101111111110010;
    rom[38430] = 25'b0000001001110011010000110;
    rom[38431] = 25'b0000001001110110100011010;
    rom[38432] = 25'b0000001001111001110101101;
    rom[38433] = 25'b0000001001111101000111110;
    rom[38434] = 25'b0000001010000000011001110;
    rom[38435] = 25'b0000001010000011101011101;
    rom[38436] = 25'b0000001010000110111101011;
    rom[38437] = 25'b0000001010001010001110110;
    rom[38438] = 25'b0000001010001101100000001;
    rom[38439] = 25'b0000001010010000110001011;
    rom[38440] = 25'b0000001010010100000010011;
    rom[38441] = 25'b0000001010010111010011010;
    rom[38442] = 25'b0000001010011010100100000;
    rom[38443] = 25'b0000001010011101110100100;
    rom[38444] = 25'b0000001010100001000100111;
    rom[38445] = 25'b0000001010100100010101001;
    rom[38446] = 25'b0000001010100111100101001;
    rom[38447] = 25'b0000001010101010110101000;
    rom[38448] = 25'b0000001010101110000100111;
    rom[38449] = 25'b0000001010110001010100011;
    rom[38450] = 25'b0000001010110100100011110;
    rom[38451] = 25'b0000001010110111110011000;
    rom[38452] = 25'b0000001010111011000010001;
    rom[38453] = 25'b0000001010111110010001000;
    rom[38454] = 25'b0000001011000001011111111;
    rom[38455] = 25'b0000001011000100101110011;
    rom[38456] = 25'b0000001011000111111100110;
    rom[38457] = 25'b0000001011001011001011001;
    rom[38458] = 25'b0000001011001110011001001;
    rom[38459] = 25'b0000001011010001100111001;
    rom[38460] = 25'b0000001011010100110100111;
    rom[38461] = 25'b0000001011011000000010100;
    rom[38462] = 25'b0000001011011011001111111;
    rom[38463] = 25'b0000001011011110011101001;
    rom[38464] = 25'b0000001011100001101010010;
    rom[38465] = 25'b0000001011100100110111010;
    rom[38466] = 25'b0000001011101000000100000;
    rom[38467] = 25'b0000001011101011010000100;
    rom[38468] = 25'b0000001011101110011101001;
    rom[38469] = 25'b0000001011110001101001010;
    rom[38470] = 25'b0000001011110100110101100;
    rom[38471] = 25'b0000001011111000000001011;
    rom[38472] = 25'b0000001011111011001101001;
    rom[38473] = 25'b0000001011111110011000110;
    rom[38474] = 25'b0000001100000001100100001;
    rom[38475] = 25'b0000001100000100101111100;
    rom[38476] = 25'b0000001100000111111010100;
    rom[38477] = 25'b0000001100001011000101011;
    rom[38478] = 25'b0000001100001110010000010;
    rom[38479] = 25'b0000001100010001011010110;
    rom[38480] = 25'b0000001100010100100101010;
    rom[38481] = 25'b0000001100010111101111100;
    rom[38482] = 25'b0000001100011010111001100;
    rom[38483] = 25'b0000001100011110000011100;
    rom[38484] = 25'b0000001100100001001101010;
    rom[38485] = 25'b0000001100100100010110111;
    rom[38486] = 25'b0000001100100111100000010;
    rom[38487] = 25'b0000001100101010101001100;
    rom[38488] = 25'b0000001100101101110010100;
    rom[38489] = 25'b0000001100110000111011100;
    rom[38490] = 25'b0000001100110100000100010;
    rom[38491] = 25'b0000001100110111001100110;
    rom[38492] = 25'b0000001100111010010101001;
    rom[38493] = 25'b0000001100111101011101011;
    rom[38494] = 25'b0000001101000000100101011;
    rom[38495] = 25'b0000001101000011101101010;
    rom[38496] = 25'b0000001101000110110101000;
    rom[38497] = 25'b0000001101001001111100100;
    rom[38498] = 25'b0000001101001101000011111;
    rom[38499] = 25'b0000001101010000001011000;
    rom[38500] = 25'b0000001101010011010010000;
    rom[38501] = 25'b0000001101010110011000111;
    rom[38502] = 25'b0000001101011001011111101;
    rom[38503] = 25'b0000001101011100100110000;
    rom[38504] = 25'b0000001101011111101100011;
    rom[38505] = 25'b0000001101100010110010100;
    rom[38506] = 25'b0000001101100101111000100;
    rom[38507] = 25'b0000001101101000111110010;
    rom[38508] = 25'b0000001101101100000011111;
    rom[38509] = 25'b0000001101101111001001011;
    rom[38510] = 25'b0000001101110010001110101;
    rom[38511] = 25'b0000001101110101010011110;
    rom[38512] = 25'b0000001101111000011000101;
    rom[38513] = 25'b0000001101111011011101011;
    rom[38514] = 25'b0000001101111110100010000;
    rom[38515] = 25'b0000001110000001100110011;
    rom[38516] = 25'b0000001110000100101010101;
    rom[38517] = 25'b0000001110000111101110110;
    rom[38518] = 25'b0000001110001010110010100;
    rom[38519] = 25'b0000001110001101110110010;
    rom[38520] = 25'b0000001110010000111001111;
    rom[38521] = 25'b0000001110010011111101001;
    rom[38522] = 25'b0000001110010111000000010;
    rom[38523] = 25'b0000001110011010000011010;
    rom[38524] = 25'b0000001110011101000110001;
    rom[38525] = 25'b0000001110100000001000110;
    rom[38526] = 25'b0000001110100011001011010;
    rom[38527] = 25'b0000001110100110001101101;
    rom[38528] = 25'b0000001110101001001111101;
    rom[38529] = 25'b0000001110101100010001101;
    rom[38530] = 25'b0000001110101111010011011;
    rom[38531] = 25'b0000001110110010010101000;
    rom[38532] = 25'b0000001110110101010110011;
    rom[38533] = 25'b0000001110111000010111101;
    rom[38534] = 25'b0000001110111011011000101;
    rom[38535] = 25'b0000001110111110011001100;
    rom[38536] = 25'b0000001111000001011010010;
    rom[38537] = 25'b0000001111000100011010101;
    rom[38538] = 25'b0000001111000111011011001;
    rom[38539] = 25'b0000001111001010011011001;
    rom[38540] = 25'b0000001111001101011011001;
    rom[38541] = 25'b0000001111010000011011000;
    rom[38542] = 25'b0000001111010011011010100;
    rom[38543] = 25'b0000001111010110011010000;
    rom[38544] = 25'b0000001111011001011001010;
    rom[38545] = 25'b0000001111011100011000010;
    rom[38546] = 25'b0000001111011111010111001;
    rom[38547] = 25'b0000001111100010010110000;
    rom[38548] = 25'b0000001111100101010100100;
    rom[38549] = 25'b0000001111101000010010110;
    rom[38550] = 25'b0000001111101011010001000;
    rom[38551] = 25'b0000001111101110001111000;
    rom[38552] = 25'b0000001111110001001100110;
    rom[38553] = 25'b0000001111110100001010011;
    rom[38554] = 25'b0000001111110111000111111;
    rom[38555] = 25'b0000001111111010000101001;
    rom[38556] = 25'b0000001111111101000010010;
    rom[38557] = 25'b0000001111111111111111001;
    rom[38558] = 25'b0000010000000010111011111;
    rom[38559] = 25'b0000010000000101111000010;
    rom[38560] = 25'b0000010000001000110100101;
    rom[38561] = 25'b0000010000001011110000111;
    rom[38562] = 25'b0000010000001110101100111;
    rom[38563] = 25'b0000010000010001101000101;
    rom[38564] = 25'b0000010000010100100100010;
    rom[38565] = 25'b0000010000010111011111110;
    rom[38566] = 25'b0000010000011010011011000;
    rom[38567] = 25'b0000010000011101010110001;
    rom[38568] = 25'b0000010000100000010000111;
    rom[38569] = 25'b0000010000100011001011101;
    rom[38570] = 25'b0000010000100110000110010;
    rom[38571] = 25'b0000010000101001000000100;
    rom[38572] = 25'b0000010000101011111010101;
    rom[38573] = 25'b0000010000101110110100101;
    rom[38574] = 25'b0000010000110001101110011;
    rom[38575] = 25'b0000010000110100101000000;
    rom[38576] = 25'b0000010000110111100001011;
    rom[38577] = 25'b0000010000111010011010101;
    rom[38578] = 25'b0000010000111101010011110;
    rom[38579] = 25'b0000010001000000001100100;
    rom[38580] = 25'b0000010001000011000101001;
    rom[38581] = 25'b0000010001000101111101101;
    rom[38582] = 25'b0000010001001000110101111;
    rom[38583] = 25'b0000010001001011101110001;
    rom[38584] = 25'b0000010001001110100110000;
    rom[38585] = 25'b0000010001010001011101110;
    rom[38586] = 25'b0000010001010100010101010;
    rom[38587] = 25'b0000010001010111001100101;
    rom[38588] = 25'b0000010001011010000011110;
    rom[38589] = 25'b0000010001011100111010111;
    rom[38590] = 25'b0000010001011111110001101;
    rom[38591] = 25'b0000010001100010101000010;
    rom[38592] = 25'b0000010001100101011110101;
    rom[38593] = 25'b0000010001101000010101000;
    rom[38594] = 25'b0000010001101011001011000;
    rom[38595] = 25'b0000010001101110000000111;
    rom[38596] = 25'b0000010001110000110110100;
    rom[38597] = 25'b0000010001110011101100000;
    rom[38598] = 25'b0000010001110110100001011;
    rom[38599] = 25'b0000010001111001010110011;
    rom[38600] = 25'b0000010001111100001011011;
    rom[38601] = 25'b0000010001111111000000001;
    rom[38602] = 25'b0000010010000001110100101;
    rom[38603] = 25'b0000010010000100101001000;
    rom[38604] = 25'b0000010010000111011101001;
    rom[38605] = 25'b0000010010001010010001001;
    rom[38606] = 25'b0000010010001101000100111;
    rom[38607] = 25'b0000010010001111111000101;
    rom[38608] = 25'b0000010010010010101100000;
    rom[38609] = 25'b0000010010010101011111001;
    rom[38610] = 25'b0000010010011000010010010;
    rom[38611] = 25'b0000010010011011000101000;
    rom[38612] = 25'b0000010010011101110111101;
    rom[38613] = 25'b0000010010100000101010001;
    rom[38614] = 25'b0000010010100011011100011;
    rom[38615] = 25'b0000010010100110001110100;
    rom[38616] = 25'b0000010010101001000000011;
    rom[38617] = 25'b0000010010101011110010000;
    rom[38618] = 25'b0000010010101110100011101;
    rom[38619] = 25'b0000010010110001010100111;
    rom[38620] = 25'b0000010010110100000110000;
    rom[38621] = 25'b0000010010110110110111000;
    rom[38622] = 25'b0000010010111001100111101;
    rom[38623] = 25'b0000010010111100011000010;
    rom[38624] = 25'b0000010010111111001000100;
    rom[38625] = 25'b0000010011000001111000110;
    rom[38626] = 25'b0000010011000100101000110;
    rom[38627] = 25'b0000010011000111011000100;
    rom[38628] = 25'b0000010011001010001000000;
    rom[38629] = 25'b0000010011001100110111011;
    rom[38630] = 25'b0000010011001111100110101;
    rom[38631] = 25'b0000010011010010010101101;
    rom[38632] = 25'b0000010011010101000100011;
    rom[38633] = 25'b0000010011010111110011000;
    rom[38634] = 25'b0000010011011010100001100;
    rom[38635] = 25'b0000010011011101001111110;
    rom[38636] = 25'b0000010011011111111101110;
    rom[38637] = 25'b0000010011100010101011101;
    rom[38638] = 25'b0000010011100101011001010;
    rom[38639] = 25'b0000010011101000000110110;
    rom[38640] = 25'b0000010011101010110100000;
    rom[38641] = 25'b0000010011101101100001000;
    rom[38642] = 25'b0000010011110000001101111;
    rom[38643] = 25'b0000010011110010111010101;
    rom[38644] = 25'b0000010011110101100111000;
    rom[38645] = 25'b0000010011111000010011011;
    rom[38646] = 25'b0000010011111010111111100;
    rom[38647] = 25'b0000010011111101101011011;
    rom[38648] = 25'b0000010100000000010111000;
    rom[38649] = 25'b0000010100000011000010101;
    rom[38650] = 25'b0000010100000101101101111;
    rom[38651] = 25'b0000010100001000011001000;
    rom[38652] = 25'b0000010100001011000011111;
    rom[38653] = 25'b0000010100001101101110101;
    rom[38654] = 25'b0000010100010000011001001;
    rom[38655] = 25'b0000010100010011000011100;
    rom[38656] = 25'b0000010100010101101101101;
    rom[38657] = 25'b0000010100011000010111100;
    rom[38658] = 25'b0000010100011011000001010;
    rom[38659] = 25'b0000010100011101101010110;
    rom[38660] = 25'b0000010100100000010100010;
    rom[38661] = 25'b0000010100100010111101011;
    rom[38662] = 25'b0000010100100101100110010;
    rom[38663] = 25'b0000010100101000001111000;
    rom[38664] = 25'b0000010100101010110111101;
    rom[38665] = 25'b0000010100101101100000000;
    rom[38666] = 25'b0000010100110000001000001;
    rom[38667] = 25'b0000010100110010110000000;
    rom[38668] = 25'b0000010100110101010111111;
    rom[38669] = 25'b0000010100110111111111011;
    rom[38670] = 25'b0000010100111010100110111;
    rom[38671] = 25'b0000010100111101001110000;
    rom[38672] = 25'b0000010100111111110101000;
    rom[38673] = 25'b0000010101000010011011110;
    rom[38674] = 25'b0000010101000101000010010;
    rom[38675] = 25'b0000010101000111101000110;
    rom[38676] = 25'b0000010101001010001110111;
    rom[38677] = 25'b0000010101001100110100111;
    rom[38678] = 25'b0000010101001111011010101;
    rom[38679] = 25'b0000010101010010000000010;
    rom[38680] = 25'b0000010101010100100101101;
    rom[38681] = 25'b0000010101010111001010110;
    rom[38682] = 25'b0000010101011001101111110;
    rom[38683] = 25'b0000010101011100010100100;
    rom[38684] = 25'b0000010101011110111001001;
    rom[38685] = 25'b0000010101100001011101100;
    rom[38686] = 25'b0000010101100100000001110;
    rom[38687] = 25'b0000010101100110100101110;
    rom[38688] = 25'b0000010101101001001001011;
    rom[38689] = 25'b0000010101101011101101000;
    rom[38690] = 25'b0000010101101110010000011;
    rom[38691] = 25'b0000010101110000110011101;
    rom[38692] = 25'b0000010101110011010110101;
    rom[38693] = 25'b0000010101110101111001011;
    rom[38694] = 25'b0000010101111000011100000;
    rom[38695] = 25'b0000010101111010111110011;
    rom[38696] = 25'b0000010101111101100000100;
    rom[38697] = 25'b0000010110000000000010100;
    rom[38698] = 25'b0000010110000010100100010;
    rom[38699] = 25'b0000010110000101000101110;
    rom[38700] = 25'b0000010110000111100111001;
    rom[38701] = 25'b0000010110001010001000011;
    rom[38702] = 25'b0000010110001100101001011;
    rom[38703] = 25'b0000010110001111001010001;
    rom[38704] = 25'b0000010110010001101010101;
    rom[38705] = 25'b0000010110010100001011000;
    rom[38706] = 25'b0000010110010110101011010;
    rom[38707] = 25'b0000010110011001001011001;
    rom[38708] = 25'b0000010110011011101010111;
    rom[38709] = 25'b0000010110011110001010011;
    rom[38710] = 25'b0000010110100000101001110;
    rom[38711] = 25'b0000010110100011001000111;
    rom[38712] = 25'b0000010110100101100111111;
    rom[38713] = 25'b0000010110101000000110101;
    rom[38714] = 25'b0000010110101010100101001;
    rom[38715] = 25'b0000010110101101000011011;
    rom[38716] = 25'b0000010110101111100001101;
    rom[38717] = 25'b0000010110110001111111100;
    rom[38718] = 25'b0000010110110100011101010;
    rom[38719] = 25'b0000010110110110111010101;
    rom[38720] = 25'b0000010110111001011000000;
    rom[38721] = 25'b0000010110111011110101001;
    rom[38722] = 25'b0000010110111110010010000;
    rom[38723] = 25'b0000010111000000101110110;
    rom[38724] = 25'b0000010111000011001011010;
    rom[38725] = 25'b0000010111000101100111100;
    rom[38726] = 25'b0000010111001000000011101;
    rom[38727] = 25'b0000010111001010011111100;
    rom[38728] = 25'b0000010111001100111011001;
    rom[38729] = 25'b0000010111001111010110101;
    rom[38730] = 25'b0000010111010001110001111;
    rom[38731] = 25'b0000010111010100001101000;
    rom[38732] = 25'b0000010111010110100111110;
    rom[38733] = 25'b0000010111011001000010100;
    rom[38734] = 25'b0000010111011011011100111;
    rom[38735] = 25'b0000010111011101110111001;
    rom[38736] = 25'b0000010111100000010001001;
    rom[38737] = 25'b0000010111100010101011000;
    rom[38738] = 25'b0000010111100101000100101;
    rom[38739] = 25'b0000010111100111011110000;
    rom[38740] = 25'b0000010111101001110111010;
    rom[38741] = 25'b0000010111101100010000001;
    rom[38742] = 25'b0000010111101110101001000;
    rom[38743] = 25'b0000010111110001000001100;
    rom[38744] = 25'b0000010111110011011010000;
    rom[38745] = 25'b0000010111110101110010001;
    rom[38746] = 25'b0000010111111000001010001;
    rom[38747] = 25'b0000010111111010100001111;
    rom[38748] = 25'b0000010111111100111001011;
    rom[38749] = 25'b0000010111111111010000110;
    rom[38750] = 25'b0000011000000001100111111;
    rom[38751] = 25'b0000011000000011111110111;
    rom[38752] = 25'b0000011000000110010101100;
    rom[38753] = 25'b0000011000001000101100001;
    rom[38754] = 25'b0000011000001011000010011;
    rom[38755] = 25'b0000011000001101011000100;
    rom[38756] = 25'b0000011000001111101110011;
    rom[38757] = 25'b0000011000010010000100001;
    rom[38758] = 25'b0000011000010100011001100;
    rom[38759] = 25'b0000011000010110101110111;
    rom[38760] = 25'b0000011000011001000011111;
    rom[38761] = 25'b0000011000011011011000110;
    rom[38762] = 25'b0000011000011101101101011;
    rom[38763] = 25'b0000011000100000000001111;
    rom[38764] = 25'b0000011000100010010110000;
    rom[38765] = 25'b0000011000100100101010000;
    rom[38766] = 25'b0000011000100110111101111;
    rom[38767] = 25'b0000011000101001010001011;
    rom[38768] = 25'b0000011000101011100100111;
    rom[38769] = 25'b0000011000101101111000000;
    rom[38770] = 25'b0000011000110000001011000;
    rom[38771] = 25'b0000011000110010011101110;
    rom[38772] = 25'b0000011000110100110000011;
    rom[38773] = 25'b0000011000110111000010110;
    rom[38774] = 25'b0000011000111001010100111;
    rom[38775] = 25'b0000011000111011100110110;
    rom[38776] = 25'b0000011000111101111000100;
    rom[38777] = 25'b0000011001000000001010000;
    rom[38778] = 25'b0000011001000010011011011;
    rom[38779] = 25'b0000011001000100101100011;
    rom[38780] = 25'b0000011001000110111101010;
    rom[38781] = 25'b0000011001001001001110000;
    rom[38782] = 25'b0000011001001011011110011;
    rom[38783] = 25'b0000011001001101101110101;
    rom[38784] = 25'b0000011001001111111110110;
    rom[38785] = 25'b0000011001010010001110100;
    rom[38786] = 25'b0000011001010100011110001;
    rom[38787] = 25'b0000011001010110101101100;
    rom[38788] = 25'b0000011001011000111100101;
    rom[38789] = 25'b0000011001011011001011110;
    rom[38790] = 25'b0000011001011101011010011;
    rom[38791] = 25'b0000011001011111101001000;
    rom[38792] = 25'b0000011001100001110111011;
    rom[38793] = 25'b0000011001100100000101100;
    rom[38794] = 25'b0000011001100110010011011;
    rom[38795] = 25'b0000011001101000100001010;
    rom[38796] = 25'b0000011001101010101110101;
    rom[38797] = 25'b0000011001101100111100000;
    rom[38798] = 25'b0000011001101111001001001;
    rom[38799] = 25'b0000011001110001010101111;
    rom[38800] = 25'b0000011001110011100010100;
    rom[38801] = 25'b0000011001110101101111000;
    rom[38802] = 25'b0000011001110111111011010;
    rom[38803] = 25'b0000011001111010000111010;
    rom[38804] = 25'b0000011001111100010011000;
    rom[38805] = 25'b0000011001111110011110101;
    rom[38806] = 25'b0000011010000000101010001;
    rom[38807] = 25'b0000011010000010110101010;
    rom[38808] = 25'b0000011010000101000000010;
    rom[38809] = 25'b0000011010000111001011000;
    rom[38810] = 25'b0000011010001001010101100;
    rom[38811] = 25'b0000011010001011011111111;
    rom[38812] = 25'b0000011010001101101001111;
    rom[38813] = 25'b0000011010001111110011111;
    rom[38814] = 25'b0000011010010001111101100;
    rom[38815] = 25'b0000011010010100000111000;
    rom[38816] = 25'b0000011010010110010000010;
    rom[38817] = 25'b0000011010011000011001010;
    rom[38818] = 25'b0000011010011010100010001;
    rom[38819] = 25'b0000011010011100101010110;
    rom[38820] = 25'b0000011010011110110011001;
    rom[38821] = 25'b0000011010100000111011011;
    rom[38822] = 25'b0000011010100011000011011;
    rom[38823] = 25'b0000011010100101001011001;
    rom[38824] = 25'b0000011010100111010010101;
    rom[38825] = 25'b0000011010101001011010000;
    rom[38826] = 25'b0000011010101011100001001;
    rom[38827] = 25'b0000011010101101101000000;
    rom[38828] = 25'b0000011010101111101110110;
    rom[38829] = 25'b0000011010110001110101010;
    rom[38830] = 25'b0000011010110011111011011;
    rom[38831] = 25'b0000011010110110000001100;
    rom[38832] = 25'b0000011010111000000111011;
    rom[38833] = 25'b0000011010111010001101000;
    rom[38834] = 25'b0000011010111100010010011;
    rom[38835] = 25'b0000011010111110010111101;
    rom[38836] = 25'b0000011011000000011100101;
    rom[38837] = 25'b0000011011000010100001010;
    rom[38838] = 25'b0000011011000100100101111;
    rom[38839] = 25'b0000011011000110101010010;
    rom[38840] = 25'b0000011011001000101110011;
    rom[38841] = 25'b0000011011001010110010010;
    rom[38842] = 25'b0000011011001100110101111;
    rom[38843] = 25'b0000011011001110111001011;
    rom[38844] = 25'b0000011011010000111100110;
    rom[38845] = 25'b0000011011010010111111110;
    rom[38846] = 25'b0000011011010101000010101;
    rom[38847] = 25'b0000011011010111000101010;
    rom[38848] = 25'b0000011011011001000111101;
    rom[38849] = 25'b0000011011011011001001110;
    rom[38850] = 25'b0000011011011101001011110;
    rom[38851] = 25'b0000011011011111001101100;
    rom[38852] = 25'b0000011011100001001111000;
    rom[38853] = 25'b0000011011100011010000011;
    rom[38854] = 25'b0000011011100101010001100;
    rom[38855] = 25'b0000011011100111010010011;
    rom[38856] = 25'b0000011011101001010011000;
    rom[38857] = 25'b0000011011101011010011100;
    rom[38858] = 25'b0000011011101101010011101;
    rom[38859] = 25'b0000011011101111010011110;
    rom[38860] = 25'b0000011011110001010011101;
    rom[38861] = 25'b0000011011110011010011001;
    rom[38862] = 25'b0000011011110101010010100;
    rom[38863] = 25'b0000011011110111010001110;
    rom[38864] = 25'b0000011011111001010000101;
    rom[38865] = 25'b0000011011111011001111011;
    rom[38866] = 25'b0000011011111101001101111;
    rom[38867] = 25'b0000011011111111001100001;
    rom[38868] = 25'b0000011100000001001010010;
    rom[38869] = 25'b0000011100000011001000001;
    rom[38870] = 25'b0000011100000101000101110;
    rom[38871] = 25'b0000011100000111000011010;
    rom[38872] = 25'b0000011100001001000000011;
    rom[38873] = 25'b0000011100001010111101011;
    rom[38874] = 25'b0000011100001100111010001;
    rom[38875] = 25'b0000011100001110110110110;
    rom[38876] = 25'b0000011100010000110011000;
    rom[38877] = 25'b0000011100010010101111001;
    rom[38878] = 25'b0000011100010100101011001;
    rom[38879] = 25'b0000011100010110100110111;
    rom[38880] = 25'b0000011100011000100010010;
    rom[38881] = 25'b0000011100011010011101100;
    rom[38882] = 25'b0000011100011100011000100;
    rom[38883] = 25'b0000011100011110010011011;
    rom[38884] = 25'b0000011100100000001110000;
    rom[38885] = 25'b0000011100100010001000010;
    rom[38886] = 25'b0000011100100100000010100;
    rom[38887] = 25'b0000011100100101111100011;
    rom[38888] = 25'b0000011100100111110110010;
    rom[38889] = 25'b0000011100101001101111101;
    rom[38890] = 25'b0000011100101011101001000;
    rom[38891] = 25'b0000011100101101100010000;
    rom[38892] = 25'b0000011100101111011010111;
    rom[38893] = 25'b0000011100110001010011100;
    rom[38894] = 25'b0000011100110011001100000;
    rom[38895] = 25'b0000011100110101000100001;
    rom[38896] = 25'b0000011100110110111100001;
    rom[38897] = 25'b0000011100111000110011111;
    rom[38898] = 25'b0000011100111010101011100;
    rom[38899] = 25'b0000011100111100100010110;
    rom[38900] = 25'b0000011100111110011001111;
    rom[38901] = 25'b0000011101000000010000111;
    rom[38902] = 25'b0000011101000010000111011;
    rom[38903] = 25'b0000011101000011111110000;
    rom[38904] = 25'b0000011101000101110100001;
    rom[38905] = 25'b0000011101000111101010001;
    rom[38906] = 25'b0000011101001001100000000;
    rom[38907] = 25'b0000011101001011010101100;
    rom[38908] = 25'b0000011101001101001010111;
    rom[38909] = 25'b0000011101001111000000000;
    rom[38910] = 25'b0000011101010000110101000;
    rom[38911] = 25'b0000011101010010101001101;
    rom[38912] = 25'b0000011101010100011110001;
    rom[38913] = 25'b0000011101010110010010011;
    rom[38914] = 25'b0000011101011000000110011;
    rom[38915] = 25'b0000011101011001111010010;
    rom[38916] = 25'b0000011101011011101101111;
    rom[38917] = 25'b0000011101011101100001010;
    rom[38918] = 25'b0000011101011111010100011;
    rom[38919] = 25'b0000011101100001000111011;
    rom[38920] = 25'b0000011101100010111010001;
    rom[38921] = 25'b0000011101100100101100101;
    rom[38922] = 25'b0000011101100110011110111;
    rom[38923] = 25'b0000011101101000010001000;
    rom[38924] = 25'b0000011101101010000010110;
    rom[38925] = 25'b0000011101101011110100011;
    rom[38926] = 25'b0000011101101101100101110;
    rom[38927] = 25'b0000011101101111010111000;
    rom[38928] = 25'b0000011101110001001000000;
    rom[38929] = 25'b0000011101110010111000110;
    rom[38930] = 25'b0000011101110100101001010;
    rom[38931] = 25'b0000011101110110011001101;
    rom[38932] = 25'b0000011101111000001001101;
    rom[38933] = 25'b0000011101111001111001100;
    rom[38934] = 25'b0000011101111011101001001;
    rom[38935] = 25'b0000011101111101011000100;
    rom[38936] = 25'b0000011101111111000111110;
    rom[38937] = 25'b0000011110000000110110110;
    rom[38938] = 25'b0000011110000010100101100;
    rom[38939] = 25'b0000011110000100010100000;
    rom[38940] = 25'b0000011110000110000010011;
    rom[38941] = 25'b0000011110000111110000100;
    rom[38942] = 25'b0000011110001001011110011;
    rom[38943] = 25'b0000011110001011001100001;
    rom[38944] = 25'b0000011110001100111001011;
    rom[38945] = 25'b0000011110001110100110110;
    rom[38946] = 25'b0000011110010000010011101;
    rom[38947] = 25'b0000011110010010000000100;
    rom[38948] = 25'b0000011110010011101101000;
    rom[38949] = 25'b0000011110010101011001010;
    rom[38950] = 25'b0000011110010111000101100;
    rom[38951] = 25'b0000011110011000110001011;
    rom[38952] = 25'b0000011110011010011101000;
    rom[38953] = 25'b0000011110011100001000100;
    rom[38954] = 25'b0000011110011101110011110;
    rom[38955] = 25'b0000011110011111011110110;
    rom[38956] = 25'b0000011110100001001001100;
    rom[38957] = 25'b0000011110100010110100001;
    rom[38958] = 25'b0000011110100100011110100;
    rom[38959] = 25'b0000011110100110001000100;
    rom[38960] = 25'b0000011110100111110010100;
    rom[38961] = 25'b0000011110101001011100001;
    rom[38962] = 25'b0000011110101011000101101;
    rom[38963] = 25'b0000011110101100101110111;
    rom[38964] = 25'b0000011110101110010111111;
    rom[38965] = 25'b0000011110110000000000110;
    rom[38966] = 25'b0000011110110001101001010;
    rom[38967] = 25'b0000011110110011010001101;
    rom[38968] = 25'b0000011110110100111001110;
    rom[38969] = 25'b0000011110110110100001101;
    rom[38970] = 25'b0000011110111000001001011;
    rom[38971] = 25'b0000011110111001110000110;
    rom[38972] = 25'b0000011110111011011000000;
    rom[38973] = 25'b0000011110111100111111001;
    rom[38974] = 25'b0000011110111110100101111;
    rom[38975] = 25'b0000011111000000001100100;
    rom[38976] = 25'b0000011111000001110010110;
    rom[38977] = 25'b0000011111000011011001000;
    rom[38978] = 25'b0000011111000100111110111;
    rom[38979] = 25'b0000011111000110100100100;
    rom[38980] = 25'b0000011111001000001010000;
    rom[38981] = 25'b0000011111001001101111010;
    rom[38982] = 25'b0000011111001011010100011;
    rom[38983] = 25'b0000011111001100111001001;
    rom[38984] = 25'b0000011111001110011101101;
    rom[38985] = 25'b0000011111010000000010001;
    rom[38986] = 25'b0000011111010001100110001;
    rom[38987] = 25'b0000011111010011001010001;
    rom[38988] = 25'b0000011111010100101101110;
    rom[38989] = 25'b0000011111010110010001010;
    rom[38990] = 25'b0000011111010111110100100;
    rom[38991] = 25'b0000011111011001010111100;
    rom[38992] = 25'b0000011111011010111010011;
    rom[38993] = 25'b0000011111011100011101000;
    rom[38994] = 25'b0000011111011101111111011;
    rom[38995] = 25'b0000011111011111100001100;
    rom[38996] = 25'b0000011111100001000011011;
    rom[38997] = 25'b0000011111100010100101000;
    rom[38998] = 25'b0000011111100100000110100;
    rom[38999] = 25'b0000011111100101100111110;
    rom[39000] = 25'b0000011111100111001000110;
    rom[39001] = 25'b0000011111101000101001101;
    rom[39002] = 25'b0000011111101010001010001;
    rom[39003] = 25'b0000011111101011101010100;
    rom[39004] = 25'b0000011111101101001010101;
    rom[39005] = 25'b0000011111101110101010101;
    rom[39006] = 25'b0000011111110000001010010;
    rom[39007] = 25'b0000011111110001101001110;
    rom[39008] = 25'b0000011111110011001001000;
    rom[39009] = 25'b0000011111110100101000000;
    rom[39010] = 25'b0000011111110110000110111;
    rom[39011] = 25'b0000011111110111100101011;
    rom[39012] = 25'b0000011111111001000011110;
    rom[39013] = 25'b0000011111111010100001111;
    rom[39014] = 25'b0000011111111011111111111;
    rom[39015] = 25'b0000011111111101011101100;
    rom[39016] = 25'b0000011111111110111011000;
    rom[39017] = 25'b0000100000000000011000001;
    rom[39018] = 25'b0000100000000001110101001;
    rom[39019] = 25'b0000100000000011010010000;
    rom[39020] = 25'b0000100000000100101110100;
    rom[39021] = 25'b0000100000000110001010111;
    rom[39022] = 25'b0000100000000111100111001;
    rom[39023] = 25'b0000100000001001000011000;
    rom[39024] = 25'b0000100000001010011110101;
    rom[39025] = 25'b0000100000001011111010001;
    rom[39026] = 25'b0000100000001101010101011;
    rom[39027] = 25'b0000100000001110110000011;
    rom[39028] = 25'b0000100000010000001011001;
    rom[39029] = 25'b0000100000010001100101110;
    rom[39030] = 25'b0000100000010011000000001;
    rom[39031] = 25'b0000100000010100011010001;
    rom[39032] = 25'b0000100000010101110100001;
    rom[39033] = 25'b0000100000010111001101110;
    rom[39034] = 25'b0000100000011000100111010;
    rom[39035] = 25'b0000100000011010000000011;
    rom[39036] = 25'b0000100000011011011001100;
    rom[39037] = 25'b0000100000011100110010010;
    rom[39038] = 25'b0000100000011110001010111;
    rom[39039] = 25'b0000100000011111100011001;
    rom[39040] = 25'b0000100000100000111011010;
    rom[39041] = 25'b0000100000100010010011001;
    rom[39042] = 25'b0000100000100011101010111;
    rom[39043] = 25'b0000100000100101000010010;
    rom[39044] = 25'b0000100000100110011001100;
    rom[39045] = 25'b0000100000100111110000100;
    rom[39046] = 25'b0000100000101001000111010;
    rom[39047] = 25'b0000100000101010011101111;
    rom[39048] = 25'b0000100000101011110100001;
    rom[39049] = 25'b0000100000101101001010010;
    rom[39050] = 25'b0000100000101110100000001;
    rom[39051] = 25'b0000100000101111110101110;
    rom[39052] = 25'b0000100000110001001011010;
    rom[39053] = 25'b0000100000110010100000100;
    rom[39054] = 25'b0000100000110011110101100;
    rom[39055] = 25'b0000100000110101001010001;
    rom[39056] = 25'b0000100000110110011110110;
    rom[39057] = 25'b0000100000110111110011001;
    rom[39058] = 25'b0000100000111001000111001;
    rom[39059] = 25'b0000100000111010011011000;
    rom[39060] = 25'b0000100000111011101110101;
    rom[39061] = 25'b0000100000111101000010001;
    rom[39062] = 25'b0000100000111110010101010;
    rom[39063] = 25'b0000100000111111101000010;
    rom[39064] = 25'b0000100001000000111011000;
    rom[39065] = 25'b0000100001000010001101101;
    rom[39066] = 25'b0000100001000011011111111;
    rom[39067] = 25'b0000100001000100110010000;
    rom[39068] = 25'b0000100001000110000011111;
    rom[39069] = 25'b0000100001000111010101100;
    rom[39070] = 25'b0000100001001000100110111;
    rom[39071] = 25'b0000100001001001111000001;
    rom[39072] = 25'b0000100001001011001001000;
    rom[39073] = 25'b0000100001001100011001111;
    rom[39074] = 25'b0000100001001101101010011;
    rom[39075] = 25'b0000100001001110111010101;
    rom[39076] = 25'b0000100001010000001010110;
    rom[39077] = 25'b0000100001010001011010101;
    rom[39078] = 25'b0000100001010010101010001;
    rom[39079] = 25'b0000100001010011111001101;
    rom[39080] = 25'b0000100001010101001000111;
    rom[39081] = 25'b0000100001010110010111110;
    rom[39082] = 25'b0000100001010111100110100;
    rom[39083] = 25'b0000100001011000110101000;
    rom[39084] = 25'b0000100001011010000011010;
    rom[39085] = 25'b0000100001011011010001011;
    rom[39086] = 25'b0000100001011100011111010;
    rom[39087] = 25'b0000100001011101101100111;
    rom[39088] = 25'b0000100001011110111010010;
    rom[39089] = 25'b0000100001100000000111011;
    rom[39090] = 25'b0000100001100001010100011;
    rom[39091] = 25'b0000100001100010100001001;
    rom[39092] = 25'b0000100001100011101101101;
    rom[39093] = 25'b0000100001100100111001111;
    rom[39094] = 25'b0000100001100110000101111;
    rom[39095] = 25'b0000100001100111010001111;
    rom[39096] = 25'b0000100001101000011101011;
    rom[39097] = 25'b0000100001101001101000110;
    rom[39098] = 25'b0000100001101010110011111;
    rom[39099] = 25'b0000100001101011111110111;
    rom[39100] = 25'b0000100001101101001001101;
    rom[39101] = 25'b0000100001101110010100001;
    rom[39102] = 25'b0000100001101111011110011;
    rom[39103] = 25'b0000100001110000101000011;
    rom[39104] = 25'b0000100001110001110010010;
    rom[39105] = 25'b0000100001110010111011111;
    rom[39106] = 25'b0000100001110100000101010;
    rom[39107] = 25'b0000100001110101001110011;
    rom[39108] = 25'b0000100001110110010111011;
    rom[39109] = 25'b0000100001110111100000000;
    rom[39110] = 25'b0000100001111000101000101;
    rom[39111] = 25'b0000100001111001110000110;
    rom[39112] = 25'b0000100001111010111000111;
    rom[39113] = 25'b0000100001111100000000101;
    rom[39114] = 25'b0000100001111101001000010;
    rom[39115] = 25'b0000100001111110001111101;
    rom[39116] = 25'b0000100001111111010110110;
    rom[39117] = 25'b0000100010000000011101101;
    rom[39118] = 25'b0000100010000001100100011;
    rom[39119] = 25'b0000100010000010101010111;
    rom[39120] = 25'b0000100010000011110001001;
    rom[39121] = 25'b0000100010000100110111001;
    rom[39122] = 25'b0000100010000101111101000;
    rom[39123] = 25'b0000100010000111000010101;
    rom[39124] = 25'b0000100010001000001000000;
    rom[39125] = 25'b0000100010001001001101001;
    rom[39126] = 25'b0000100010001010010010000;
    rom[39127] = 25'b0000100010001011010110101;
    rom[39128] = 25'b0000100010001100011011001;
    rom[39129] = 25'b0000100010001101011111011;
    rom[39130] = 25'b0000100010001110100011011;
    rom[39131] = 25'b0000100010001111100111010;
    rom[39132] = 25'b0000100010010000101010111;
    rom[39133] = 25'b0000100010010001101110001;
    rom[39134] = 25'b0000100010010010110001011;
    rom[39135] = 25'b0000100010010011110100001;
    rom[39136] = 25'b0000100010010100110110111;
    rom[39137] = 25'b0000100010010101111001011;
    rom[39138] = 25'b0000100010010110111011101;
    rom[39139] = 25'b0000100010010111111101101;
    rom[39140] = 25'b0000100010011000111111011;
    rom[39141] = 25'b0000100010011010000001000;
    rom[39142] = 25'b0000100010011011000010011;
    rom[39143] = 25'b0000100010011100000011100;
    rom[39144] = 25'b0000100010011101000100100;
    rom[39145] = 25'b0000100010011110000101001;
    rom[39146] = 25'b0000100010011111000101100;
    rom[39147] = 25'b0000100010100000000101110;
    rom[39148] = 25'b0000100010100001000101111;
    rom[39149] = 25'b0000100010100010000101101;
    rom[39150] = 25'b0000100010100011000101010;
    rom[39151] = 25'b0000100010100100000100100;
    rom[39152] = 25'b0000100010100101000011101;
    rom[39153] = 25'b0000100010100110000010101;
    rom[39154] = 25'b0000100010100111000001010;
    rom[39155] = 25'b0000100010100111111111110;
    rom[39156] = 25'b0000100010101000111101111;
    rom[39157] = 25'b0000100010101001111011111;
    rom[39158] = 25'b0000100010101010111001110;
    rom[39159] = 25'b0000100010101011110111010;
    rom[39160] = 25'b0000100010101100110100101;
    rom[39161] = 25'b0000100010101101110001111;
    rom[39162] = 25'b0000100010101110101110110;
    rom[39163] = 25'b0000100010101111101011011;
    rom[39164] = 25'b0000100010110000100111111;
    rom[39165] = 25'b0000100010110001100100000;
    rom[39166] = 25'b0000100010110010100000001;
    rom[39167] = 25'b0000100010110011011011111;
    rom[39168] = 25'b0000100010110100010111100;
    rom[39169] = 25'b0000100010110101010010110;
    rom[39170] = 25'b0000100010110110001101111;
    rom[39171] = 25'b0000100010110111001000110;
    rom[39172] = 25'b0000100010111000000011100;
    rom[39173] = 25'b0000100010111000111110000;
    rom[39174] = 25'b0000100010111001111000001;
    rom[39175] = 25'b0000100010111010110010001;
    rom[39176] = 25'b0000100010111011101100000;
    rom[39177] = 25'b0000100010111100100101101;
    rom[39178] = 25'b0000100010111101011111000;
    rom[39179] = 25'b0000100010111110011000001;
    rom[39180] = 25'b0000100010111111010001000;
    rom[39181] = 25'b0000100011000000001001101;
    rom[39182] = 25'b0000100011000001000010001;
    rom[39183] = 25'b0000100011000001111010011;
    rom[39184] = 25'b0000100011000010110010011;
    rom[39185] = 25'b0000100011000011101010001;
    rom[39186] = 25'b0000100011000100100001110;
    rom[39187] = 25'b0000100011000101011001001;
    rom[39188] = 25'b0000100011000110010000010;
    rom[39189] = 25'b0000100011000111000111001;
    rom[39190] = 25'b0000100011000111111101111;
    rom[39191] = 25'b0000100011001000110100010;
    rom[39192] = 25'b0000100011001001101010100;
    rom[39193] = 25'b0000100011001010100000101;
    rom[39194] = 25'b0000100011001011010110011;
    rom[39195] = 25'b0000100011001100001100000;
    rom[39196] = 25'b0000100011001101000001011;
    rom[39197] = 25'b0000100011001101110110100;
    rom[39198] = 25'b0000100011001110101011011;
    rom[39199] = 25'b0000100011001111100000001;
    rom[39200] = 25'b0000100011010000010100101;
    rom[39201] = 25'b0000100011010001001000111;
    rom[39202] = 25'b0000100011010001111100111;
    rom[39203] = 25'b0000100011010010110000110;
    rom[39204] = 25'b0000100011010011100100010;
    rom[39205] = 25'b0000100011010100010111101;
    rom[39206] = 25'b0000100011010101001010110;
    rom[39207] = 25'b0000100011010101111101110;
    rom[39208] = 25'b0000100011010110110000011;
    rom[39209] = 25'b0000100011010111100010111;
    rom[39210] = 25'b0000100011011000010101001;
    rom[39211] = 25'b0000100011011001000111010;
    rom[39212] = 25'b0000100011011001111001001;
    rom[39213] = 25'b0000100011011010101010101;
    rom[39214] = 25'b0000100011011011011100001;
    rom[39215] = 25'b0000100011011100001101010;
    rom[39216] = 25'b0000100011011100111110001;
    rom[39217] = 25'b0000100011011101101110111;
    rom[39218] = 25'b0000100011011110011111011;
    rom[39219] = 25'b0000100011011111001111101;
    rom[39220] = 25'b0000100011011111111111110;
    rom[39221] = 25'b0000100011100000101111100;
    rom[39222] = 25'b0000100011100001011111001;
    rom[39223] = 25'b0000100011100010001110101;
    rom[39224] = 25'b0000100011100010111101110;
    rom[39225] = 25'b0000100011100011101100110;
    rom[39226] = 25'b0000100011100100011011100;
    rom[39227] = 25'b0000100011100101001010000;
    rom[39228] = 25'b0000100011100101111000010;
    rom[39229] = 25'b0000100011100110100110011;
    rom[39230] = 25'b0000100011100111010100010;
    rom[39231] = 25'b0000100011101000000001111;
    rom[39232] = 25'b0000100011101000101111010;
    rom[39233] = 25'b0000100011101001011100100;
    rom[39234] = 25'b0000100011101010001001100;
    rom[39235] = 25'b0000100011101010110110010;
    rom[39236] = 25'b0000100011101011100010110;
    rom[39237] = 25'b0000100011101100001111001;
    rom[39238] = 25'b0000100011101100111011010;
    rom[39239] = 25'b0000100011101101100111001;
    rom[39240] = 25'b0000100011101110010010110;
    rom[39241] = 25'b0000100011101110111110001;
    rom[39242] = 25'b0000100011101111101001011;
    rom[39243] = 25'b0000100011110000010100100;
    rom[39244] = 25'b0000100011110000111111010;
    rom[39245] = 25'b0000100011110001101001110;
    rom[39246] = 25'b0000100011110010010100001;
    rom[39247] = 25'b0000100011110010111110010;
    rom[39248] = 25'b0000100011110011101000001;
    rom[39249] = 25'b0000100011110100010001110;
    rom[39250] = 25'b0000100011110100111011011;
    rom[39251] = 25'b0000100011110101100100100;
    rom[39252] = 25'b0000100011110110001101101;
    rom[39253] = 25'b0000100011110110110110100;
    rom[39254] = 25'b0000100011110111011111000;
    rom[39255] = 25'b0000100011111000000111011;
    rom[39256] = 25'b0000100011111000101111101;
    rom[39257] = 25'b0000100011111001010111100;
    rom[39258] = 25'b0000100011111001111111010;
    rom[39259] = 25'b0000100011111010100110110;
    rom[39260] = 25'b0000100011111011001110000;
    rom[39261] = 25'b0000100011111011110101001;
    rom[39262] = 25'b0000100011111100011011111;
    rom[39263] = 25'b0000100011111101000010100;
    rom[39264] = 25'b0000100011111101101000111;
    rom[39265] = 25'b0000100011111110001111001;
    rom[39266] = 25'b0000100011111110110101001;
    rom[39267] = 25'b0000100011111111011010111;
    rom[39268] = 25'b0000100100000000000000011;
    rom[39269] = 25'b0000100100000000100101110;
    rom[39270] = 25'b0000100100000001001010110;
    rom[39271] = 25'b0000100100000001101111101;
    rom[39272] = 25'b0000100100000010010100011;
    rom[39273] = 25'b0000100100000010111000110;
    rom[39274] = 25'b0000100100000011011101000;
    rom[39275] = 25'b0000100100000100000001000;
    rom[39276] = 25'b0000100100000100100100111;
    rom[39277] = 25'b0000100100000101001000011;
    rom[39278] = 25'b0000100100000101101011110;
    rom[39279] = 25'b0000100100000110001110111;
    rom[39280] = 25'b0000100100000110110001110;
    rom[39281] = 25'b0000100100000111010100100;
    rom[39282] = 25'b0000100100000111110111000;
    rom[39283] = 25'b0000100100001000011001010;
    rom[39284] = 25'b0000100100001000111011011;
    rom[39285] = 25'b0000100100001001011101001;
    rom[39286] = 25'b0000100100001001111110110;
    rom[39287] = 25'b0000100100001010100000001;
    rom[39288] = 25'b0000100100001011000001011;
    rom[39289] = 25'b0000100100001011100010010;
    rom[39290] = 25'b0000100100001100000011001;
    rom[39291] = 25'b0000100100001100100011101;
    rom[39292] = 25'b0000100100001101000011111;
    rom[39293] = 25'b0000100100001101100100000;
    rom[39294] = 25'b0000100100001110000011111;
    rom[39295] = 25'b0000100100001110100011100;
    rom[39296] = 25'b0000100100001111000011000;
    rom[39297] = 25'b0000100100001111100010010;
    rom[39298] = 25'b0000100100010000000001010;
    rom[39299] = 25'b0000100100010000100000000;
    rom[39300] = 25'b0000100100010000111110101;
    rom[39301] = 25'b0000100100010001011101000;
    rom[39302] = 25'b0000100100010001111011001;
    rom[39303] = 25'b0000100100010010011001001;
    rom[39304] = 25'b0000100100010010110110111;
    rom[39305] = 25'b0000100100010011010100011;
    rom[39306] = 25'b0000100100010011110001101;
    rom[39307] = 25'b0000100100010100001110110;
    rom[39308] = 25'b0000100100010100101011100;
    rom[39309] = 25'b0000100100010101001000001;
    rom[39310] = 25'b0000100100010101100100101;
    rom[39311] = 25'b0000100100010110000000111;
    rom[39312] = 25'b0000100100010110011100110;
    rom[39313] = 25'b0000100100010110111000101;
    rom[39314] = 25'b0000100100010111010100001;
    rom[39315] = 25'b0000100100010111101111100;
    rom[39316] = 25'b0000100100011000001010101;
    rom[39317] = 25'b0000100100011000100101100;
    rom[39318] = 25'b0000100100011001000000001;
    rom[39319] = 25'b0000100100011001011010110;
    rom[39320] = 25'b0000100100011001110100111;
    rom[39321] = 25'b0000100100011010001111000;
    rom[39322] = 25'b0000100100011010101000111;
    rom[39323] = 25'b0000100100011011000010100;
    rom[39324] = 25'b0000100100011011011011111;
    rom[39325] = 25'b0000100100011011110101001;
    rom[39326] = 25'b0000100100011100001110001;
    rom[39327] = 25'b0000100100011100100110111;
    rom[39328] = 25'b0000100100011100111111011;
    rom[39329] = 25'b0000100100011101010111101;
    rom[39330] = 25'b0000100100011101101111111;
    rom[39331] = 25'b0000100100011110000111110;
    rom[39332] = 25'b0000100100011110011111011;
    rom[39333] = 25'b0000100100011110110110111;
    rom[39334] = 25'b0000100100011111001110010;
    rom[39335] = 25'b0000100100011111100101010;
    rom[39336] = 25'b0000100100011111111100000;
    rom[39337] = 25'b0000100100100000010010110;
    rom[39338] = 25'b0000100100100000101001001;
    rom[39339] = 25'b0000100100100000111111010;
    rom[39340] = 25'b0000100100100001010101011;
    rom[39341] = 25'b0000100100100001101011001;
    rom[39342] = 25'b0000100100100010000000101;
    rom[39343] = 25'b0000100100100010010110000;
    rom[39344] = 25'b0000100100100010101011000;
    rom[39345] = 25'b0000100100100011000000000;
    rom[39346] = 25'b0000100100100011010100110;
    rom[39347] = 25'b0000100100100011101001001;
    rom[39348] = 25'b0000100100100011111101011;
    rom[39349] = 25'b0000100100100100010001100;
    rom[39350] = 25'b0000100100100100100101011;
    rom[39351] = 25'b0000100100100100111001000;
    rom[39352] = 25'b0000100100100101001100011;
    rom[39353] = 25'b0000100100100101011111101;
    rom[39354] = 25'b0000100100100101110010101;
    rom[39355] = 25'b0000100100100110000101011;
    rom[39356] = 25'b0000100100100110011000000;
    rom[39357] = 25'b0000100100100110101010011;
    rom[39358] = 25'b0000100100100110111100100;
    rom[39359] = 25'b0000100100100111001110011;
    rom[39360] = 25'b0000100100100111100000001;
    rom[39361] = 25'b0000100100100111110001101;
    rom[39362] = 25'b0000100100101000000011000;
    rom[39363] = 25'b0000100100101000010100001;
    rom[39364] = 25'b0000100100101000100100111;
    rom[39365] = 25'b0000100100101000110101101;
    rom[39366] = 25'b0000100100101001000110000;
    rom[39367] = 25'b0000100100101001010110010;
    rom[39368] = 25'b0000100100101001100110011;
    rom[39369] = 25'b0000100100101001110110001;
    rom[39370] = 25'b0000100100101010000101110;
    rom[39371] = 25'b0000100100101010010101001;
    rom[39372] = 25'b0000100100101010100100010;
    rom[39373] = 25'b0000100100101010110011010;
    rom[39374] = 25'b0000100100101011000010000;
    rom[39375] = 25'b0000100100101011010000101;
    rom[39376] = 25'b0000100100101011011110111;
    rom[39377] = 25'b0000100100101011101101000;
    rom[39378] = 25'b0000100100101011111010111;
    rom[39379] = 25'b0000100100101100001000101;
    rom[39380] = 25'b0000100100101100010110010;
    rom[39381] = 25'b0000100100101100100011100;
    rom[39382] = 25'b0000100100101100110000100;
    rom[39383] = 25'b0000100100101100111101011;
    rom[39384] = 25'b0000100100101101001010000;
    rom[39385] = 25'b0000100100101101010110100;
    rom[39386] = 25'b0000100100101101100010110;
    rom[39387] = 25'b0000100100101101101110110;
    rom[39388] = 25'b0000100100101101111010101;
    rom[39389] = 25'b0000100100101110000110001;
    rom[39390] = 25'b0000100100101110010001101;
    rom[39391] = 25'b0000100100101110011100110;
    rom[39392] = 25'b0000100100101110100111110;
    rom[39393] = 25'b0000100100101110110010100;
    rom[39394] = 25'b0000100100101110111101000;
    rom[39395] = 25'b0000100100101111000111011;
    rom[39396] = 25'b0000100100101111010001100;
    rom[39397] = 25'b0000100100101111011011011;
    rom[39398] = 25'b0000100100101111100101001;
    rom[39399] = 25'b0000100100101111101110101;
    rom[39400] = 25'b0000100100101111110111111;
    rom[39401] = 25'b0000100100110000000001001;
    rom[39402] = 25'b0000100100110000001010000;
    rom[39403] = 25'b0000100100110000010010101;
    rom[39404] = 25'b0000100100110000011011000;
    rom[39405] = 25'b0000100100110000100011011;
    rom[39406] = 25'b0000100100110000101011011;
    rom[39407] = 25'b0000100100110000110011010;
    rom[39408] = 25'b0000100100110000111010111;
    rom[39409] = 25'b0000100100110001000010010;
    rom[39410] = 25'b0000100100110001001001100;
    rom[39411] = 25'b0000100100110001010000100;
    rom[39412] = 25'b0000100100110001010111010;
    rom[39413] = 25'b0000100100110001011101111;
    rom[39414] = 25'b0000100100110001100100010;
    rom[39415] = 25'b0000100100110001101010011;
    rom[39416] = 25'b0000100100110001110000011;
    rom[39417] = 25'b0000100100110001110110001;
    rom[39418] = 25'b0000100100110001111011110;
    rom[39419] = 25'b0000100100110010000001000;
    rom[39420] = 25'b0000100100110010000110001;
    rom[39421] = 25'b0000100100110010001011001;
    rom[39422] = 25'b0000100100110010001111111;
    rom[39423] = 25'b0000100100110010010100011;
    rom[39424] = 25'b0000100100110010011000101;
    rom[39425] = 25'b0000100100110010011100110;
    rom[39426] = 25'b0000100100110010100000101;
    rom[39427] = 25'b0000100100110010100100011;
    rom[39428] = 25'b0000100100110010100111111;
    rom[39429] = 25'b0000100100110010101011001;
    rom[39430] = 25'b0000100100110010101110010;
    rom[39431] = 25'b0000100100110010110001000;
    rom[39432] = 25'b0000100100110010110011110;
    rom[39433] = 25'b0000100100110010110110001;
    rom[39434] = 25'b0000100100110010111000011;
    rom[39435] = 25'b0000100100110010111010100;
    rom[39436] = 25'b0000100100110010111100011;
    rom[39437] = 25'b0000100100110010111101111;
    rom[39438] = 25'b0000100100110010111111010;
    rom[39439] = 25'b0000100100110011000000100;
    rom[39440] = 25'b0000100100110011000001100;
    rom[39441] = 25'b0000100100110011000010011;
    rom[39442] = 25'b0000100100110011000011000;
    rom[39443] = 25'b0000100100110011000011011;
    rom[39444] = 25'b0000100100110011000011101;
    rom[39445] = 25'b0000100100110011000011101;
    rom[39446] = 25'b0000100100110011000011011;
    rom[39447] = 25'b0000100100110011000011000;
    rom[39448] = 25'b0000100100110011000010010;
    rom[39449] = 25'b0000100100110011000001100;
    rom[39450] = 25'b0000100100110011000000011;
    rom[39451] = 25'b0000100100110010111111010;
    rom[39452] = 25'b0000100100110010111101110;
    rom[39453] = 25'b0000100100110010111100001;
    rom[39454] = 25'b0000100100110010111010010;
    rom[39455] = 25'b0000100100110010111000010;
    rom[39456] = 25'b0000100100110010110101111;
    rom[39457] = 25'b0000100100110010110011100;
    rom[39458] = 25'b0000100100110010110000111;
    rom[39459] = 25'b0000100100110010101101111;
    rom[39460] = 25'b0000100100110010101010111;
    rom[39461] = 25'b0000100100110010100111101;
    rom[39462] = 25'b0000100100110010100100000;
    rom[39463] = 25'b0000100100110010100000011;
    rom[39464] = 25'b0000100100110010011100100;
    rom[39465] = 25'b0000100100110010011000100;
    rom[39466] = 25'b0000100100110010010100001;
    rom[39467] = 25'b0000100100110010001111101;
    rom[39468] = 25'b0000100100110010001010111;
    rom[39469] = 25'b0000100100110010000110000;
    rom[39470] = 25'b0000100100110010000000111;
    rom[39471] = 25'b0000100100110001111011101;
    rom[39472] = 25'b0000100100110001110110001;
    rom[39473] = 25'b0000100100110001110000011;
    rom[39474] = 25'b0000100100110001101010100;
    rom[39475] = 25'b0000100100110001100100011;
    rom[39476] = 25'b0000100100110001011110001;
    rom[39477] = 25'b0000100100110001010111100;
    rom[39478] = 25'b0000100100110001010000111;
    rom[39479] = 25'b0000100100110001001001111;
    rom[39480] = 25'b0000100100110001000010110;
    rom[39481] = 25'b0000100100110000111011100;
    rom[39482] = 25'b0000100100110000110011111;
    rom[39483] = 25'b0000100100110000101100010;
    rom[39484] = 25'b0000100100110000100100010;
    rom[39485] = 25'b0000100100110000011100001;
    rom[39486] = 25'b0000100100110000010011111;
    rom[39487] = 25'b0000100100110000001011010;
    rom[39488] = 25'b0000100100110000000010101;
    rom[39489] = 25'b0000100100101111111001101;
    rom[39490] = 25'b0000100100101111110000100;
    rom[39491] = 25'b0000100100101111100111001;
    rom[39492] = 25'b0000100100101111011101101;
    rom[39493] = 25'b0000100100101111010011111;
    rom[39494] = 25'b0000100100101111001010000;
    rom[39495] = 25'b0000100100101110111111110;
    rom[39496] = 25'b0000100100101110110101100;
    rom[39497] = 25'b0000100100101110101011000;
    rom[39498] = 25'b0000100100101110100000010;
    rom[39499] = 25'b0000100100101110010101010;
    rom[39500] = 25'b0000100100101110001010010;
    rom[39501] = 25'b0000100100101101111110111;
    rom[39502] = 25'b0000100100101101110011010;
    rom[39503] = 25'b0000100100101101100111101;
    rom[39504] = 25'b0000100100101101011011101;
    rom[39505] = 25'b0000100100101101001111100;
    rom[39506] = 25'b0000100100101101000011010;
    rom[39507] = 25'b0000100100101100110110110;
    rom[39508] = 25'b0000100100101100101010000;
    rom[39509] = 25'b0000100100101100011101001;
    rom[39510] = 25'b0000100100101100010000000;
    rom[39511] = 25'b0000100100101100000010101;
    rom[39512] = 25'b0000100100101011110101001;
    rom[39513] = 25'b0000100100101011100111011;
    rom[39514] = 25'b0000100100101011011001100;
    rom[39515] = 25'b0000100100101011001011011;
    rom[39516] = 25'b0000100100101010111101001;
    rom[39517] = 25'b0000100100101010101110101;
    rom[39518] = 25'b0000100100101010011111111;
    rom[39519] = 25'b0000100100101010010001000;
    rom[39520] = 25'b0000100100101010000001111;
    rom[39521] = 25'b0000100100101001110010101;
    rom[39522] = 25'b0000100100101001100011001;
    rom[39523] = 25'b0000100100101001010011100;
    rom[39524] = 25'b0000100100101001000011101;
    rom[39525] = 25'b0000100100101000110011100;
    rom[39526] = 25'b0000100100101000100011010;
    rom[39527] = 25'b0000100100101000010010110;
    rom[39528] = 25'b0000100100101000000010001;
    rom[39529] = 25'b0000100100100111110001010;
    rom[39530] = 25'b0000100100100111100000001;
    rom[39531] = 25'b0000100100100111001111000;
    rom[39532] = 25'b0000100100100110111101100;
    rom[39533] = 25'b0000100100100110101011111;
    rom[39534] = 25'b0000100100100110011010000;
    rom[39535] = 25'b0000100100100110001000000;
    rom[39536] = 25'b0000100100100101110101110;
    rom[39537] = 25'b0000100100100101100011010;
    rom[39538] = 25'b0000100100100101010000110;
    rom[39539] = 25'b0000100100100100111101111;
    rom[39540] = 25'b0000100100100100101010111;
    rom[39541] = 25'b0000100100100100010111101;
    rom[39542] = 25'b0000100100100100000100011;
    rom[39543] = 25'b0000100100100011110000110;
    rom[39544] = 25'b0000100100100011011100111;
    rom[39545] = 25'b0000100100100011001000111;
    rom[39546] = 25'b0000100100100010110100110;
    rom[39547] = 25'b0000100100100010100000011;
    rom[39548] = 25'b0000100100100010001011111;
    rom[39549] = 25'b0000100100100001110111000;
    rom[39550] = 25'b0000100100100001100010001;
    rom[39551] = 25'b0000100100100001001101000;
    rom[39552] = 25'b0000100100100000110111101;
    rom[39553] = 25'b0000100100100000100010001;
    rom[39554] = 25'b0000100100100000001100011;
    rom[39555] = 25'b0000100100011111110110011;
    rom[39556] = 25'b0000100100011111100000010;
    rom[39557] = 25'b0000100100011111001010001;
    rom[39558] = 25'b0000100100011110110011101;
    rom[39559] = 25'b0000100100011110011100111;
    rom[39560] = 25'b0000100100011110000110000;
    rom[39561] = 25'b0000100100011101101110111;
    rom[39562] = 25'b0000100100011101010111101;
    rom[39563] = 25'b0000100100011101000000001;
    rom[39564] = 25'b0000100100011100101000100;
    rom[39565] = 25'b0000100100011100010000110;
    rom[39566] = 25'b0000100100011011111000110;
    rom[39567] = 25'b0000100100011011100000011;
    rom[39568] = 25'b0000100100011011001000000;
    rom[39569] = 25'b0000100100011010101111011;
    rom[39570] = 25'b0000100100011010010110101;
    rom[39571] = 25'b0000100100011001111101101;
    rom[39572] = 25'b0000100100011001100100011;
    rom[39573] = 25'b0000100100011001001011001;
    rom[39574] = 25'b0000100100011000110001100;
    rom[39575] = 25'b0000100100011000010111110;
    rom[39576] = 25'b0000100100010111111101111;
    rom[39577] = 25'b0000100100010111100011110;
    rom[39578] = 25'b0000100100010111001001011;
    rom[39579] = 25'b0000100100010110101110111;
    rom[39580] = 25'b0000100100010110010100001;
    rom[39581] = 25'b0000100100010101111001010;
    rom[39582] = 25'b0000100100010101011110001;
    rom[39583] = 25'b0000100100010101000010111;
    rom[39584] = 25'b0000100100010100100111100;
    rom[39585] = 25'b0000100100010100001011110;
    rom[39586] = 25'b0000100100010011110000000;
    rom[39587] = 25'b0000100100010011010100000;
    rom[39588] = 25'b0000100100010010110111101;
    rom[39589] = 25'b0000100100010010011011010;
    rom[39590] = 25'b0000100100010001111110110;
    rom[39591] = 25'b0000100100010001100001111;
    rom[39592] = 25'b0000100100010001000100111;
    rom[39593] = 25'b0000100100010000100111110;
    rom[39594] = 25'b0000100100010000001010011;
    rom[39595] = 25'b0000100100001111101100111;
    rom[39596] = 25'b0000100100001111001111001;
    rom[39597] = 25'b0000100100001110110001010;
    rom[39598] = 25'b0000100100001110010011001;
    rom[39599] = 25'b0000100100001101110100111;
    rom[39600] = 25'b0000100100001101010110011;
    rom[39601] = 25'b0000100100001100110111110;
    rom[39602] = 25'b0000100100001100011000111;
    rom[39603] = 25'b0000100100001011111001111;
    rom[39604] = 25'b0000100100001011011010101;
    rom[39605] = 25'b0000100100001010111011001;
    rom[39606] = 25'b0000100100001010011011101;
    rom[39607] = 25'b0000100100001001111011110;
    rom[39608] = 25'b0000100100001001011011111;
    rom[39609] = 25'b0000100100001000111011110;
    rom[39610] = 25'b0000100100001000011011010;
    rom[39611] = 25'b0000100100000111111010110;
    rom[39612] = 25'b0000100100000111011010001;
    rom[39613] = 25'b0000100100000110111001001;
    rom[39614] = 25'b0000100100000110011000001;
    rom[39615] = 25'b0000100100000101110110111;
    rom[39616] = 25'b0000100100000101010101011;
    rom[39617] = 25'b0000100100000100110011110;
    rom[39618] = 25'b0000100100000100010001111;
    rom[39619] = 25'b0000100100000011101111111;
    rom[39620] = 25'b0000100100000011001101110;
    rom[39621] = 25'b0000100100000010101011010;
    rom[39622] = 25'b0000100100000010001000110;
    rom[39623] = 25'b0000100100000001100110000;
    rom[39624] = 25'b0000100100000001000011000;
    rom[39625] = 25'b0000100100000000011111111;
    rom[39626] = 25'b0000100011111111111100101;
    rom[39627] = 25'b0000100011111111011001001;
    rom[39628] = 25'b0000100011111110110101100;
    rom[39629] = 25'b0000100011111110010001101;
    rom[39630] = 25'b0000100011111101101101100;
    rom[39631] = 25'b0000100011111101001001011;
    rom[39632] = 25'b0000100011111100100100111;
    rom[39633] = 25'b0000100011111100000000011;
    rom[39634] = 25'b0000100011111011011011101;
    rom[39635] = 25'b0000100011111010110110101;
    rom[39636] = 25'b0000100011111010010001100;
    rom[39637] = 25'b0000100011111001101100001;
    rom[39638] = 25'b0000100011111001000110101;
    rom[39639] = 25'b0000100011111000100001000;
    rom[39640] = 25'b0000100011110111111011001;
    rom[39641] = 25'b0000100011110111010101001;
    rom[39642] = 25'b0000100011110110101110110;
    rom[39643] = 25'b0000100011110110001000011;
    rom[39644] = 25'b0000100011110101100001111;
    rom[39645] = 25'b0000100011110100111011000;
    rom[39646] = 25'b0000100011110100010100000;
    rom[39647] = 25'b0000100011110011101100111;
    rom[39648] = 25'b0000100011110011000101101;
    rom[39649] = 25'b0000100011110010011110001;
    rom[39650] = 25'b0000100011110001110110011;
    rom[39651] = 25'b0000100011110001001110100;
    rom[39652] = 25'b0000100011110000100110101;
    rom[39653] = 25'b0000100011101111111110011;
    rom[39654] = 25'b0000100011101111010101111;
    rom[39655] = 25'b0000100011101110101101011;
    rom[39656] = 25'b0000100011101110000100100;
    rom[39657] = 25'b0000100011101101011011101;
    rom[39658] = 25'b0000100011101100110010100;
    rom[39659] = 25'b0000100011101100001001001;
    rom[39660] = 25'b0000100011101011011111110;
    rom[39661] = 25'b0000100011101010110110000;
    rom[39662] = 25'b0000100011101010001100010;
    rom[39663] = 25'b0000100011101001100010010;
    rom[39664] = 25'b0000100011101000111000000;
    rom[39665] = 25'b0000100011101000001101101;
    rom[39666] = 25'b0000100011100111100011000;
    rom[39667] = 25'b0000100011100110111000011;
    rom[39668] = 25'b0000100011100110001101011;
    rom[39669] = 25'b0000100011100101100010011;
    rom[39670] = 25'b0000100011100100110111001;
    rom[39671] = 25'b0000100011100100001011100;
    rom[39672] = 25'b0000100011100011100000000;
    rom[39673] = 25'b0000100011100010110100001;
    rom[39674] = 25'b0000100011100010001000001;
    rom[39675] = 25'b0000100011100001011100000;
    rom[39676] = 25'b0000100011100000101111110;
    rom[39677] = 25'b0000100011100000000011001;
    rom[39678] = 25'b0000100011011111010110100;
    rom[39679] = 25'b0000100011011110101001101;
    rom[39680] = 25'b0000100011011101111100101;
    rom[39681] = 25'b0000100011011101001111011;
    rom[39682] = 25'b0000100011011100100001111;
    rom[39683] = 25'b0000100011011011110100011;
    rom[39684] = 25'b0000100011011011000110110;
    rom[39685] = 25'b0000100011011010011000110;
    rom[39686] = 25'b0000100011011001101010101;
    rom[39687] = 25'b0000100011011000111100011;
    rom[39688] = 25'b0000100011011000001101111;
    rom[39689] = 25'b0000100011010111011111010;
    rom[39690] = 25'b0000100011010110110000100;
    rom[39691] = 25'b0000100011010110000001100;
    rom[39692] = 25'b0000100011010101010010011;
    rom[39693] = 25'b0000100011010100100011000;
    rom[39694] = 25'b0000100011010011110011101;
    rom[39695] = 25'b0000100011010011000011111;
    rom[39696] = 25'b0000100011010010010100000;
    rom[39697] = 25'b0000100011010001100100000;
    rom[39698] = 25'b0000100011010000110011110;
    rom[39699] = 25'b0000100011010000000011011;
    rom[39700] = 25'b0000100011001111010010111;
    rom[39701] = 25'b0000100011001110100010001;
    rom[39702] = 25'b0000100011001101110001010;
    rom[39703] = 25'b0000100011001101000000010;
    rom[39704] = 25'b0000100011001100001111000;
    rom[39705] = 25'b0000100011001011011101101;
    rom[39706] = 25'b0000100011001010101100000;
    rom[39707] = 25'b0000100011001001111010010;
    rom[39708] = 25'b0000100011001001001000010;
    rom[39709] = 25'b0000100011001000010110010;
    rom[39710] = 25'b0000100011000111100100000;
    rom[39711] = 25'b0000100011000110110001100;
    rom[39712] = 25'b0000100011000101111110111;
    rom[39713] = 25'b0000100011000101001100000;
    rom[39714] = 25'b0000100011000100011001001;
    rom[39715] = 25'b0000100011000011100110000;
    rom[39716] = 25'b0000100011000010110010101;
    rom[39717] = 25'b0000100011000001111111010;
    rom[39718] = 25'b0000100011000001001011101;
    rom[39719] = 25'b0000100011000000010111110;
    rom[39720] = 25'b0000100010111111100011110;
    rom[39721] = 25'b0000100010111110101111101;
    rom[39722] = 25'b0000100010111101111011010;
    rom[39723] = 25'b0000100010111101000110110;
    rom[39724] = 25'b0000100010111100010010001;
    rom[39725] = 25'b0000100010111011011101010;
    rom[39726] = 25'b0000100010111010101000010;
    rom[39727] = 25'b0000100010111001110011000;
    rom[39728] = 25'b0000100010111000111101110;
    rom[39729] = 25'b0000100010111000001000010;
    rom[39730] = 25'b0000100010110111010010100;
    rom[39731] = 25'b0000100010110110011100101;
    rom[39732] = 25'b0000100010110101100110101;
    rom[39733] = 25'b0000100010110100110000011;
    rom[39734] = 25'b0000100010110011111010000;
    rom[39735] = 25'b0000100010110011000011100;
    rom[39736] = 25'b0000100010110010001100111;
    rom[39737] = 25'b0000100010110001010110000;
    rom[39738] = 25'b0000100010110000011111000;
    rom[39739] = 25'b0000100010101111100111110;
    rom[39740] = 25'b0000100010101110110000011;
    rom[39741] = 25'b0000100010101101111000111;
    rom[39742] = 25'b0000100010101101000001001;
    rom[39743] = 25'b0000100010101100001001010;
    rom[39744] = 25'b0000100010101011010001010;
    rom[39745] = 25'b0000100010101010011001000;
    rom[39746] = 25'b0000100010101001100000101;
    rom[39747] = 25'b0000100010101000101000001;
    rom[39748] = 25'b0000100010100111101111011;
    rom[39749] = 25'b0000100010100110110110100;
    rom[39750] = 25'b0000100010100101111101100;
    rom[39751] = 25'b0000100010100101000100010;
    rom[39752] = 25'b0000100010100100001010111;
    rom[39753] = 25'b0000100010100011010001011;
    rom[39754] = 25'b0000100010100010010111101;
    rom[39755] = 25'b0000100010100001011101110;
    rom[39756] = 25'b0000100010100000100011110;
    rom[39757] = 25'b0000100010011111101001100;
    rom[39758] = 25'b0000100010011110101111001;
    rom[39759] = 25'b0000100010011101110100101;
    rom[39760] = 25'b0000100010011100111001111;
    rom[39761] = 25'b0000100010011011111111000;
    rom[39762] = 25'b0000100010011011000100000;
    rom[39763] = 25'b0000100010011010001000111;
    rom[39764] = 25'b0000100010011001001101100;
    rom[39765] = 25'b0000100010011000010010000;
    rom[39766] = 25'b0000100010010111010110010;
    rom[39767] = 25'b0000100010010110011010011;
    rom[39768] = 25'b0000100010010101011110100;
    rom[39769] = 25'b0000100010010100100010010;
    rom[39770] = 25'b0000100010010011100101111;
    rom[39771] = 25'b0000100010010010101001100;
    rom[39772] = 25'b0000100010010001101100110;
    rom[39773] = 25'b0000100010010000110000000;
    rom[39774] = 25'b0000100010001111110011000;
    rom[39775] = 25'b0000100010001110110101111;
    rom[39776] = 25'b0000100010001101111000100;
    rom[39777] = 25'b0000100010001100111011000;
    rom[39778] = 25'b0000100010001011111101011;
    rom[39779] = 25'b0000100010001010111111101;
    rom[39780] = 25'b0000100010001010000001101;
    rom[39781] = 25'b0000100010001001000011100;
    rom[39782] = 25'b0000100010001000000101010;
    rom[39783] = 25'b0000100010000111000110110;
    rom[39784] = 25'b0000100010000110001000010;
    rom[39785] = 25'b0000100010000101001001100;
    rom[39786] = 25'b0000100010000100001010100;
    rom[39787] = 25'b0000100010000011001011100;
    rom[39788] = 25'b0000100010000010001100010;
    rom[39789] = 25'b0000100010000001001100111;
    rom[39790] = 25'b0000100010000000001101010;
    rom[39791] = 25'b0000100001111111001101100;
    rom[39792] = 25'b0000100001111110001101101;
    rom[39793] = 25'b0000100001111101001101101;
    rom[39794] = 25'b0000100001111100001101011;
    rom[39795] = 25'b0000100001111011001101000;
    rom[39796] = 25'b0000100001111010001100100;
    rom[39797] = 25'b0000100001111001001011111;
    rom[39798] = 25'b0000100001111000001011000;
    rom[39799] = 25'b0000100001110111001010000;
    rom[39800] = 25'b0000100001110110001000111;
    rom[39801] = 25'b0000100001110101000111100;
    rom[39802] = 25'b0000100001110100000110000;
    rom[39803] = 25'b0000100001110011000100011;
    rom[39804] = 25'b0000100001110010000010101;
    rom[39805] = 25'b0000100001110001000000110;
    rom[39806] = 25'b0000100001101111111110101;
    rom[39807] = 25'b0000100001101110111100010;
    rom[39808] = 25'b0000100001101101111001111;
    rom[39809] = 25'b0000100001101100110111010;
    rom[39810] = 25'b0000100001101011110100101;
    rom[39811] = 25'b0000100001101010110001110;
    rom[39812] = 25'b0000100001101001101110110;
    rom[39813] = 25'b0000100001101000101011100;
    rom[39814] = 25'b0000100001100111101000001;
    rom[39815] = 25'b0000100001100110100100101;
    rom[39816] = 25'b0000100001100101100000111;
    rom[39817] = 25'b0000100001100100011101001;
    rom[39818] = 25'b0000100001100011011001001;
    rom[39819] = 25'b0000100001100010010101000;
    rom[39820] = 25'b0000100001100001010000110;
    rom[39821] = 25'b0000100001100000001100011;
    rom[39822] = 25'b0000100001011111000111110;
    rom[39823] = 25'b0000100001011110000011000;
    rom[39824] = 25'b0000100001011100111110000;
    rom[39825] = 25'b0000100001011011111000111;
    rom[39826] = 25'b0000100001011010110011110;
    rom[39827] = 25'b0000100001011001101110011;
    rom[39828] = 25'b0000100001011000101000111;
    rom[39829] = 25'b0000100001010111100011010;
    rom[39830] = 25'b0000100001010110011101011;
    rom[39831] = 25'b0000100001010101010111011;
    rom[39832] = 25'b0000100001010100010001010;
    rom[39833] = 25'b0000100001010011001011000;
    rom[39834] = 25'b0000100001010010000100100;
    rom[39835] = 25'b0000100001010000111101111;
    rom[39836] = 25'b0000100001001111110111001;
    rom[39837] = 25'b0000100001001110110000010;
    rom[39838] = 25'b0000100001001101101001010;
    rom[39839] = 25'b0000100001001100100010000;
    rom[39840] = 25'b0000100001001011011010101;
    rom[39841] = 25'b0000100001001010010011001;
    rom[39842] = 25'b0000100001001001001011011;
    rom[39843] = 25'b0000100001001000000011101;
    rom[39844] = 25'b0000100001000110111011110;
    rom[39845] = 25'b0000100001000101110011101;
    rom[39846] = 25'b0000100001000100101011011;
    rom[39847] = 25'b0000100001000011100010111;
    rom[39848] = 25'b0000100001000010011010010;
    rom[39849] = 25'b0000100001000001010001101;
    rom[39850] = 25'b0000100001000000001000110;
    rom[39851] = 25'b0000100000111110111111110;
    rom[39852] = 25'b0000100000111101110110101;
    rom[39853] = 25'b0000100000111100101101010;
    rom[39854] = 25'b0000100000111011100011110;
    rom[39855] = 25'b0000100000111010011010001;
    rom[39856] = 25'b0000100000111001010000011;
    rom[39857] = 25'b0000100000111000000110100;
    rom[39858] = 25'b0000100000110110111100100;
    rom[39859] = 25'b0000100000110101110010010;
    rom[39860] = 25'b0000100000110100100111111;
    rom[39861] = 25'b0000100000110011011101011;
    rom[39862] = 25'b0000100000110010010010110;
    rom[39863] = 25'b0000100000110001001000000;
    rom[39864] = 25'b0000100000101111111101000;
    rom[39865] = 25'b0000100000101110110001111;
    rom[39866] = 25'b0000100000101101100110101;
    rom[39867] = 25'b0000100000101100011011010;
    rom[39868] = 25'b0000100000101011001111110;
    rom[39869] = 25'b0000100000101010000100000;
    rom[39870] = 25'b0000100000101000111000001;
    rom[39871] = 25'b0000100000100111101100010;
    rom[39872] = 25'b0000100000100110100000001;
    rom[39873] = 25'b0000100000100101010011110;
    rom[39874] = 25'b0000100000100100000111011;
    rom[39875] = 25'b0000100000100010111010111;
    rom[39876] = 25'b0000100000100001101110000;
    rom[39877] = 25'b0000100000100000100001010;
    rom[39878] = 25'b0000100000011111010100010;
    rom[39879] = 25'b0000100000011110000111001;
    rom[39880] = 25'b0000100000011100111001110;
    rom[39881] = 25'b0000100000011011101100011;
    rom[39882] = 25'b0000100000011010011110110;
    rom[39883] = 25'b0000100000011001010001001;
    rom[39884] = 25'b0000100000011000000011001;
    rom[39885] = 25'b0000100000010110110101001;
    rom[39886] = 25'b0000100000010101100111000;
    rom[39887] = 25'b0000100000010100011000110;
    rom[39888] = 25'b0000100000010011001010010;
    rom[39889] = 25'b0000100000010001111011101;
    rom[39890] = 25'b0000100000010000101100111;
    rom[39891] = 25'b0000100000001111011110001;
    rom[39892] = 25'b0000100000001110001111000;
    rom[39893] = 25'b0000100000001100111111111;
    rom[39894] = 25'b0000100000001011110000101;
    rom[39895] = 25'b0000100000001010100001001;
    rom[39896] = 25'b0000100000001001010001100;
    rom[39897] = 25'b0000100000001000000001110;
    rom[39898] = 25'b0000100000000110110001111;
    rom[39899] = 25'b0000100000000101100001111;
    rom[39900] = 25'b0000100000000100010001110;
    rom[39901] = 25'b0000100000000011000001011;
    rom[39902] = 25'b0000100000000001110001000;
    rom[39903] = 25'b0000100000000000100000011;
    rom[39904] = 25'b0000011111111111001111110;
    rom[39905] = 25'b0000011111111101111110111;
    rom[39906] = 25'b0000011111111100101101110;
    rom[39907] = 25'b0000011111111011011100101;
    rom[39908] = 25'b0000011111111010001011011;
    rom[39909] = 25'b0000011111111000111001111;
    rom[39910] = 25'b0000011111110111101000011;
    rom[39911] = 25'b0000011111110110010110110;
    rom[39912] = 25'b0000011111110101000100110;
    rom[39913] = 25'b0000011111110011110010111;
    rom[39914] = 25'b0000011111110010100000110;
    rom[39915] = 25'b0000011111110001001110011;
    rom[39916] = 25'b0000011111101111111100001;
    rom[39917] = 25'b0000011111101110101001100;
    rom[39918] = 25'b0000011111101101010110111;
    rom[39919] = 25'b0000011111101100000100000;
    rom[39920] = 25'b0000011111101010110001001;
    rom[39921] = 25'b0000011111101001011110000;
    rom[39922] = 25'b0000011111101000001010110;
    rom[39923] = 25'b0000011111100110110111011;
    rom[39924] = 25'b0000011111100101100011111;
    rom[39925] = 25'b0000011111100100010000010;
    rom[39926] = 25'b0000011111100010111100100;
    rom[39927] = 25'b0000011111100001101000100;
    rom[39928] = 25'b0000011111100000010100100;
    rom[39929] = 25'b0000011111011111000000011;
    rom[39930] = 25'b0000011111011101101100000;
    rom[39931] = 25'b0000011111011100010111100;
    rom[39932] = 25'b0000011111011011000010111;
    rom[39933] = 25'b0000011111011001101110001;
    rom[39934] = 25'b0000011111011000011001010;
    rom[39935] = 25'b0000011111010111000100010;
    rom[39936] = 25'b0000011111010101101111001;
    rom[39937] = 25'b0000011111010100011001111;
    rom[39938] = 25'b0000011111010011000100011;
    rom[39939] = 25'b0000011111010001101110111;
    rom[39940] = 25'b0000011111010000011001010;
    rom[39941] = 25'b0000011111001111000011011;
    rom[39942] = 25'b0000011111001101101101100;
    rom[39943] = 25'b0000011111001100010111011;
    rom[39944] = 25'b0000011111001011000001001;
    rom[39945] = 25'b0000011111001001101010110;
    rom[39946] = 25'b0000011111001000010100011;
    rom[39947] = 25'b0000011111000110111101101;
    rom[39948] = 25'b0000011111000101100110111;
    rom[39949] = 25'b0000011111000100010000000;
    rom[39950] = 25'b0000011111000010111001000;
    rom[39951] = 25'b0000011111000001100001111;
    rom[39952] = 25'b0000011111000000001010101;
    rom[39953] = 25'b0000011110111110110011001;
    rom[39954] = 25'b0000011110111101011011101;
    rom[39955] = 25'b0000011110111100000100000;
    rom[39956] = 25'b0000011110111010101100001;
    rom[39957] = 25'b0000011110111001010100010;
    rom[39958] = 25'b0000011110110111111100001;
    rom[39959] = 25'b0000011110110110100011111;
    rom[39960] = 25'b0000011110110101001011100;
    rom[39961] = 25'b0000011110110011110011001;
    rom[39962] = 25'b0000011110110010011010100;
    rom[39963] = 25'b0000011110110001000001110;
    rom[39964] = 25'b0000011110101111101000111;
    rom[39965] = 25'b0000011110101110001111111;
    rom[39966] = 25'b0000011110101100110110110;
    rom[39967] = 25'b0000011110101011011101100;
    rom[39968] = 25'b0000011110101010000100001;
    rom[39969] = 25'b0000011110101000101010101;
    rom[39970] = 25'b0000011110100111010001000;
    rom[39971] = 25'b0000011110100101110111010;
    rom[39972] = 25'b0000011110100100011101011;
    rom[39973] = 25'b0000011110100011000011011;
    rom[39974] = 25'b0000011110100001101001010;
    rom[39975] = 25'b0000011110100000001110111;
    rom[39976] = 25'b0000011110011110110100100;
    rom[39977] = 25'b0000011110011101011001111;
    rom[39978] = 25'b0000011110011011111111011;
    rom[39979] = 25'b0000011110011010100100100;
    rom[39980] = 25'b0000011110011001001001101;
    rom[39981] = 25'b0000011110010111101110100;
    rom[39982] = 25'b0000011110010110010011010;
    rom[39983] = 25'b0000011110010100111000001;
    rom[39984] = 25'b0000011110010011011100101;
    rom[39985] = 25'b0000011110010010000001000;
    rom[39986] = 25'b0000011110010000100101011;
    rom[39987] = 25'b0000011110001111001001100;
    rom[39988] = 25'b0000011110001101101101101;
    rom[39989] = 25'b0000011110001100010001100;
    rom[39990] = 25'b0000011110001010110101011;
    rom[39991] = 25'b0000011110001001011001001;
    rom[39992] = 25'b0000011110000111111100101;
    rom[39993] = 25'b0000011110000110100000001;
    rom[39994] = 25'b0000011110000101000011011;
    rom[39995] = 25'b0000011110000011100110100;
    rom[39996] = 25'b0000011110000010001001101;
    rom[39997] = 25'b0000011110000000101100101;
    rom[39998] = 25'b0000011101111111001111011;
    rom[39999] = 25'b0000011101111101110010001;
    rom[40000] = 25'b0000011101111100010100101;
    rom[40001] = 25'b0000011101111010110111001;
    rom[40002] = 25'b0000011101111001011001011;
    rom[40003] = 25'b0000011101110111111011101;
    rom[40004] = 25'b0000011101110110011101110;
    rom[40005] = 25'b0000011101110100111111101;
    rom[40006] = 25'b0000011101110011100001011;
    rom[40007] = 25'b0000011101110010000011010;
    rom[40008] = 25'b0000011101110000100100110;
    rom[40009] = 25'b0000011101101111000110001;
    rom[40010] = 25'b0000011101101101100111101;
    rom[40011] = 25'b0000011101101100001000110;
    rom[40012] = 25'b0000011101101010101001111;
    rom[40013] = 25'b0000011101101001001010111;
    rom[40014] = 25'b0000011101100111101011101;
    rom[40015] = 25'b0000011101100110001100011;
    rom[40016] = 25'b0000011101100100101101000;
    rom[40017] = 25'b0000011101100011001101100;
    rom[40018] = 25'b0000011101100001101101111;
    rom[40019] = 25'b0000011101100000001110001;
    rom[40020] = 25'b0000011101011110101110010;
    rom[40021] = 25'b0000011101011101001110010;
    rom[40022] = 25'b0000011101011011101110010;
    rom[40023] = 25'b0000011101011010001101111;
    rom[40024] = 25'b0000011101011000101101101;
    rom[40025] = 25'b0000011101010111001101001;
    rom[40026] = 25'b0000011101010101101100100;
    rom[40027] = 25'b0000011101010100001011111;
    rom[40028] = 25'b0000011101010010101011000;
    rom[40029] = 25'b0000011101010001001010001;
    rom[40030] = 25'b0000011101001111101001000;
    rom[40031] = 25'b0000011101001110000111111;
    rom[40032] = 25'b0000011101001100100110100;
    rom[40033] = 25'b0000011101001011000101001;
    rom[40034] = 25'b0000011101001001100011100;
    rom[40035] = 25'b0000011101001000000001111;
    rom[40036] = 25'b0000011101000110100000001;
    rom[40037] = 25'b0000011101000100111110010;
    rom[40038] = 25'b0000011101000011011100010;
    rom[40039] = 25'b0000011101000001111010001;
    rom[40040] = 25'b0000011101000000010111111;
    rom[40041] = 25'b0000011100111110110101100;
    rom[40042] = 25'b0000011100111101010011001;
    rom[40043] = 25'b0000011100111011110000100;
    rom[40044] = 25'b0000011100111010001101111;
    rom[40045] = 25'b0000011100111000101011000;
    rom[40046] = 25'b0000011100110111001000000;
    rom[40047] = 25'b0000011100110101100101000;
    rom[40048] = 25'b0000011100110100000001111;
    rom[40049] = 25'b0000011100110010011110101;
    rom[40050] = 25'b0000011100110000111011001;
    rom[40051] = 25'b0000011100101111010111110;
    rom[40052] = 25'b0000011100101101110100000;
    rom[40053] = 25'b0000011100101100010000010;
    rom[40054] = 25'b0000011100101010101100100;
    rom[40055] = 25'b0000011100101001001000100;
    rom[40056] = 25'b0000011100100111100100100;
    rom[40057] = 25'b0000011100100110000000010;
    rom[40058] = 25'b0000011100100100011100000;
    rom[40059] = 25'b0000011100100010110111100;
    rom[40060] = 25'b0000011100100001010011000;
    rom[40061] = 25'b0000011100011111101110011;
    rom[40062] = 25'b0000011100011110001001101;
    rom[40063] = 25'b0000011100011100100100110;
    rom[40064] = 25'b0000011100011010111111111;
    rom[40065] = 25'b0000011100011001011010101;
    rom[40066] = 25'b0000011100010111110101100;
    rom[40067] = 25'b0000011100010110010000010;
    rom[40068] = 25'b0000011100010100101010110;
    rom[40069] = 25'b0000011100010011000101010;
    rom[40070] = 25'b0000011100010001011111101;
    rom[40071] = 25'b0000011100001111111001110;
    rom[40072] = 25'b0000011100001110010100000;
    rom[40073] = 25'b0000011100001100101110000;
    rom[40074] = 25'b0000011100001011001000000;
    rom[40075] = 25'b0000011100001001100001110;
    rom[40076] = 25'b0000011100000111111011100;
    rom[40077] = 25'b0000011100000110010101000;
    rom[40078] = 25'b0000011100000100101110100;
    rom[40079] = 25'b0000011100000011000111111;
    rom[40080] = 25'b0000011100000001100001001;
    rom[40081] = 25'b0000011011111111111010010;
    rom[40082] = 25'b0000011011111110010011010;
    rom[40083] = 25'b0000011011111100101100010;
    rom[40084] = 25'b0000011011111011000101001;
    rom[40085] = 25'b0000011011111001011101110;
    rom[40086] = 25'b0000011011110111110110011;
    rom[40087] = 25'b0000011011110110001110111;
    rom[40088] = 25'b0000011011110100100111010;
    rom[40089] = 25'b0000011011110010111111100;
    rom[40090] = 25'b0000011011110001010111110;
    rom[40091] = 25'b0000011011101111101111111;
    rom[40092] = 25'b0000011011101110000111110;
    rom[40093] = 25'b0000011011101100011111101;
    rom[40094] = 25'b0000011011101010110111011;
    rom[40095] = 25'b0000011011101001001111000;
    rom[40096] = 25'b0000011011100111100110100;
    rom[40097] = 25'b0000011011100101111110000;
    rom[40098] = 25'b0000011011100100010101011;
    rom[40099] = 25'b0000011011100010101100101;
    rom[40100] = 25'b0000011011100001000011110;
    rom[40101] = 25'b0000011011011111011010110;
    rom[40102] = 25'b0000011011011101110001101;
    rom[40103] = 25'b0000011011011100001000011;
    rom[40104] = 25'b0000011011011010011111001;
    rom[40105] = 25'b0000011011011000110101110;
    rom[40106] = 25'b0000011011010111001100010;
    rom[40107] = 25'b0000011011010101100010101;
    rom[40108] = 25'b0000011011010011111000111;
    rom[40109] = 25'b0000011011010010001111001;
    rom[40110] = 25'b0000011011010000100101001;
    rom[40111] = 25'b0000011011001110111011001;
    rom[40112] = 25'b0000011011001101010001000;
    rom[40113] = 25'b0000011011001011100110110;
    rom[40114] = 25'b0000011011001001111100100;
    rom[40115] = 25'b0000011011001000010010000;
    rom[40116] = 25'b0000011011000110100111011;
    rom[40117] = 25'b0000011011000100111100110;
    rom[40118] = 25'b0000011011000011010010000;
    rom[40119] = 25'b0000011011000001100111010;
    rom[40120] = 25'b0000011010111111111100010;
    rom[40121] = 25'b0000011010111110010001010;
    rom[40122] = 25'b0000011010111100100110000;
    rom[40123] = 25'b0000011010111010111010111;
    rom[40124] = 25'b0000011010111001001111100;
    rom[40125] = 25'b0000011010110111100100000;
    rom[40126] = 25'b0000011010110101111000100;
    rom[40127] = 25'b0000011010110100001100110;
    rom[40128] = 25'b0000011010110010100001001;
    rom[40129] = 25'b0000011010110000110101010;
    rom[40130] = 25'b0000011010101111001001010;
    rom[40131] = 25'b0000011010101101011101010;
    rom[40132] = 25'b0000011010101011110001001;
    rom[40133] = 25'b0000011010101010000100111;
    rom[40134] = 25'b0000011010101000011000100;
    rom[40135] = 25'b0000011010100110101100000;
    rom[40136] = 25'b0000011010100100111111100;
    rom[40137] = 25'b0000011010100011010010111;
    rom[40138] = 25'b0000011010100001100110001;
    rom[40139] = 25'b0000011010011111111001011;
    rom[40140] = 25'b0000011010011110001100011;
    rom[40141] = 25'b0000011010011100011111011;
    rom[40142] = 25'b0000011010011010110010001;
    rom[40143] = 25'b0000011010011001000101000;
    rom[40144] = 25'b0000011010010111010111101;
    rom[40145] = 25'b0000011010010101101010010;
    rom[40146] = 25'b0000011010010011111100110;
    rom[40147] = 25'b0000011010010010001111001;
    rom[40148] = 25'b0000011010010000100001011;
    rom[40149] = 25'b0000011010001110110011101;
    rom[40150] = 25'b0000011010001101000101110;
    rom[40151] = 25'b0000011010001011010111110;
    rom[40152] = 25'b0000011010001001101001101;
    rom[40153] = 25'b0000011010000111111011011;
    rom[40154] = 25'b0000011010000110001101001;
    rom[40155] = 25'b0000011010000100011110110;
    rom[40156] = 25'b0000011010000010110000010;
    rom[40157] = 25'b0000011010000001000001110;
    rom[40158] = 25'b0000011001111111010011001;
    rom[40159] = 25'b0000011001111101100100011;
    rom[40160] = 25'b0000011001111011110101100;
    rom[40161] = 25'b0000011001111010000110101;
    rom[40162] = 25'b0000011001111000010111100;
    rom[40163] = 25'b0000011001110110101000011;
    rom[40164] = 25'b0000011001110100111001010;
    rom[40165] = 25'b0000011001110011001001111;
    rom[40166] = 25'b0000011001110001011010100;
    rom[40167] = 25'b0000011001101111101011000;
    rom[40168] = 25'b0000011001101101111011011;
    rom[40169] = 25'b0000011001101100001011110;
    rom[40170] = 25'b0000011001101010011100000;
    rom[40171] = 25'b0000011001101000101100001;
    rom[40172] = 25'b0000011001100110111100001;
    rom[40173] = 25'b0000011001100101001100001;
    rom[40174] = 25'b0000011001100011011100000;
    rom[40175] = 25'b0000011001100001101011110;
    rom[40176] = 25'b0000011001011111111011011;
    rom[40177] = 25'b0000011001011110001011000;
    rom[40178] = 25'b0000011001011100011010100;
    rom[40179] = 25'b0000011001011010101001111;
    rom[40180] = 25'b0000011001011000111001010;
    rom[40181] = 25'b0000011001010111001000100;
    rom[40182] = 25'b0000011001010101010111101;
    rom[40183] = 25'b0000011001010011100110101;
    rom[40184] = 25'b0000011001010001110101101;
    rom[40185] = 25'b0000011001010000000100100;
    rom[40186] = 25'b0000011001001110010011010;
    rom[40187] = 25'b0000011001001100100010000;
    rom[40188] = 25'b0000011001001010110000101;
    rom[40189] = 25'b0000011001001000111111001;
    rom[40190] = 25'b0000011001000111001101100;
    rom[40191] = 25'b0000011001000101011011111;
    rom[40192] = 25'b0000011001000011101010001;
    rom[40193] = 25'b0000011001000001111000011;
    rom[40194] = 25'b0000011001000000000110100;
    rom[40195] = 25'b0000011000111110010100011;
    rom[40196] = 25'b0000011000111100100010011;
    rom[40197] = 25'b0000011000111010110000010;
    rom[40198] = 25'b0000011000111000111101111;
    rom[40199] = 25'b0000011000110111001011101;
    rom[40200] = 25'b0000011000110101011001001;
    rom[40201] = 25'b0000011000110011100110101;
    rom[40202] = 25'b0000011000110001110100000;
    rom[40203] = 25'b0000011000110000000001011;
    rom[40204] = 25'b0000011000101110001110101;
    rom[40205] = 25'b0000011000101100011011110;
    rom[40206] = 25'b0000011000101010101000110;
    rom[40207] = 25'b0000011000101000110101101;
    rom[40208] = 25'b0000011000100111000010100;
    rom[40209] = 25'b0000011000100101001111011;
    rom[40210] = 25'b0000011000100011011100000;
    rom[40211] = 25'b0000011000100001101000110;
    rom[40212] = 25'b0000011000011111110101010;
    rom[40213] = 25'b0000011000011110000001110;
    rom[40214] = 25'b0000011000011100001110001;
    rom[40215] = 25'b0000011000011010011010011;
    rom[40216] = 25'b0000011000011000100110101;
    rom[40217] = 25'b0000011000010110110010110;
    rom[40218] = 25'b0000011000010100111110110;
    rom[40219] = 25'b0000011000010011001010110;
    rom[40220] = 25'b0000011000010001010110101;
    rom[40221] = 25'b0000011000001111100010100;
    rom[40222] = 25'b0000011000001101101110001;
    rom[40223] = 25'b0000011000001011111001111;
    rom[40224] = 25'b0000011000001010000101011;
    rom[40225] = 25'b0000011000001000010000111;
    rom[40226] = 25'b0000011000000110011100010;
    rom[40227] = 25'b0000011000000100100111100;
    rom[40228] = 25'b0000011000000010110010110;
    rom[40229] = 25'b0000011000000000111110000;
    rom[40230] = 25'b0000010111111111001001000;
    rom[40231] = 25'b0000010111111101010100000;
    rom[40232] = 25'b0000010111111011011110111;
    rom[40233] = 25'b0000010111111001101001111;
    rom[40234] = 25'b0000010111110111110100100;
    rom[40235] = 25'b0000010111110101111111010;
    rom[40236] = 25'b0000010111110100001001111;
    rom[40237] = 25'b0000010111110010010100011;
    rom[40238] = 25'b0000010111110000011110110;
    rom[40239] = 25'b0000010111101110101001001;
    rom[40240] = 25'b0000010111101100110011100;
    rom[40241] = 25'b0000010111101010111101101;
    rom[40242] = 25'b0000010111101001000111110;
    rom[40243] = 25'b0000010111100111010001110;
    rom[40244] = 25'b0000010111100101011011110;
    rom[40245] = 25'b0000010111100011100101101;
    rom[40246] = 25'b0000010111100001101111100;
    rom[40247] = 25'b0000010111011111111001010;
    rom[40248] = 25'b0000010111011110000011000;
    rom[40249] = 25'b0000010111011100001100100;
    rom[40250] = 25'b0000010111011010010110000;
    rom[40251] = 25'b0000010111011000011111011;
    rom[40252] = 25'b0000010111010110101000111;
    rom[40253] = 25'b0000010111010100110010001;
    rom[40254] = 25'b0000010111010010111011011;
    rom[40255] = 25'b0000010111010001000100100;
    rom[40256] = 25'b0000010111001111001101100;
    rom[40257] = 25'b0000010111001101010110100;
    rom[40258] = 25'b0000010111001011011111011;
    rom[40259] = 25'b0000010111001001101000001;
    rom[40260] = 25'b0000010111000111110001000;
    rom[40261] = 25'b0000010111000101111001101;
    rom[40262] = 25'b0000010111000100000010010;
    rom[40263] = 25'b0000010111000010001010110;
    rom[40264] = 25'b0000010111000000010011010;
    rom[40265] = 25'b0000010110111110011011101;
    rom[40266] = 25'b0000010110111100100100000;
    rom[40267] = 25'b0000010110111010101100010;
    rom[40268] = 25'b0000010110111000110100011;
    rom[40269] = 25'b0000010110110110111100100;
    rom[40270] = 25'b0000010110110101000100100;
    rom[40271] = 25'b0000010110110011001100100;
    rom[40272] = 25'b0000010110110001010100011;
    rom[40273] = 25'b0000010110101111011100001;
    rom[40274] = 25'b0000010110101101100011111;
    rom[40275] = 25'b0000010110101011101011101;
    rom[40276] = 25'b0000010110101001110011010;
    rom[40277] = 25'b0000010110100111111010110;
    rom[40278] = 25'b0000010110100110000010010;
    rom[40279] = 25'b0000010110100100001001100;
    rom[40280] = 25'b0000010110100010010000111;
    rom[40281] = 25'b0000010110100000011000001;
    rom[40282] = 25'b0000010110011110011111010;
    rom[40283] = 25'b0000010110011100100110011;
    rom[40284] = 25'b0000010110011010101101011;
    rom[40285] = 25'b0000010110011000110100011;
    rom[40286] = 25'b0000010110010110111011010;
    rom[40287] = 25'b0000010110010101000010001;
    rom[40288] = 25'b0000010110010011001000111;
    rom[40289] = 25'b0000010110010001001111100;
    rom[40290] = 25'b0000010110001111010110010;
    rom[40291] = 25'b0000010110001101011100110;
    rom[40292] = 25'b0000010110001011100011010;
    rom[40293] = 25'b0000010110001001101001101;
    rom[40294] = 25'b0000010110000111110000000;
    rom[40295] = 25'b0000010110000101110110010;
    rom[40296] = 25'b0000010110000011111100100;
    rom[40297] = 25'b0000010110000010000010101;
    rom[40298] = 25'b0000010110000000001000110;
    rom[40299] = 25'b0000010101111110001110110;
    rom[40300] = 25'b0000010101111100010100101;
    rom[40301] = 25'b0000010101111010011010101;
    rom[40302] = 25'b0000010101111000100000011;
    rom[40303] = 25'b0000010101110110100110001;
    rom[40304] = 25'b0000010101110100101011110;
    rom[40305] = 25'b0000010101110010110001011;
    rom[40306] = 25'b0000010101110000110111000;
    rom[40307] = 25'b0000010101101110111100100;
    rom[40308] = 25'b0000010101101101000001111;
    rom[40309] = 25'b0000010101101011000111010;
    rom[40310] = 25'b0000010101101001001100100;
    rom[40311] = 25'b0000010101100111010001110;
    rom[40312] = 25'b0000010101100101010110111;
    rom[40313] = 25'b0000010101100011011100000;
    rom[40314] = 25'b0000010101100001100001000;
    rom[40315] = 25'b0000010101011111100110000;
    rom[40316] = 25'b0000010101011101101011000;
    rom[40317] = 25'b0000010101011011101111110;
    rom[40318] = 25'b0000010101011001110100101;
    rom[40319] = 25'b0000010101010111111001010;
    rom[40320] = 25'b0000010101010101111110000;
    rom[40321] = 25'b0000010101010100000010100;
    rom[40322] = 25'b0000010101010010000111000;
    rom[40323] = 25'b0000010101010000001011100;
    rom[40324] = 25'b0000010101001110001111111;
    rom[40325] = 25'b0000010101001100010100010;
    rom[40326] = 25'b0000010101001010011000100;
    rom[40327] = 25'b0000010101001000011100111;
    rom[40328] = 25'b0000010101000110100001000;
    rom[40329] = 25'b0000010101000100100101000;
    rom[40330] = 25'b0000010101000010101001001;
    rom[40331] = 25'b0000010101000000101101001;
    rom[40332] = 25'b0000010100111110110001000;
    rom[40333] = 25'b0000010100111100110100111;
    rom[40334] = 25'b0000010100111010111000110;
    rom[40335] = 25'b0000010100111000111100011;
    rom[40336] = 25'b0000010100110111000000001;
    rom[40337] = 25'b0000010100110101000011110;
    rom[40338] = 25'b0000010100110011000111010;
    rom[40339] = 25'b0000010100110001001010110;
    rom[40340] = 25'b0000010100101111001110010;
    rom[40341] = 25'b0000010100101101010001101;
    rom[40342] = 25'b0000010100101011010100111;
    rom[40343] = 25'b0000010100101001011000010;
    rom[40344] = 25'b0000010100100111011011011;
    rom[40345] = 25'b0000010100100101011110101;
    rom[40346] = 25'b0000010100100011100001101;
    rom[40347] = 25'b0000010100100001100100110;
    rom[40348] = 25'b0000010100011111100111101;
    rom[40349] = 25'b0000010100011101101010101;
    rom[40350] = 25'b0000010100011011101101100;
    rom[40351] = 25'b0000010100011001110000011;
    rom[40352] = 25'b0000010100010111110011000;
    rom[40353] = 25'b0000010100010101110101110;
    rom[40354] = 25'b0000010100010011111000011;
    rom[40355] = 25'b0000010100010001111011000;
    rom[40356] = 25'b0000010100001111111101100;
    rom[40357] = 25'b0000010100001110000000000;
    rom[40358] = 25'b0000010100001100000010011;
    rom[40359] = 25'b0000010100001010000100110;
    rom[40360] = 25'b0000010100001000000111001;
    rom[40361] = 25'b0000010100000110001001010;
    rom[40362] = 25'b0000010100000100001011100;
    rom[40363] = 25'b0000010100000010001101110;
    rom[40364] = 25'b0000010100000000001111110;
    rom[40365] = 25'b0000010011111110010001111;
    rom[40366] = 25'b0000010011111100010011110;
    rom[40367] = 25'b0000010011111010010101110;
    rom[40368] = 25'b0000010011111000010111101;
    rom[40369] = 25'b0000010011110110011001100;
    rom[40370] = 25'b0000010011110100011011010;
    rom[40371] = 25'b0000010011110010011101000;
    rom[40372] = 25'b0000010011110000011110101;
    rom[40373] = 25'b0000010011101110100000010;
    rom[40374] = 25'b0000010011101100100001110;
    rom[40375] = 25'b0000010011101010100011011;
    rom[40376] = 25'b0000010011101000100100111;
    rom[40377] = 25'b0000010011100110100110010;
    rom[40378] = 25'b0000010011100100100111100;
    rom[40379] = 25'b0000010011100010101000111;
    rom[40380] = 25'b0000010011100000101010001;
    rom[40381] = 25'b0000010011011110101011010;
    rom[40382] = 25'b0000010011011100101100100;
    rom[40383] = 25'b0000010011011010101101100;
    rom[40384] = 25'b0000010011011000101110101;
    rom[40385] = 25'b0000010011010110101111101;
    rom[40386] = 25'b0000010011010100110000101;
    rom[40387] = 25'b0000010011010010110001100;
    rom[40388] = 25'b0000010011010000110010011;
    rom[40389] = 25'b0000010011001110110011001;
    rom[40390] = 25'b0000010011001100110100000;
    rom[40391] = 25'b0000010011001010110100101;
    rom[40392] = 25'b0000010011001000110101010;
    rom[40393] = 25'b0000010011000110110101111;
    rom[40394] = 25'b0000010011000100110110011;
    rom[40395] = 25'b0000010011000010110111000;
    rom[40396] = 25'b0000010011000000110111100;
    rom[40397] = 25'b0000010010111110110111111;
    rom[40398] = 25'b0000010010111100111000010;
    rom[40399] = 25'b0000010010111010111000101;
    rom[40400] = 25'b0000010010111000111000111;
    rom[40401] = 25'b0000010010110110111001001;
    rom[40402] = 25'b0000010010110100111001010;
    rom[40403] = 25'b0000010010110010111001011;
    rom[40404] = 25'b0000010010110000111001100;
    rom[40405] = 25'b0000010010101110111001100;
    rom[40406] = 25'b0000010010101100111001100;
    rom[40407] = 25'b0000010010101010111001100;
    rom[40408] = 25'b0000010010101000111001011;
    rom[40409] = 25'b0000010010100110111001010;
    rom[40410] = 25'b0000010010100100111001001;
    rom[40411] = 25'b0000010010100010111000111;
    rom[40412] = 25'b0000010010100000111000100;
    rom[40413] = 25'b0000010010011110111000010;
    rom[40414] = 25'b0000010010011100110111111;
    rom[40415] = 25'b0000010010011010110111100;
    rom[40416] = 25'b0000010010011000110111001;
    rom[40417] = 25'b0000010010010110110110101;
    rom[40418] = 25'b0000010010010100110110000;
    rom[40419] = 25'b0000010010010010110101011;
    rom[40420] = 25'b0000010010010000110100110;
    rom[40421] = 25'b0000010010001110110100001;
    rom[40422] = 25'b0000010010001100110011011;
    rom[40423] = 25'b0000010010001010110010101;
    rom[40424] = 25'b0000010010001000110001111;
    rom[40425] = 25'b0000010010000110110001001;
    rom[40426] = 25'b0000010010000100110000010;
    rom[40427] = 25'b0000010010000010101111010;
    rom[40428] = 25'b0000010010000000101110010;
    rom[40429] = 25'b0000010001111110101101011;
    rom[40430] = 25'b0000010001111100101100010;
    rom[40431] = 25'b0000010001111010101011010;
    rom[40432] = 25'b0000010001111000101010000;
    rom[40433] = 25'b0000010001110110101000111;
    rom[40434] = 25'b0000010001110100100111110;
    rom[40435] = 25'b0000010001110010100110100;
    rom[40436] = 25'b0000010001110000100101001;
    rom[40437] = 25'b0000010001101110100011110;
    rom[40438] = 25'b0000010001101100100010100;
    rom[40439] = 25'b0000010001101010100001000;
    rom[40440] = 25'b0000010001101000011111101;
    rom[40441] = 25'b0000010001100110011110001;
    rom[40442] = 25'b0000010001100100011100101;
    rom[40443] = 25'b0000010001100010011011000;
    rom[40444] = 25'b0000010001100000011001100;
    rom[40445] = 25'b0000010001011110010111110;
    rom[40446] = 25'b0000010001011100010110001;
    rom[40447] = 25'b0000010001011010010100011;
    rom[40448] = 25'b0000010001011000010010101;
    rom[40449] = 25'b0000010001010110010000111;
    rom[40450] = 25'b0000010001010100001111000;
    rom[40451] = 25'b0000010001010010001101010;
    rom[40452] = 25'b0000010001010000001011010;
    rom[40453] = 25'b0000010001001110001001010;
    rom[40454] = 25'b0000010001001100000111011;
    rom[40455] = 25'b0000010001001010000101010;
    rom[40456] = 25'b0000010001001000000011011;
    rom[40457] = 25'b0000010001000110000001010;
    rom[40458] = 25'b0000010001000011111111001;
    rom[40459] = 25'b0000010001000001111101000;
    rom[40460] = 25'b0000010000111111111010110;
    rom[40461] = 25'b0000010000111101111000100;
    rom[40462] = 25'b0000010000111011110110010;
    rom[40463] = 25'b0000010000111001110100000;
    rom[40464] = 25'b0000010000110111110001101;
    rom[40465] = 25'b0000010000110101101111010;
    rom[40466] = 25'b0000010000110011101100111;
    rom[40467] = 25'b0000010000110001101010100;
    rom[40468] = 25'b0000010000101111101000000;
    rom[40469] = 25'b0000010000101101100101100;
    rom[40470] = 25'b0000010000101011100010111;
    rom[40471] = 25'b0000010000101001100000011;
    rom[40472] = 25'b0000010000100111011101110;
    rom[40473] = 25'b0000010000100101011011001;
    rom[40474] = 25'b0000010000100011011000100;
    rom[40475] = 25'b0000010000100001010101110;
    rom[40476] = 25'b0000010000011111010011000;
    rom[40477] = 25'b0000010000011101010000010;
    rom[40478] = 25'b0000010000011011001101100;
    rom[40479] = 25'b0000010000011001001010110;
    rom[40480] = 25'b0000010000010111000111110;
    rom[40481] = 25'b0000010000010101000100111;
    rom[40482] = 25'b0000010000010011000010000;
    rom[40483] = 25'b0000010000010000111111000;
    rom[40484] = 25'b0000010000001110111100000;
    rom[40485] = 25'b0000010000001100111001000;
    rom[40486] = 25'b0000010000001010110110000;
    rom[40487] = 25'b0000010000001000110010111;
    rom[40488] = 25'b0000010000000110101111110;
    rom[40489] = 25'b0000010000000100101100101;
    rom[40490] = 25'b0000010000000010101001100;
    rom[40491] = 25'b0000010000000000100110011;
    rom[40492] = 25'b0000001111111110100011000;
    rom[40493] = 25'b0000001111111100011111111;
    rom[40494] = 25'b0000001111111010011100100;
    rom[40495] = 25'b0000001111111000011001010;
    rom[40496] = 25'b0000001111110110010101111;
    rom[40497] = 25'b0000001111110100010010100;
    rom[40498] = 25'b0000001111110010001111001;
    rom[40499] = 25'b0000001111110000001011110;
    rom[40500] = 25'b0000001111101110001000010;
    rom[40501] = 25'b0000001111101100000100110;
    rom[40502] = 25'b0000001111101010000001010;
    rom[40503] = 25'b0000001111100111111101110;
    rom[40504] = 25'b0000001111100101111010010;
    rom[40505] = 25'b0000001111100011110110101;
    rom[40506] = 25'b0000001111100001110011000;
    rom[40507] = 25'b0000001111011111101111011;
    rom[40508] = 25'b0000001111011101101011101;
    rom[40509] = 25'b0000001111011011101000000;
    rom[40510] = 25'b0000001111011001100100010;
    rom[40511] = 25'b0000001111010111100000100;
    rom[40512] = 25'b0000001111010101011100110;
    rom[40513] = 25'b0000001111010011011000111;
    rom[40514] = 25'b0000001111010001010101001;
    rom[40515] = 25'b0000001111001111010001010;
    rom[40516] = 25'b0000001111001101001101011;
    rom[40517] = 25'b0000001111001011001001100;
    rom[40518] = 25'b0000001111001001000101101;
    rom[40519] = 25'b0000001111000111000001101;
    rom[40520] = 25'b0000001111000100111101110;
    rom[40521] = 25'b0000001111000010111001101;
    rom[40522] = 25'b0000001111000000110101110;
    rom[40523] = 25'b0000001110111110110001101;
    rom[40524] = 25'b0000001110111100101101101;
    rom[40525] = 25'b0000001110111010101001100;
    rom[40526] = 25'b0000001110111000100101011;
    rom[40527] = 25'b0000001110110110100001010;
    rom[40528] = 25'b0000001110110100011101001;
    rom[40529] = 25'b0000001110110010011000111;
    rom[40530] = 25'b0000001110110000010100110;
    rom[40531] = 25'b0000001110101110010000100;
    rom[40532] = 25'b0000001110101100001100010;
    rom[40533] = 25'b0000001110101010001000000;
    rom[40534] = 25'b0000001110101000000011110;
    rom[40535] = 25'b0000001110100101111111011;
    rom[40536] = 25'b0000001110100011111011000;
    rom[40537] = 25'b0000001110100001110110110;
    rom[40538] = 25'b0000001110011111110010011;
    rom[40539] = 25'b0000001110011101101110000;
    rom[40540] = 25'b0000001110011011101001100;
    rom[40541] = 25'b0000001110011001100101001;
    rom[40542] = 25'b0000001110010111100000110;
    rom[40543] = 25'b0000001110010101011100010;
    rom[40544] = 25'b0000001110010011010111110;
    rom[40545] = 25'b0000001110010001010011010;
    rom[40546] = 25'b0000001110001111001110110;
    rom[40547] = 25'b0000001110001101001010010;
    rom[40548] = 25'b0000001110001011000101101;
    rom[40549] = 25'b0000001110001001000001000;
    rom[40550] = 25'b0000001110000110111100100;
    rom[40551] = 25'b0000001110000100110111110;
    rom[40552] = 25'b0000001110000010110011001;
    rom[40553] = 25'b0000001110000000101110100;
    rom[40554] = 25'b0000001101111110101001111;
    rom[40555] = 25'b0000001101111100100101001;
    rom[40556] = 25'b0000001101111010100000100;
    rom[40557] = 25'b0000001101111000011011110;
    rom[40558] = 25'b0000001101110110010111000;
    rom[40559] = 25'b0000001101110100010010010;
    rom[40560] = 25'b0000001101110010001101100;
    rom[40561] = 25'b0000001101110000001000101;
    rom[40562] = 25'b0000001101101110000011111;
    rom[40563] = 25'b0000001101101011111111000;
    rom[40564] = 25'b0000001101101001111010010;
    rom[40565] = 25'b0000001101100111110101011;
    rom[40566] = 25'b0000001101100101110000100;
    rom[40567] = 25'b0000001101100011101011101;
    rom[40568] = 25'b0000001101100001100110110;
    rom[40569] = 25'b0000001101011111100001111;
    rom[40570] = 25'b0000001101011101011100111;
    rom[40571] = 25'b0000001101011011011000000;
    rom[40572] = 25'b0000001101011001010011000;
    rom[40573] = 25'b0000001101010111001110000;
    rom[40574] = 25'b0000001101010101001001000;
    rom[40575] = 25'b0000001101010011000100000;
    rom[40576] = 25'b0000001101010000111111000;
    rom[40577] = 25'b0000001101001110111010000;
    rom[40578] = 25'b0000001101001100110101000;
    rom[40579] = 25'b0000001101001010101111111;
    rom[40580] = 25'b0000001101001000101010111;
    rom[40581] = 25'b0000001101000110100101110;
    rom[40582] = 25'b0000001101000100100000101;
    rom[40583] = 25'b0000001101000010011011101;
    rom[40584] = 25'b0000001101000000010110100;
    rom[40585] = 25'b0000001100111110010001011;
    rom[40586] = 25'b0000001100111100001100001;
    rom[40587] = 25'b0000001100111010000111001;
    rom[40588] = 25'b0000001100111000000001111;
    rom[40589] = 25'b0000001100110101111100110;
    rom[40590] = 25'b0000001100110011110111101;
    rom[40591] = 25'b0000001100110001110010011;
    rom[40592] = 25'b0000001100101111101101001;
    rom[40593] = 25'b0000001100101101101000000;
    rom[40594] = 25'b0000001100101011100010110;
    rom[40595] = 25'b0000001100101001011101100;
    rom[40596] = 25'b0000001100100111011000010;
    rom[40597] = 25'b0000001100100101010011000;
    rom[40598] = 25'b0000001100100011001101110;
    rom[40599] = 25'b0000001100100001001000100;
    rom[40600] = 25'b0000001100011111000011010;
    rom[40601] = 25'b0000001100011100111101111;
    rom[40602] = 25'b0000001100011010111000101;
    rom[40603] = 25'b0000001100011000110011011;
    rom[40604] = 25'b0000001100010110101110000;
    rom[40605] = 25'b0000001100010100101000101;
    rom[40606] = 25'b0000001100010010100011011;
    rom[40607] = 25'b0000001100010000011110000;
    rom[40608] = 25'b0000001100001110011000101;
    rom[40609] = 25'b0000001100001100010011010;
    rom[40610] = 25'b0000001100001010001110000;
    rom[40611] = 25'b0000001100001000001000101;
    rom[40612] = 25'b0000001100000110000011010;
    rom[40613] = 25'b0000001100000011111101111;
    rom[40614] = 25'b0000001100000001111000011;
    rom[40615] = 25'b0000001011111111110011001;
    rom[40616] = 25'b0000001011111101101101110;
    rom[40617] = 25'b0000001011111011101000010;
    rom[40618] = 25'b0000001011111001100010110;
    rom[40619] = 25'b0000001011110111011101100;
    rom[40620] = 25'b0000001011110101011000000;
    rom[40621] = 25'b0000001011110011010010100;
    rom[40622] = 25'b0000001011110001001101010;
    rom[40623] = 25'b0000001011101111000111110;
    rom[40624] = 25'b0000001011101101000010010;
    rom[40625] = 25'b0000001011101010111100111;
    rom[40626] = 25'b0000001011101000110111011;
    rom[40627] = 25'b0000001011100110110010000;
    rom[40628] = 25'b0000001011100100101100100;
    rom[40629] = 25'b0000001011100010100111000;
    rom[40630] = 25'b0000001011100000100001101;
    rom[40631] = 25'b0000001011011110011100000;
    rom[40632] = 25'b0000001011011100010110101;
    rom[40633] = 25'b0000001011011010010001001;
    rom[40634] = 25'b0000001011011000001011110;
    rom[40635] = 25'b0000001011010110000110001;
    rom[40636] = 25'b0000001011010100000000110;
    rom[40637] = 25'b0000001011010001111011010;
    rom[40638] = 25'b0000001011001111110101110;
    rom[40639] = 25'b0000001011001101110000010;
    rom[40640] = 25'b0000001011001011101010110;
    rom[40641] = 25'b0000001011001001100101010;
    rom[40642] = 25'b0000001011000111011111111;
    rom[40643] = 25'b0000001011000101011010010;
    rom[40644] = 25'b0000001011000011010100111;
    rom[40645] = 25'b0000001011000001001111010;
    rom[40646] = 25'b0000001010111111001001111;
    rom[40647] = 25'b0000001010111101000100010;
    rom[40648] = 25'b0000001010111010111110111;
    rom[40649] = 25'b0000001010111000111001010;
    rom[40650] = 25'b0000001010110110110011111;
    rom[40651] = 25'b0000001010110100101110010;
    rom[40652] = 25'b0000001010110010101000111;
    rom[40653] = 25'b0000001010110000100011010;
    rom[40654] = 25'b0000001010101110011101111;
    rom[40655] = 25'b0000001010101100011000011;
    rom[40656] = 25'b0000001010101010010010111;
    rom[40657] = 25'b0000001010101000001101011;
    rom[40658] = 25'b0000001010100110000111111;
    rom[40659] = 25'b0000001010100100000010011;
    rom[40660] = 25'b0000001010100001111100111;
    rom[40661] = 25'b0000001010011111110111011;
    rom[40662] = 25'b0000001010011101110010000;
    rom[40663] = 25'b0000001010011011101100011;
    rom[40664] = 25'b0000001010011001100111000;
    rom[40665] = 25'b0000001010010111100001100;
    rom[40666] = 25'b0000001010010101011100000;
    rom[40667] = 25'b0000001010010011010110100;
    rom[40668] = 25'b0000001010010001010001001;
    rom[40669] = 25'b0000001010001111001011101;
    rom[40670] = 25'b0000001010001101000110010;
    rom[40671] = 25'b0000001010001011000000110;
    rom[40672] = 25'b0000001010001000111011010;
    rom[40673] = 25'b0000001010000110110101111;
    rom[40674] = 25'b0000001010000100110000011;
    rom[40675] = 25'b0000001010000010101011000;
    rom[40676] = 25'b0000001010000000100101101;
    rom[40677] = 25'b0000001001111110100000001;
    rom[40678] = 25'b0000001001111100011010101;
    rom[40679] = 25'b0000001001111010010101011;
    rom[40680] = 25'b0000001001111000001111111;
    rom[40681] = 25'b0000001001110110001010011;
    rom[40682] = 25'b0000001001110100000101001;
    rom[40683] = 25'b0000001001110001111111110;
    rom[40684] = 25'b0000001001101111111010010;
    rom[40685] = 25'b0000001001101101110100111;
    rom[40686] = 25'b0000001001101011101111100;
    rom[40687] = 25'b0000001001101001101010010;
    rom[40688] = 25'b0000001001100111100100111;
    rom[40689] = 25'b0000001001100101011111100;
    rom[40690] = 25'b0000001001100011011010001;
    rom[40691] = 25'b0000001001100001010100110;
    rom[40692] = 25'b0000001001011111001111011;
    rom[40693] = 25'b0000001001011101001010001;
    rom[40694] = 25'b0000001001011011000100110;
    rom[40695] = 25'b0000001001011000111111100;
    rom[40696] = 25'b0000001001010110111010001;
    rom[40697] = 25'b0000001001010100110100111;
    rom[40698] = 25'b0000001001010010101111101;
    rom[40699] = 25'b0000001001010000101010011;
    rom[40700] = 25'b0000001001001110100101001;
    rom[40701] = 25'b0000001001001100011111111;
    rom[40702] = 25'b0000001001001010011010101;
    rom[40703] = 25'b0000001001001000010101011;
    rom[40704] = 25'b0000001001000110010000001;
    rom[40705] = 25'b0000001001000100001011000;
    rom[40706] = 25'b0000001001000010000101110;
    rom[40707] = 25'b0000001001000000000000100;
    rom[40708] = 25'b0000001000111101111011011;
    rom[40709] = 25'b0000001000111011110110010;
    rom[40710] = 25'b0000001000111001110001000;
    rom[40711] = 25'b0000001000110111101011111;
    rom[40712] = 25'b0000001000110101100110110;
    rom[40713] = 25'b0000001000110011100001101;
    rom[40714] = 25'b0000001000110001011100100;
    rom[40715] = 25'b0000001000101111010111011;
    rom[40716] = 25'b0000001000101101010010010;
    rom[40717] = 25'b0000001000101011001101010;
    rom[40718] = 25'b0000001000101001001000001;
    rom[40719] = 25'b0000001000100111000011001;
    rom[40720] = 25'b0000001000100100111110000;
    rom[40721] = 25'b0000001000100010111001000;
    rom[40722] = 25'b0000001000100000110100000;
    rom[40723] = 25'b0000001000011110101111000;
    rom[40724] = 25'b0000001000011100101010000;
    rom[40725] = 25'b0000001000011010100101000;
    rom[40726] = 25'b0000001000011000100000000;
    rom[40727] = 25'b0000001000010110011011001;
    rom[40728] = 25'b0000001000010100010110001;
    rom[40729] = 25'b0000001000010010010001010;
    rom[40730] = 25'b0000001000010000001100011;
    rom[40731] = 25'b0000001000001110000111100;
    rom[40732] = 25'b0000001000001100000010101;
    rom[40733] = 25'b0000001000001001111101110;
    rom[40734] = 25'b0000001000000111111000110;
    rom[40735] = 25'b0000001000000101110100000;
    rom[40736] = 25'b0000001000000011101111010;
    rom[40737] = 25'b0000001000000001101010011;
    rom[40738] = 25'b0000000111111111100101101;
    rom[40739] = 25'b0000000111111101100000111;
    rom[40740] = 25'b0000000111111011011100000;
    rom[40741] = 25'b0000000111111001010111011;
    rom[40742] = 25'b0000000111110111010010101;
    rom[40743] = 25'b0000000111110101001101111;
    rom[40744] = 25'b0000000111110011001001010;
    rom[40745] = 25'b0000000111110001000100100;
    rom[40746] = 25'b0000000111101110111111111;
    rom[40747] = 25'b0000000111101100111011010;
    rom[40748] = 25'b0000000111101010110110101;
    rom[40749] = 25'b0000000111101000110010000;
    rom[40750] = 25'b0000000111100110101101100;
    rom[40751] = 25'b0000000111100100101000111;
    rom[40752] = 25'b0000000111100010100100011;
    rom[40753] = 25'b0000000111100000011111110;
    rom[40754] = 25'b0000000111011110011011010;
    rom[40755] = 25'b0000000111011100010110110;
    rom[40756] = 25'b0000000111011010010010010;
    rom[40757] = 25'b0000000111011000001101111;
    rom[40758] = 25'b0000000111010110001001011;
    rom[40759] = 25'b0000000111010100000101000;
    rom[40760] = 25'b0000000111010010000000101;
    rom[40761] = 25'b0000000111001111111100001;
    rom[40762] = 25'b0000000111001101110111111;
    rom[40763] = 25'b0000000111001011110011100;
    rom[40764] = 25'b0000000111001001101111001;
    rom[40765] = 25'b0000000111000111101010111;
    rom[40766] = 25'b0000000111000101100110101;
    rom[40767] = 25'b0000000111000011100010010;
    rom[40768] = 25'b0000000111000001011110000;
    rom[40769] = 25'b0000000110111111011001111;
    rom[40770] = 25'b0000000110111101010101101;
    rom[40771] = 25'b0000000110111011010001100;
    rom[40772] = 25'b0000000110111001001101011;
    rom[40773] = 25'b0000000110110111001001010;
    rom[40774] = 25'b0000000110110101000101001;
    rom[40775] = 25'b0000000110110011000001000;
    rom[40776] = 25'b0000000110110000111101000;
    rom[40777] = 25'b0000000110101110111000111;
    rom[40778] = 25'b0000000110101100110100111;
    rom[40779] = 25'b0000000110101010110000111;
    rom[40780] = 25'b0000000110101000101100111;
    rom[40781] = 25'b0000000110100110101000111;
    rom[40782] = 25'b0000000110100100100101001;
    rom[40783] = 25'b0000000110100010100001001;
    rom[40784] = 25'b0000000110100000011101010;
    rom[40785] = 25'b0000000110011110011001011;
    rom[40786] = 25'b0000000110011100010101100;
    rom[40787] = 25'b0000000110011010010001110;
    rom[40788] = 25'b0000000110011000001110000;
    rom[40789] = 25'b0000000110010110001010010;
    rom[40790] = 25'b0000000110010100000110100;
    rom[40791] = 25'b0000000110010010000010110;
    rom[40792] = 25'b0000000110001111111111001;
    rom[40793] = 25'b0000000110001101111011011;
    rom[40794] = 25'b0000000110001011110111110;
    rom[40795] = 25'b0000000110001001110100001;
    rom[40796] = 25'b0000000110000111110000101;
    rom[40797] = 25'b0000000110000101101101000;
    rom[40798] = 25'b0000000110000011101001011;
    rom[40799] = 25'b0000000110000001100101111;
    rom[40800] = 25'b0000000101111111100010011;
    rom[40801] = 25'b0000000101111101011111000;
    rom[40802] = 25'b0000000101111011011011100;
    rom[40803] = 25'b0000000101111001011000001;
    rom[40804] = 25'b0000000101110111010100110;
    rom[40805] = 25'b0000000101110101010001100;
    rom[40806] = 25'b0000000101110011001110001;
    rom[40807] = 25'b0000000101110001001010111;
    rom[40808] = 25'b0000000101101111000111100;
    rom[40809] = 25'b0000000101101101000100011;
    rom[40810] = 25'b0000000101101011000001001;
    rom[40811] = 25'b0000000101101000111101111;
    rom[40812] = 25'b0000000101100110111010110;
    rom[40813] = 25'b0000000101100100110111101;
    rom[40814] = 25'b0000000101100010110100101;
    rom[40815] = 25'b0000000101100000110001100;
    rom[40816] = 25'b0000000101011110101110100;
    rom[40817] = 25'b0000000101011100101011011;
    rom[40818] = 25'b0000000101011010101000011;
    rom[40819] = 25'b0000000101011000100101100;
    rom[40820] = 25'b0000000101010110100010100;
    rom[40821] = 25'b0000000101010100011111110;
    rom[40822] = 25'b0000000101010010011100110;
    rom[40823] = 25'b0000000101010000011010000;
    rom[40824] = 25'b0000000101001110010111010;
    rom[40825] = 25'b0000000101001100010100011;
    rom[40826] = 25'b0000000101001010010001101;
    rom[40827] = 25'b0000000101001000001111000;
    rom[40828] = 25'b0000000101000110001100010;
    rom[40829] = 25'b0000000101000100001001101;
    rom[40830] = 25'b0000000101000010000111000;
    rom[40831] = 25'b0000000101000000000100011;
    rom[40832] = 25'b0000000100111110000001111;
    rom[40833] = 25'b0000000100111011111111010;
    rom[40834] = 25'b0000000100111001111100110;
    rom[40835] = 25'b0000000100110111111010011;
    rom[40836] = 25'b0000000100110101111000000;
    rom[40837] = 25'b0000000100110011110101100;
    rom[40838] = 25'b0000000100110001110011001;
    rom[40839] = 25'b0000000100101111110000111;
    rom[40840] = 25'b0000000100101101101110100;
    rom[40841] = 25'b0000000100101011101100010;
    rom[40842] = 25'b0000000100101001101010000;
    rom[40843] = 25'b0000000100100111100111111;
    rom[40844] = 25'b0000000100100101100101101;
    rom[40845] = 25'b0000000100100011100011100;
    rom[40846] = 25'b0000000100100001100001011;
    rom[40847] = 25'b0000000100011111011111011;
    rom[40848] = 25'b0000000100011101011101011;
    rom[40849] = 25'b0000000100011011011011011;
    rom[40850] = 25'b0000000100011001011001011;
    rom[40851] = 25'b0000000100010111010111100;
    rom[40852] = 25'b0000000100010101010101100;
    rom[40853] = 25'b0000000100010011010011110;
    rom[40854] = 25'b0000000100010001010001111;
    rom[40855] = 25'b0000000100001111010000001;
    rom[40856] = 25'b0000000100001101001110010;
    rom[40857] = 25'b0000000100001011001100101;
    rom[40858] = 25'b0000000100001001001011000;
    rom[40859] = 25'b0000000100000111001001010;
    rom[40860] = 25'b0000000100000101000111110;
    rom[40861] = 25'b0000000100000011000110001;
    rom[40862] = 25'b0000000100000001000100101;
    rom[40863] = 25'b0000000011111111000011000;
    rom[40864] = 25'b0000000011111101000001101;
    rom[40865] = 25'b0000000011111011000000001;
    rom[40866] = 25'b0000000011111000111110110;
    rom[40867] = 25'b0000000011110110111101011;
    rom[40868] = 25'b0000000011110100111100001;
    rom[40869] = 25'b0000000011110010111010111;
    rom[40870] = 25'b0000000011110000111001101;
    rom[40871] = 25'b0000000011101110111000011;
    rom[40872] = 25'b0000000011101100110111010;
    rom[40873] = 25'b0000000011101010110110001;
    rom[40874] = 25'b0000000011101000110101000;
    rom[40875] = 25'b0000000011100110110100000;
    rom[40876] = 25'b0000000011100100110010111;
    rom[40877] = 25'b0000000011100010110010000;
    rom[40878] = 25'b0000000011100000110001001;
    rom[40879] = 25'b0000000011011110110000001;
    rom[40880] = 25'b0000000011011100101111010;
    rom[40881] = 25'b0000000011011010101110100;
    rom[40882] = 25'b0000000011011000101101101;
    rom[40883] = 25'b0000000011010110101101000;
    rom[40884] = 25'b0000000011010100101100010;
    rom[40885] = 25'b0000000011010010101011101;
    rom[40886] = 25'b0000000011010000101010111;
    rom[40887] = 25'b0000000011001110101010011;
    rom[40888] = 25'b0000000011001100101001111;
    rom[40889] = 25'b0000000011001010101001011;
    rom[40890] = 25'b0000000011001000101000111;
    rom[40891] = 25'b0000000011000110101000100;
    rom[40892] = 25'b0000000011000100101000001;
    rom[40893] = 25'b0000000011000010100111110;
    rom[40894] = 25'b0000000011000000100111100;
    rom[40895] = 25'b0000000010111110100111010;
    rom[40896] = 25'b0000000010111100100111000;
    rom[40897] = 25'b0000000010111010100110111;
    rom[40898] = 25'b0000000010111000100110110;
    rom[40899] = 25'b0000000010110110100110101;
    rom[40900] = 25'b0000000010110100100110101;
    rom[40901] = 25'b0000000010110010100110101;
    rom[40902] = 25'b0000000010110000100110101;
    rom[40903] = 25'b0000000010101110100110110;
    rom[40904] = 25'b0000000010101100100110111;
    rom[40905] = 25'b0000000010101010100111000;
    rom[40906] = 25'b0000000010101000100111010;
    rom[40907] = 25'b0000000010100110100111100;
    rom[40908] = 25'b0000000010100100100111111;
    rom[40909] = 25'b0000000010100010101000010;
    rom[40910] = 25'b0000000010100000101000100;
    rom[40911] = 25'b0000000010011110101001000;
    rom[40912] = 25'b0000000010011100101001100;
    rom[40913] = 25'b0000000010011010101010000;
    rom[40914] = 25'b0000000010011000101010100;
    rom[40915] = 25'b0000000010010110101011001;
    rom[40916] = 25'b0000000010010100101011111;
    rom[40917] = 25'b0000000010010010101100100;
    rom[40918] = 25'b0000000010010000101101011;
    rom[40919] = 25'b0000000010001110101110001;
    rom[40920] = 25'b0000000010001100101110111;
    rom[40921] = 25'b0000000010001010101111111;
    rom[40922] = 25'b0000000010001000110000110;
    rom[40923] = 25'b0000000010000110110001110;
    rom[40924] = 25'b0000000010000100110010110;
    rom[40925] = 25'b0000000010000010110011110;
    rom[40926] = 25'b0000000010000000110100111;
    rom[40927] = 25'b0000000001111110110110001;
    rom[40928] = 25'b0000000001111100110111010;
    rom[40929] = 25'b0000000001111010111000100;
    rom[40930] = 25'b0000000001111000111001110;
    rom[40931] = 25'b0000000001110110111011001;
    rom[40932] = 25'b0000000001110100111100100;
    rom[40933] = 25'b0000000001110010111110000;
    rom[40934] = 25'b0000000001110000111111100;
    rom[40935] = 25'b0000000001101111000001000;
    rom[40936] = 25'b0000000001101101000010101;
    rom[40937] = 25'b0000000001101011000100010;
    rom[40938] = 25'b0000000001101001000110000;
    rom[40939] = 25'b0000000001100111000111101;
    rom[40940] = 25'b0000000001100101001001011;
    rom[40941] = 25'b0000000001100011001011010;
    rom[40942] = 25'b0000000001100001001101001;
    rom[40943] = 25'b0000000001011111001111000;
    rom[40944] = 25'b0000000001011101010001000;
    rom[40945] = 25'b0000000001011011010011001;
    rom[40946] = 25'b0000000001011001010101001;
    rom[40947] = 25'b0000000001010111010111010;
    rom[40948] = 25'b0000000001010101011001011;
    rom[40949] = 25'b0000000001010011011011101;
    rom[40950] = 25'b0000000001010001011101111;
    rom[40951] = 25'b0000000001001111100000010;
    rom[40952] = 25'b0000000001001101100010100;
    rom[40953] = 25'b0000000001001011100101000;
    rom[40954] = 25'b0000000001001001100111011;
    rom[40955] = 25'b0000000001000111101010000;
    rom[40956] = 25'b0000000001000101101100101;
    rom[40957] = 25'b0000000001000011101111001;
    rom[40958] = 25'b0000000001000001110001111;
    rom[40959] = 25'b0000000000111111110100100;
    rom[40960] = 25'b0000000000111101110111011;
    rom[40961] = 25'b0000000000111011111010001;
    rom[40962] = 25'b0000000000111001111101000;
    rom[40963] = 25'b0000000000111000000000000;
    rom[40964] = 25'b0000000000110110000010111;
    rom[40965] = 25'b0000000000110100000110000;
    rom[40966] = 25'b0000000000110010001001001;
    rom[40967] = 25'b0000000000110000001100010;
    rom[40968] = 25'b0000000000101110001111011;
    rom[40969] = 25'b0000000000101100010010101;
    rom[40970] = 25'b0000000000101010010101111;
    rom[40971] = 25'b0000000000101000011001010;
    rom[40972] = 25'b0000000000100110011100101;
    rom[40973] = 25'b0000000000100100100000001;
    rom[40974] = 25'b0000000000100010100011101;
    rom[40975] = 25'b0000000000100000100111010;
    rom[40976] = 25'b0000000000011110101010111;
    rom[40977] = 25'b0000000000011100101110100;
    rom[40978] = 25'b0000000000011010110010010;
    rom[40979] = 25'b0000000000011000110110000;
    rom[40980] = 25'b0000000000010110111001111;
    rom[40981] = 25'b0000000000010100111101110;
    rom[40982] = 25'b0000000000010011000001101;
    rom[40983] = 25'b0000000000010001000101101;
    rom[40984] = 25'b0000000000001111001001101;
    rom[40985] = 25'b0000000000001101001101110;
    rom[40986] = 25'b0000000000001011010001111;
    rom[40987] = 25'b0000000000001001010110001;
    rom[40988] = 25'b0000000000000111011010011;
    rom[40989] = 25'b0000000000000101011110110;
    rom[40990] = 25'b0000000000000011100011001;
    rom[40991] = 25'b0000000000000001100111101;
    rom[40992] = 25'b1111111111111111101100001;
    rom[40993] = 25'b1111111111111101110000101;
    rom[40994] = 25'b1111111111111011110101011;
    rom[40995] = 25'b1111111111111001111010000;
    rom[40996] = 25'b1111111111110111111110101;
    rom[40997] = 25'b1111111111110110000011100;
    rom[40998] = 25'b1111111111110100001000011;
    rom[40999] = 25'b1111111111110010001101001;
    rom[41000] = 25'b1111111111110000010010001;
    rom[41001] = 25'b1111111111101110010111001;
    rom[41002] = 25'b1111111111101100011100001;
    rom[41003] = 25'b1111111111101010100001010;
    rom[41004] = 25'b1111111111101000100110100;
    rom[41005] = 25'b1111111111100110101011110;
    rom[41006] = 25'b1111111111100100110001000;
    rom[41007] = 25'b1111111111100010110110011;
    rom[41008] = 25'b1111111111100000111011111;
    rom[41009] = 25'b1111111111011111000001010;
    rom[41010] = 25'b1111111111011101000110110;
    rom[41011] = 25'b1111111111011011001100011;
    rom[41012] = 25'b1111111111011001010010000;
    rom[41013] = 25'b1111111111010111010111101;
    rom[41014] = 25'b1111111111010101011101011;
    rom[41015] = 25'b1111111111010011100011010;
    rom[41016] = 25'b1111111111010001101001001;
    rom[41017] = 25'b1111111111001111101111001;
    rom[41018] = 25'b1111111111001101110101001;
    rom[41019] = 25'b1111111111001011111011001;
    rom[41020] = 25'b1111111111001010000001010;
    rom[41021] = 25'b1111111111001000000111011;
    rom[41022] = 25'b1111111111000110001101110;
    rom[41023] = 25'b1111111111000100010100000;
    rom[41024] = 25'b1111111111000010011010011;
    rom[41025] = 25'b1111111111000000100000110;
    rom[41026] = 25'b1111111110111110100111010;
    rom[41027] = 25'b1111111110111100101101110;
    rom[41028] = 25'b1111111110111010110100011;
    rom[41029] = 25'b1111111110111000111011000;
    rom[41030] = 25'b1111111110110111000001110;
    rom[41031] = 25'b1111111110110101001000100;
    rom[41032] = 25'b1111111110110011001111011;
    rom[41033] = 25'b1111111110110001010110010;
    rom[41034] = 25'b1111111110101111011101010;
    rom[41035] = 25'b1111111110101101100100011;
    rom[41036] = 25'b1111111110101011101011011;
    rom[41037] = 25'b1111111110101001110010100;
    rom[41038] = 25'b1111111110100111111001110;
    rom[41039] = 25'b1111111110100110000001000;
    rom[41040] = 25'b1111111110100100001000011;
    rom[41041] = 25'b1111111110100010001111111;
    rom[41042] = 25'b1111111110100000010111010;
    rom[41043] = 25'b1111111110011110011110110;
    rom[41044] = 25'b1111111110011100100110011;
    rom[41045] = 25'b1111111110011010101110000;
    rom[41046] = 25'b1111111110011000110101110;
    rom[41047] = 25'b1111111110010110111101101;
    rom[41048] = 25'b1111111110010101000101100;
    rom[41049] = 25'b1111111110010011001101011;
    rom[41050] = 25'b1111111110010001010101010;
    rom[41051] = 25'b1111111110001111011101011;
    rom[41052] = 25'b1111111110001101100101100;
    rom[41053] = 25'b1111111110001011101101101;
    rom[41054] = 25'b1111111110001001110101111;
    rom[41055] = 25'b1111111110000111111110010;
    rom[41056] = 25'b1111111110000110000110101;
    rom[41057] = 25'b1111111110000100001111000;
    rom[41058] = 25'b1111111110000010010111100;
    rom[41059] = 25'b1111111110000000100000000;
    rom[41060] = 25'b1111111101111110101000101;
    rom[41061] = 25'b1111111101111100110001011;
    rom[41062] = 25'b1111111101111010111010001;
    rom[41063] = 25'b1111111101111001000011000;
    rom[41064] = 25'b1111111101110111001011110;
    rom[41065] = 25'b1111111101110101010100110;
    rom[41066] = 25'b1111111101110011011101110;
    rom[41067] = 25'b1111111101110001100110111;
    rom[41068] = 25'b1111111101101111110000000;
    rom[41069] = 25'b1111111101101101111001010;
    rom[41070] = 25'b1111111101101100000010100;
    rom[41071] = 25'b1111111101101010001011111;
    rom[41072] = 25'b1111111101101000010101010;
    rom[41073] = 25'b1111111101100110011110110;
    rom[41074] = 25'b1111111101100100101000011;
    rom[41075] = 25'b1111111101100010110010000;
    rom[41076] = 25'b1111111101100000111011101;
    rom[41077] = 25'b1111111101011111000101011;
    rom[41078] = 25'b1111111101011101001111001;
    rom[41079] = 25'b1111111101011011011001001;
    rom[41080] = 25'b1111111101011001100011001;
    rom[41081] = 25'b1111111101010111101101000;
    rom[41082] = 25'b1111111101010101110111010;
    rom[41083] = 25'b1111111101010100000001011;
    rom[41084] = 25'b1111111101010010001011101;
    rom[41085] = 25'b1111111101010000010101111;
    rom[41086] = 25'b1111111101001110100000010;
    rom[41087] = 25'b1111111101001100101010101;
    rom[41088] = 25'b1111111101001010110101010;
    rom[41089] = 25'b1111111101001000111111110;
    rom[41090] = 25'b1111111101000111001010011;
    rom[41091] = 25'b1111111101000101010101001;
    rom[41092] = 25'b1111111101000011011111111;
    rom[41093] = 25'b1111111101000001101010111;
    rom[41094] = 25'b1111111100111111110101110;
    rom[41095] = 25'b1111111100111110000000110;
    rom[41096] = 25'b1111111100111100001011110;
    rom[41097] = 25'b1111111100111010010110111;
    rom[41098] = 25'b1111111100111000100010001;
    rom[41099] = 25'b1111111100110110101101011;
    rom[41100] = 25'b1111111100110100111000110;
    rom[41101] = 25'b1111111100110011000100001;
    rom[41102] = 25'b1111111100110001001111101;
    rom[41103] = 25'b1111111100101111011011010;
    rom[41104] = 25'b1111111100101101100110111;
    rom[41105] = 25'b1111111100101011110010100;
    rom[41106] = 25'b1111111100101001111110010;
    rom[41107] = 25'b1111111100101000001010001;
    rom[41108] = 25'b1111111100100110010110000;
    rom[41109] = 25'b1111111100100100100010000;
    rom[41110] = 25'b1111111100100010101110001;
    rom[41111] = 25'b1111111100100000111010001;
    rom[41112] = 25'b1111111100011111000110011;
    rom[41113] = 25'b1111111100011101010010101;
    rom[41114] = 25'b1111111100011011011111000;
    rom[41115] = 25'b1111111100011001101011100;
    rom[41116] = 25'b1111111100010111110111111;
    rom[41117] = 25'b1111111100010110000100100;
    rom[41118] = 25'b1111111100010100010001001;
    rom[41119] = 25'b1111111100010010011101111;
    rom[41120] = 25'b1111111100010000101010101;
    rom[41121] = 25'b1111111100001110110111100;
    rom[41122] = 25'b1111111100001101000100011;
    rom[41123] = 25'b1111111100001011010001011;
    rom[41124] = 25'b1111111100001001011110100;
    rom[41125] = 25'b1111111100000111101011101;
    rom[41126] = 25'b1111111100000101111000111;
    rom[41127] = 25'b1111111100000100000110001;
    rom[41128] = 25'b1111111100000010010011100;
    rom[41129] = 25'b1111111100000000100001000;
    rom[41130] = 25'b1111111011111110101110100;
    rom[41131] = 25'b1111111011111100111100001;
    rom[41132] = 25'b1111111011111011001001110;
    rom[41133] = 25'b1111111011111001010111100;
    rom[41134] = 25'b1111111011110111100101010;
    rom[41135] = 25'b1111111011110101110011001;
    rom[41136] = 25'b1111111011110100000001001;
    rom[41137] = 25'b1111111011110010001111010;
    rom[41138] = 25'b1111111011110000011101010;
    rom[41139] = 25'b1111111011101110101011100;
    rom[41140] = 25'b1111111011101100111001110;
    rom[41141] = 25'b1111111011101011001000001;
    rom[41142] = 25'b1111111011101001010110101;
    rom[41143] = 25'b1111111011100111100101000;
    rom[41144] = 25'b1111111011100101110011100;
    rom[41145] = 25'b1111111011100100000010010;
    rom[41146] = 25'b1111111011100010010001000;
    rom[41147] = 25'b1111111011100000011111110;
    rom[41148] = 25'b1111111011011110101110101;
    rom[41149] = 25'b1111111011011100111101101;
    rom[41150] = 25'b1111111011011011001100101;
    rom[41151] = 25'b1111111011011001011011110;
    rom[41152] = 25'b1111111011010111101010111;
    rom[41153] = 25'b1111111011010101111010001;
    rom[41154] = 25'b1111111011010100001001100;
    rom[41155] = 25'b1111111011010010011000111;
    rom[41156] = 25'b1111111011010000101000011;
    rom[41157] = 25'b1111111011001110111000000;
    rom[41158] = 25'b1111111011001101000111101;
    rom[41159] = 25'b1111111011001011010111011;
    rom[41160] = 25'b1111111011001001100111001;
    rom[41161] = 25'b1111111011000111110111000;
    rom[41162] = 25'b1111111011000110000111000;
    rom[41163] = 25'b1111111011000100010111000;
    rom[41164] = 25'b1111111011000010100111001;
    rom[41165] = 25'b1111111011000000110111011;
    rom[41166] = 25'b1111111010111111000111101;
    rom[41167] = 25'b1111111010111101011000000;
    rom[41168] = 25'b1111111010111011101000011;
    rom[41169] = 25'b1111111010111001111000111;
    rom[41170] = 25'b1111111010111000001001100;
    rom[41171] = 25'b1111111010110110011010001;
    rom[41172] = 25'b1111111010110100101010111;
    rom[41173] = 25'b1111111010110010111011110;
    rom[41174] = 25'b1111111010110001001100101;
    rom[41175] = 25'b1111111010101111011101101;
    rom[41176] = 25'b1111111010101101101110101;
    rom[41177] = 25'b1111111010101011111111111;
    rom[41178] = 25'b1111111010101010010001000;
    rom[41179] = 25'b1111111010101000100010011;
    rom[41180] = 25'b1111111010100110110011101;
    rom[41181] = 25'b1111111010100101000101001;
    rom[41182] = 25'b1111111010100011010110110;
    rom[41183] = 25'b1111111010100001101000011;
    rom[41184] = 25'b1111111010011111111010000;
    rom[41185] = 25'b1111111010011110001011111;
    rom[41186] = 25'b1111111010011100011101110;
    rom[41187] = 25'b1111111010011010101111101;
    rom[41188] = 25'b1111111010011001000001101;
    rom[41189] = 25'b1111111010010111010011110;
    rom[41190] = 25'b1111111010010101100110000;
    rom[41191] = 25'b1111111010010011111000010;
    rom[41192] = 25'b1111111010010010001010101;
    rom[41193] = 25'b1111111010010000011101000;
    rom[41194] = 25'b1111111010001110101111100;
    rom[41195] = 25'b1111111010001101000010001;
    rom[41196] = 25'b1111111010001011010100110;
    rom[41197] = 25'b1111111010001001100111100;
    rom[41198] = 25'b1111111010000111111010100;
    rom[41199] = 25'b1111111010000110001101011;
    rom[41200] = 25'b1111111010000100100000010;
    rom[41201] = 25'b1111111010000010110011011;
    rom[41202] = 25'b1111111010000001000110101;
    rom[41203] = 25'b1111111001111111011001111;
    rom[41204] = 25'b1111111001111101101101010;
    rom[41205] = 25'b1111111001111100000000101;
    rom[41206] = 25'b1111111001111010010100001;
    rom[41207] = 25'b1111111001111000100111110;
    rom[41208] = 25'b1111111001110110111011011;
    rom[41209] = 25'b1111111001110101001111010;
    rom[41210] = 25'b1111111001110011100011000;
    rom[41211] = 25'b1111111001110001110110111;
    rom[41212] = 25'b1111111001110000001011000;
    rom[41213] = 25'b1111111001101110011111000;
    rom[41214] = 25'b1111111001101100110011010;
    rom[41215] = 25'b1111111001101011000111100;
    rom[41216] = 25'b1111111001101001011011110;
    rom[41217] = 25'b1111111001100111110000010;
    rom[41218] = 25'b1111111001100110000100110;
    rom[41219] = 25'b1111111001100100011001011;
    rom[41220] = 25'b1111111001100010101110000;
    rom[41221] = 25'b1111111001100001000010111;
    rom[41222] = 25'b1111111001011111010111101;
    rom[41223] = 25'b1111111001011101101100101;
    rom[41224] = 25'b1111111001011100000001101;
    rom[41225] = 25'b1111111001011010010110110;
    rom[41226] = 25'b1111111001011000101011111;
    rom[41227] = 25'b1111111001010111000001001;
    rom[41228] = 25'b1111111001010101010110100;
    rom[41229] = 25'b1111111001010011101100000;
    rom[41230] = 25'b1111111001010010000001100;
    rom[41231] = 25'b1111111001010000010111001;
    rom[41232] = 25'b1111111001001110101100111;
    rom[41233] = 25'b1111111001001101000010101;
    rom[41234] = 25'b1111111001001011011000100;
    rom[41235] = 25'b1111111001001001101110100;
    rom[41236] = 25'b1111111001001000000100100;
    rom[41237] = 25'b1111111001000110011010101;
    rom[41238] = 25'b1111111001000100110000111;
    rom[41239] = 25'b1111111001000011000111001;
    rom[41240] = 25'b1111111001000001011101100;
    rom[41241] = 25'b1111111000111111110100000;
    rom[41242] = 25'b1111111000111110001010101;
    rom[41243] = 25'b1111111000111100100001010;
    rom[41244] = 25'b1111111000111010111000000;
    rom[41245] = 25'b1111111000111001001110111;
    rom[41246] = 25'b1111111000110111100101110;
    rom[41247] = 25'b1111111000110101111100110;
    rom[41248] = 25'b1111111000110100010011111;
    rom[41249] = 25'b1111111000110010101011001;
    rom[41250] = 25'b1111111000110001000010010;
    rom[41251] = 25'b1111111000101111011001110;
    rom[41252] = 25'b1111111000101101110001001;
    rom[41253] = 25'b1111111000101100001000101;
    rom[41254] = 25'b1111111000101010100000010;
    rom[41255] = 25'b1111111000101000111000000;
    rom[41256] = 25'b1111111000100111001111110;
    rom[41257] = 25'b1111111000100101100111101;
    rom[41258] = 25'b1111111000100011111111101;
    rom[41259] = 25'b1111111000100010010111101;
    rom[41260] = 25'b1111111000100000101111110;
    rom[41261] = 25'b1111111000011111001000000;
    rom[41262] = 25'b1111111000011101100000011;
    rom[41263] = 25'b1111111000011011111000111;
    rom[41264] = 25'b1111111000011010010001011;
    rom[41265] = 25'b1111111000011000101001111;
    rom[41266] = 25'b1111111000010111000010101;
    rom[41267] = 25'b1111111000010101011011011;
    rom[41268] = 25'b1111111000010011110100010;
    rom[41269] = 25'b1111111000010010001101010;
    rom[41270] = 25'b1111111000010000100110010;
    rom[41271] = 25'b1111111000001110111111011;
    rom[41272] = 25'b1111111000001101011000101;
    rom[41273] = 25'b1111111000001011110001111;
    rom[41274] = 25'b1111111000001010001011010;
    rom[41275] = 25'b1111111000001000100100111;
    rom[41276] = 25'b1111111000000110111110011;
    rom[41277] = 25'b1111111000000101011000000;
    rom[41278] = 25'b1111111000000011110001111;
    rom[41279] = 25'b1111111000000010001011110;
    rom[41280] = 25'b1111111000000000100101101;
    rom[41281] = 25'b1111110111111110111111101;
    rom[41282] = 25'b1111110111111101011001110;
    rom[41283] = 25'b1111110111111011110100001;
    rom[41284] = 25'b1111110111111010001110011;
    rom[41285] = 25'b1111110111111000101000110;
    rom[41286] = 25'b1111110111110111000011010;
    rom[41287] = 25'b1111110111110101011101111;
    rom[41288] = 25'b1111110111110011111000100;
    rom[41289] = 25'b1111110111110010010011010;
    rom[41290] = 25'b1111110111110000101110001;
    rom[41291] = 25'b1111110111101111001001001;
    rom[41292] = 25'b1111110111101101100100001;
    rom[41293] = 25'b1111110111101011111111010;
    rom[41294] = 25'b1111110111101010011010100;
    rom[41295] = 25'b1111110111101000110101111;
    rom[41296] = 25'b1111110111100111010001010;
    rom[41297] = 25'b1111110111100101101100110;
    rom[41298] = 25'b1111110111100100001000011;
    rom[41299] = 25'b1111110111100010100100000;
    rom[41300] = 25'b1111110111100000111111111;
    rom[41301] = 25'b1111110111011111011011110;
    rom[41302] = 25'b1111110111011101110111110;
    rom[41303] = 25'b1111110111011100010011110;
    rom[41304] = 25'b1111110111011010101111111;
    rom[41305] = 25'b1111110111011001001100001;
    rom[41306] = 25'b1111110111010111101000100;
    rom[41307] = 25'b1111110111010110000100111;
    rom[41308] = 25'b1111110111010100100001100;
    rom[41309] = 25'b1111110111010010111110001;
    rom[41310] = 25'b1111110111010001011010111;
    rom[41311] = 25'b1111110111001111110111100;
    rom[41312] = 25'b1111110111001110010100100;
    rom[41313] = 25'b1111110111001100110001100;
    rom[41314] = 25'b1111110111001011001110101;
    rom[41315] = 25'b1111110111001001101011110;
    rom[41316] = 25'b1111110111001000001001001;
    rom[41317] = 25'b1111110111000110100110100;
    rom[41318] = 25'b1111110111000101000011111;
    rom[41319] = 25'b1111110111000011100001100;
    rom[41320] = 25'b1111110111000001111111001;
    rom[41321] = 25'b1111110111000000011100111;
    rom[41322] = 25'b1111110110111110111010101;
    rom[41323] = 25'b1111110110111101011000101;
    rom[41324] = 25'b1111110110111011110110101;
    rom[41325] = 25'b1111110110111010010100110;
    rom[41326] = 25'b1111110110111000110011000;
    rom[41327] = 25'b1111110110110111010001011;
    rom[41328] = 25'b1111110110110101101111110;
    rom[41329] = 25'b1111110110110100001110011;
    rom[41330] = 25'b1111110110110010101100111;
    rom[41331] = 25'b1111110110110001001011101;
    rom[41332] = 25'b1111110110101111101010011;
    rom[41333] = 25'b1111110110101110001001010;
    rom[41334] = 25'b1111110110101100101000010;
    rom[41335] = 25'b1111110110101011000111011;
    rom[41336] = 25'b1111110110101001100110101;
    rom[41337] = 25'b1111110110101000000101111;
    rom[41338] = 25'b1111110110100110100101010;
    rom[41339] = 25'b1111110110100101000100110;
    rom[41340] = 25'b1111110110100011100100010;
    rom[41341] = 25'b1111110110100010000100000;
    rom[41342] = 25'b1111110110100000100011101;
    rom[41343] = 25'b1111110110011111000011101;
    rom[41344] = 25'b1111110110011101100011100;
    rom[41345] = 25'b1111110110011100000011101;
    rom[41346] = 25'b1111110110011010100011101;
    rom[41347] = 25'b1111110110011001000100000;
    rom[41348] = 25'b1111110110010111100100010;
    rom[41349] = 25'b1111110110010110000100101;
    rom[41350] = 25'b1111110110010100100101010;
    rom[41351] = 25'b1111110110010011000101111;
    rom[41352] = 25'b1111110110010001100110101;
    rom[41353] = 25'b1111110110010000000111100;
    rom[41354] = 25'b1111110110001110101000011;
    rom[41355] = 25'b1111110110001101001001011;
    rom[41356] = 25'b1111110110001011101010100;
    rom[41357] = 25'b1111110110001010001011110;
    rom[41358] = 25'b1111110110001000101101001;
    rom[41359] = 25'b1111110110000111001110100;
    rom[41360] = 25'b1111110110000101110000000;
    rom[41361] = 25'b1111110110000100010001100;
    rom[41362] = 25'b1111110110000010110011011;
    rom[41363] = 25'b1111110110000001010101001;
    rom[41364] = 25'b1111110101111111110111000;
    rom[41365] = 25'b1111110101111110011001000;
    rom[41366] = 25'b1111110101111100111011001;
    rom[41367] = 25'b1111110101111011011101010;
    rom[41368] = 25'b1111110101111001111111101;
    rom[41369] = 25'b1111110101111000100010000;
    rom[41370] = 25'b1111110101110111000100100;
    rom[41371] = 25'b1111110101110101100111001;
    rom[41372] = 25'b1111110101110100001001110;
    rom[41373] = 25'b1111110101110010101100101;
    rom[41374] = 25'b1111110101110001001111100;
    rom[41375] = 25'b1111110101101111110010100;
    rom[41376] = 25'b1111110101101110010101101;
    rom[41377] = 25'b1111110101101100111000110;
    rom[41378] = 25'b1111110101101011011100001;
    rom[41379] = 25'b1111110101101001111111100;
    rom[41380] = 25'b1111110101101000100010111;
    rom[41381] = 25'b1111110101100111000110100;
    rom[41382] = 25'b1111110101100101101010010;
    rom[41383] = 25'b1111110101100100001110000;
    rom[41384] = 25'b1111110101100010110010000;
    rom[41385] = 25'b1111110101100001010101111;
    rom[41386] = 25'b1111110101011111111010000;
    rom[41387] = 25'b1111110101011110011110001;
    rom[41388] = 25'b1111110101011101000010100;
    rom[41389] = 25'b1111110101011011100110111;
    rom[41390] = 25'b1111110101011010001011011;
    rom[41391] = 25'b1111110101011000110000000;
    rom[41392] = 25'b1111110101010111010100101;
    rom[41393] = 25'b1111110101010101111001011;
    rom[41394] = 25'b1111110101010100011110011;
    rom[41395] = 25'b1111110101010011000011011;
    rom[41396] = 25'b1111110101010001101000100;
    rom[41397] = 25'b1111110101010000001101101;
    rom[41398] = 25'b1111110101001110110010111;
    rom[41399] = 25'b1111110101001101011000011;
    rom[41400] = 25'b1111110101001011111101111;
    rom[41401] = 25'b1111110101001010100011100;
    rom[41402] = 25'b1111110101001001001001001;
    rom[41403] = 25'b1111110101000111101110111;
    rom[41404] = 25'b1111110101000110010100111;
    rom[41405] = 25'b1111110101000100111010111;
    rom[41406] = 25'b1111110101000011100001000;
    rom[41407] = 25'b1111110101000010000111010;
    rom[41408] = 25'b1111110101000000101101100;
    rom[41409] = 25'b1111110100111111010100000;
    rom[41410] = 25'b1111110100111101111010011;
    rom[41411] = 25'b1111110100111100100001000;
    rom[41412] = 25'b1111110100111011000111110;
    rom[41413] = 25'b1111110100111001101110101;
    rom[41414] = 25'b1111110100111000010101101;
    rom[41415] = 25'b1111110100110110111100101;
    rom[41416] = 25'b1111110100110101100011110;
    rom[41417] = 25'b1111110100110100001011000;
    rom[41418] = 25'b1111110100110010110010011;
    rom[41419] = 25'b1111110100110001011001110;
    rom[41420] = 25'b1111110100110000000001010;
    rom[41421] = 25'b1111110100101110101001000;
    rom[41422] = 25'b1111110100101101010000110;
    rom[41423] = 25'b1111110100101011111000100;
    rom[41424] = 25'b1111110100101010100000100;
    rom[41425] = 25'b1111110100101001001000101;
    rom[41426] = 25'b1111110100100111110000110;
    rom[41427] = 25'b1111110100100110011001000;
    rom[41428] = 25'b1111110100100101000001011;
    rom[41429] = 25'b1111110100100011101001111;
    rom[41430] = 25'b1111110100100010010010011;
    rom[41431] = 25'b1111110100100000111011001;
    rom[41432] = 25'b1111110100011111100011111;
    rom[41433] = 25'b1111110100011110001100110;
    rom[41434] = 25'b1111110100011100110101110;
    rom[41435] = 25'b1111110100011011011110111;
    rom[41436] = 25'b1111110100011010001000001;
    rom[41437] = 25'b1111110100011000110001011;
    rom[41438] = 25'b1111110100010111011010110;
    rom[41439] = 25'b1111110100010110000100010;
    rom[41440] = 25'b1111110100010100101101111;
    rom[41441] = 25'b1111110100010011010111101;
    rom[41442] = 25'b1111110100010010000001100;
    rom[41443] = 25'b1111110100010000101011011;
    rom[41444] = 25'b1111110100001111010101011;
    rom[41445] = 25'b1111110100001101111111101;
    rom[41446] = 25'b1111110100001100101001110;
    rom[41447] = 25'b1111110100001011010100001;
    rom[41448] = 25'b1111110100001001111110101;
    rom[41449] = 25'b1111110100001000101001001;
    rom[41450] = 25'b1111110100000111010011111;
    rom[41451] = 25'b1111110100000101111110101;
    rom[41452] = 25'b1111110100000100101001100;
    rom[41453] = 25'b1111110100000011010100100;
    rom[41454] = 25'b1111110100000001111111101;
    rom[41455] = 25'b1111110100000000101010110;
    rom[41456] = 25'b1111110011111111010110000;
    rom[41457] = 25'b1111110011111110000001100;
    rom[41458] = 25'b1111110011111100101101000;
    rom[41459] = 25'b1111110011111011011000100;
    rom[41460] = 25'b1111110011111010000100010;
    rom[41461] = 25'b1111110011111000110000001;
    rom[41462] = 25'b1111110011110111011100000;
    rom[41463] = 25'b1111110011110110001000001;
    rom[41464] = 25'b1111110011110100110100010;
    rom[41465] = 25'b1111110011110011100000011;
    rom[41466] = 25'b1111110011110010001100110;
    rom[41467] = 25'b1111110011110000111001010;
    rom[41468] = 25'b1111110011101111100101110;
    rom[41469] = 25'b1111110011101110010010100;
    rom[41470] = 25'b1111110011101100111111010;
    rom[41471] = 25'b1111110011101011101100001;
    rom[41472] = 25'b1111110011101010011001001;
    rom[41473] = 25'b1111110011101001000110010;
    rom[41474] = 25'b1111110011100111110011100;
    rom[41475] = 25'b1111110011100110100000110;
    rom[41476] = 25'b1111110011100101001110001;
    rom[41477] = 25'b1111110011100011111011110;
    rom[41478] = 25'b1111110011100010101001011;
    rom[41479] = 25'b1111110011100001010111001;
    rom[41480] = 25'b1111110011100000000100111;
    rom[41481] = 25'b1111110011011110110010111;
    rom[41482] = 25'b1111110011011101100000111;
    rom[41483] = 25'b1111110011011100001111001;
    rom[41484] = 25'b1111110011011010111101011;
    rom[41485] = 25'b1111110011011001101011110;
    rom[41486] = 25'b1111110011011000011010010;
    rom[41487] = 25'b1111110011010111001000110;
    rom[41488] = 25'b1111110011010101110111100;
    rom[41489] = 25'b1111110011010100100110010;
    rom[41490] = 25'b1111110011010011010101010;
    rom[41491] = 25'b1111110011010010000100010;
    rom[41492] = 25'b1111110011010000110011011;
    rom[41493] = 25'b1111110011001111100010101;
    rom[41494] = 25'b1111110011001110010010000;
    rom[41495] = 25'b1111110011001101000001100;
    rom[41496] = 25'b1111110011001011110001000;
    rom[41497] = 25'b1111110011001010100000110;
    rom[41498] = 25'b1111110011001001010000100;
    rom[41499] = 25'b1111110011001000000000011;
    rom[41500] = 25'b1111110011000110110000011;
    rom[41501] = 25'b1111110011000101100000100;
    rom[41502] = 25'b1111110011000100010000101;
    rom[41503] = 25'b1111110011000011000001000;
    rom[41504] = 25'b1111110011000001110001011;
    rom[41505] = 25'b1111110011000000100010000;
    rom[41506] = 25'b1111110010111111010010101;
    rom[41507] = 25'b1111110010111110000011011;
    rom[41508] = 25'b1111110010111100110100010;
    rom[41509] = 25'b1111110010111011100101010;
    rom[41510] = 25'b1111110010111010010110010;
    rom[41511] = 25'b1111110010111001000111100;
    rom[41512] = 25'b1111110010110111111000111;
    rom[41513] = 25'b1111110010110110101010010;
    rom[41514] = 25'b1111110010110101011011110;
    rom[41515] = 25'b1111110010110100001101011;
    rom[41516] = 25'b1111110010110010111111001;
    rom[41517] = 25'b1111110010110001110001000;
    rom[41518] = 25'b1111110010110000100010111;
    rom[41519] = 25'b1111110010101111010100111;
    rom[41520] = 25'b1111110010101110000111001;
    rom[41521] = 25'b1111110010101100111001011;
    rom[41522] = 25'b1111110010101011101011111;
    rom[41523] = 25'b1111110010101010011110011;
    rom[41524] = 25'b1111110010101001010000111;
    rom[41525] = 25'b1111110010101000000011101;
    rom[41526] = 25'b1111110010100110110110100;
    rom[41527] = 25'b1111110010100101101001011;
    rom[41528] = 25'b1111110010100100011100100;
    rom[41529] = 25'b1111110010100011001111101;
    rom[41530] = 25'b1111110010100010000010111;
    rom[41531] = 25'b1111110010100000110110010;
    rom[41532] = 25'b1111110010011111101001110;
    rom[41533] = 25'b1111110010011110011101011;
    rom[41534] = 25'b1111110010011101010001001;
    rom[41535] = 25'b1111110010011100000100111;
    rom[41536] = 25'b1111110010011010111000111;
    rom[41537] = 25'b1111110010011001101100111;
    rom[41538] = 25'b1111110010011000100001000;
    rom[41539] = 25'b1111110010010111010101010;
    rom[41540] = 25'b1111110010010110001001110;
    rom[41541] = 25'b1111110010010100111110001;
    rom[41542] = 25'b1111110010010011110010110;
    rom[41543] = 25'b1111110010010010100111100;
    rom[41544] = 25'b1111110010010001011100010;
    rom[41545] = 25'b1111110010010000010001001;
    rom[41546] = 25'b1111110010001111000110010;
    rom[41547] = 25'b1111110010001101111011011;
    rom[41548] = 25'b1111110010001100110000101;
    rom[41549] = 25'b1111110010001011100110001;
    rom[41550] = 25'b1111110010001010011011100;
    rom[41551] = 25'b1111110010001001010001001;
    rom[41552] = 25'b1111110010001000000110110;
    rom[41553] = 25'b1111110010000110111100101;
    rom[41554] = 25'b1111110010000101110010101;
    rom[41555] = 25'b1111110010000100101000101;
    rom[41556] = 25'b1111110010000011011110110;
    rom[41557] = 25'b1111110010000010010101000;
    rom[41558] = 25'b1111110010000001001011011;
    rom[41559] = 25'b1111110010000000000001111;
    rom[41560] = 25'b1111110001111110111000100;
    rom[41561] = 25'b1111110001111101101111001;
    rom[41562] = 25'b1111110001111100100110000;
    rom[41563] = 25'b1111110001111011011100111;
    rom[41564] = 25'b1111110001111010010011111;
    rom[41565] = 25'b1111110001111001001011000;
    rom[41566] = 25'b1111110001111000000010010;
    rom[41567] = 25'b1111110001110110111001110;
    rom[41568] = 25'b1111110001110101110001001;
    rom[41569] = 25'b1111110001110100101000110;
    rom[41570] = 25'b1111110001110011100000100;
    rom[41571] = 25'b1111110001110010011000011;
    rom[41572] = 25'b1111110001110001010000010;
    rom[41573] = 25'b1111110001110000001000011;
    rom[41574] = 25'b1111110001101111000000100;
    rom[41575] = 25'b1111110001101101111000110;
    rom[41576] = 25'b1111110001101100110001001;
    rom[41577] = 25'b1111110001101011101001101;
    rom[41578] = 25'b1111110001101010100010010;
    rom[41579] = 25'b1111110001101001011011000;
    rom[41580] = 25'b1111110001101000010011110;
    rom[41581] = 25'b1111110001100111001100110;
    rom[41582] = 25'b1111110001100110000101111;
    rom[41583] = 25'b1111110001100100111111000;
    rom[41584] = 25'b1111110001100011111000010;
    rom[41585] = 25'b1111110001100010110001101;
    rom[41586] = 25'b1111110001100001101011001;
    rom[41587] = 25'b1111110001100000100100111;
    rom[41588] = 25'b1111110001011111011110100;
    rom[41589] = 25'b1111110001011110011000011;
    rom[41590] = 25'b1111110001011101010010011;
    rom[41591] = 25'b1111110001011100001100011;
    rom[41592] = 25'b1111110001011011000110101;
    rom[41593] = 25'b1111110001011010000001000;
    rom[41594] = 25'b1111110001011000111011010;
    rom[41595] = 25'b1111110001010111110101111;
    rom[41596] = 25'b1111110001010110110000100;
    rom[41597] = 25'b1111110001010101101011010;
    rom[41598] = 25'b1111110001010100100110001;
    rom[41599] = 25'b1111110001010011100001001;
    rom[41600] = 25'b1111110001010010011100010;
    rom[41601] = 25'b1111110001010001010111100;
    rom[41602] = 25'b1111110001010000010010110;
    rom[41603] = 25'b1111110001001111001110001;
    rom[41604] = 25'b1111110001001110001001110;
    rom[41605] = 25'b1111110001001101000101011;
    rom[41606] = 25'b1111110001001100000001010;
    rom[41607] = 25'b1111110001001010111101000;
    rom[41608] = 25'b1111110001001001111001000;
    rom[41609] = 25'b1111110001001000110101001;
    rom[41610] = 25'b1111110001000111110001011;
    rom[41611] = 25'b1111110001000110101101110;
    rom[41612] = 25'b1111110001000101101010010;
    rom[41613] = 25'b1111110001000100100110110;
    rom[41614] = 25'b1111110001000011100011100;
    rom[41615] = 25'b1111110001000010100000010;
    rom[41616] = 25'b1111110001000001011101001;
    rom[41617] = 25'b1111110001000000011010010;
    rom[41618] = 25'b1111110000111111010111011;
    rom[41619] = 25'b1111110000111110010100101;
    rom[41620] = 25'b1111110000111101010010000;
    rom[41621] = 25'b1111110000111100001111011;
    rom[41622] = 25'b1111110000111011001101000;
    rom[41623] = 25'b1111110000111010001010110;
    rom[41624] = 25'b1111110000111001001000101;
    rom[41625] = 25'b1111110000111000000110100;
    rom[41626] = 25'b1111110000110111000100101;
    rom[41627] = 25'b1111110000110110000010110;
    rom[41628] = 25'b1111110000110101000001000;
    rom[41629] = 25'b1111110000110011111111100;
    rom[41630] = 25'b1111110000110010111101111;
    rom[41631] = 25'b1111110000110001111100100;
    rom[41632] = 25'b1111110000110000111011011;
    rom[41633] = 25'b1111110000101111111010001;
    rom[41634] = 25'b1111110000101110111001010;
    rom[41635] = 25'b1111110000101101111000010;
    rom[41636] = 25'b1111110000101100110111100;
    rom[41637] = 25'b1111110000101011110110110;
    rom[41638] = 25'b1111110000101010110110010;
    rom[41639] = 25'b1111110000101001110101110;
    rom[41640] = 25'b1111110000101000110101100;
    rom[41641] = 25'b1111110000100111110101010;
    rom[41642] = 25'b1111110000100110110101000;
    rom[41643] = 25'b1111110000100101110101001;
    rom[41644] = 25'b1111110000100100110101010;
    rom[41645] = 25'b1111110000100011110101011;
    rom[41646] = 25'b1111110000100010110101110;
    rom[41647] = 25'b1111110000100001110110010;
    rom[41648] = 25'b1111110000100000110110111;
    rom[41649] = 25'b1111110000011111110111101;
    rom[41650] = 25'b1111110000011110111000011;
    rom[41651] = 25'b1111110000011101111001011;
    rom[41652] = 25'b1111110000011100111010011;
    rom[41653] = 25'b1111110000011011111011100;
    rom[41654] = 25'b1111110000011010111100110;
    rom[41655] = 25'b1111110000011001111110010;
    rom[41656] = 25'b1111110000011000111111101;
    rom[41657] = 25'b1111110000011000000001010;
    rom[41658] = 25'b1111110000010111000011000;
    rom[41659] = 25'b1111110000010110000100111;
    rom[41660] = 25'b1111110000010101000110111;
    rom[41661] = 25'b1111110000010100001000111;
    rom[41662] = 25'b1111110000010011001011001;
    rom[41663] = 25'b1111110000010010001101100;
    rom[41664] = 25'b1111110000010001001111111;
    rom[41665] = 25'b1111110000010000010010011;
    rom[41666] = 25'b1111110000001111010101001;
    rom[41667] = 25'b1111110000001110010111111;
    rom[41668] = 25'b1111110000001101011010110;
    rom[41669] = 25'b1111110000001100011101111;
    rom[41670] = 25'b1111110000001011100000111;
    rom[41671] = 25'b1111110000001010100100001;
    rom[41672] = 25'b1111110000001001100111100;
    rom[41673] = 25'b1111110000001000101011000;
    rom[41674] = 25'b1111110000000111101110101;
    rom[41675] = 25'b1111110000000110110010010;
    rom[41676] = 25'b1111110000000101110110001;
    rom[41677] = 25'b1111110000000100111010001;
    rom[41678] = 25'b1111110000000011111110001;
    rom[41679] = 25'b1111110000000011000010010;
    rom[41680] = 25'b1111110000000010000110101;
    rom[41681] = 25'b1111110000000001001011000;
    rom[41682] = 25'b1111110000000000001111100;
    rom[41683] = 25'b1111101111111111010100001;
    rom[41684] = 25'b1111101111111110011000111;
    rom[41685] = 25'b1111101111111101011101110;
    rom[41686] = 25'b1111101111111100100010110;
    rom[41687] = 25'b1111101111111011100111111;
    rom[41688] = 25'b1111101111111010101101001;
    rom[41689] = 25'b1111101111111001110010011;
    rom[41690] = 25'b1111101111111000110111111;
    rom[41691] = 25'b1111101111110111111101100;
    rom[41692] = 25'b1111101111110111000011001;
    rom[41693] = 25'b1111101111110110001000111;
    rom[41694] = 25'b1111101111110101001110111;
    rom[41695] = 25'b1111101111110100010100111;
    rom[41696] = 25'b1111101111110011011011000;
    rom[41697] = 25'b1111101111110010100001010;
    rom[41698] = 25'b1111101111110001100111101;
    rom[41699] = 25'b1111101111110000101110001;
    rom[41700] = 25'b1111101111101111110100111;
    rom[41701] = 25'b1111101111101110111011101;
    rom[41702] = 25'b1111101111101110000010011;
    rom[41703] = 25'b1111101111101101001001011;
    rom[41704] = 25'b1111101111101100010000100;
    rom[41705] = 25'b1111101111101011010111101;
    rom[41706] = 25'b1111101111101010011110111;
    rom[41707] = 25'b1111101111101001100110011;
    rom[41708] = 25'b1111101111101000101101111;
    rom[41709] = 25'b1111101111100111110101101;
    rom[41710] = 25'b1111101111100110111101011;
    rom[41711] = 25'b1111101111100110000101011;
    rom[41712] = 25'b1111101111100101001101011;
    rom[41713] = 25'b1111101111100100010101100;
    rom[41714] = 25'b1111101111100011011101110;
    rom[41715] = 25'b1111101111100010100110001;
    rom[41716] = 25'b1111101111100001101110101;
    rom[41717] = 25'b1111101111100000110111010;
    rom[41718] = 25'b1111101111100000000000000;
    rom[41719] = 25'b1111101111011111001000110;
    rom[41720] = 25'b1111101111011110010001110;
    rom[41721] = 25'b1111101111011101011010111;
    rom[41722] = 25'b1111101111011100100100000;
    rom[41723] = 25'b1111101111011011101101010;
    rom[41724] = 25'b1111101111011010110110110;
    rom[41725] = 25'b1111101111011010000000010;
    rom[41726] = 25'b1111101111011001001010000;
    rom[41727] = 25'b1111101111011000010011110;
    rom[41728] = 25'b1111101111010111011101101;
    rom[41729] = 25'b1111101111010110100111101;
    rom[41730] = 25'b1111101111010101110001111;
    rom[41731] = 25'b1111101111010100111100001;
    rom[41732] = 25'b1111101111010100000110100;
    rom[41733] = 25'b1111101111010011010001000;
    rom[41734] = 25'b1111101111010010011011100;
    rom[41735] = 25'b1111101111010001100110010;
    rom[41736] = 25'b1111101111010000110001001;
    rom[41737] = 25'b1111101111001111111100000;
    rom[41738] = 25'b1111101111001111000111001;
    rom[41739] = 25'b1111101111001110010010011;
    rom[41740] = 25'b1111101111001101011101101;
    rom[41741] = 25'b1111101111001100101001001;
    rom[41742] = 25'b1111101111001011110100101;
    rom[41743] = 25'b1111101111001011000000010;
    rom[41744] = 25'b1111101111001010001100001;
    rom[41745] = 25'b1111101111001001011000000;
    rom[41746] = 25'b1111101111001000100100000;
    rom[41747] = 25'b1111101111000111110000001;
    rom[41748] = 25'b1111101111000110111100011;
    rom[41749] = 25'b1111101111000110001000110;
    rom[41750] = 25'b1111101111000101010101010;
    rom[41751] = 25'b1111101111000100100001111;
    rom[41752] = 25'b1111101111000011101110101;
    rom[41753] = 25'b1111101111000010111011011;
    rom[41754] = 25'b1111101111000010001000010;
    rom[41755] = 25'b1111101111000001010101011;
    rom[41756] = 25'b1111101111000000100010101;
    rom[41757] = 25'b1111101110111111101111111;
    rom[41758] = 25'b1111101110111110111101011;
    rom[41759] = 25'b1111101110111110001011000;
    rom[41760] = 25'b1111101110111101011000101;
    rom[41761] = 25'b1111101110111100100110011;
    rom[41762] = 25'b1111101110111011110100011;
    rom[41763] = 25'b1111101110111011000010010;
    rom[41764] = 25'b1111101110111010010000100;
    rom[41765] = 25'b1111101110111001011110110;
    rom[41766] = 25'b1111101110111000101101001;
    rom[41767] = 25'b1111101110110111111011100;
    rom[41768] = 25'b1111101110110111001010010;
    rom[41769] = 25'b1111101110110110011000111;
    rom[41770] = 25'b1111101110110101100111110;
    rom[41771] = 25'b1111101110110100110110110;
    rom[41772] = 25'b1111101110110100000101111;
    rom[41773] = 25'b1111101110110011010101000;
    rom[41774] = 25'b1111101110110010100100011;
    rom[41775] = 25'b1111101110110001110011110;
    rom[41776] = 25'b1111101110110001000011011;
    rom[41777] = 25'b1111101110110000010011000;
    rom[41778] = 25'b1111101110101111100010111;
    rom[41779] = 25'b1111101110101110110010110;
    rom[41780] = 25'b1111101110101110000010110;
    rom[41781] = 25'b1111101110101101010010111;
    rom[41782] = 25'b1111101110101100100011010;
    rom[41783] = 25'b1111101110101011110011101;
    rom[41784] = 25'b1111101110101011000100000;
    rom[41785] = 25'b1111101110101010010100110;
    rom[41786] = 25'b1111101110101001100101100;
    rom[41787] = 25'b1111101110101000110110010;
    rom[41788] = 25'b1111101110101000000111010;
    rom[41789] = 25'b1111101110100111011000011;
    rom[41790] = 25'b1111101110100110101001101;
    rom[41791] = 25'b1111101110100101111011000;
    rom[41792] = 25'b1111101110100101001100100;
    rom[41793] = 25'b1111101110100100011101111;
    rom[41794] = 25'b1111101110100011101111101;
    rom[41795] = 25'b1111101110100011000001100;
    rom[41796] = 25'b1111101110100010010011011;
    rom[41797] = 25'b1111101110100001100101011;
    rom[41798] = 25'b1111101110100000110111101;
    rom[41799] = 25'b1111101110100000001001111;
    rom[41800] = 25'b1111101110011111011100010;
    rom[41801] = 25'b1111101110011110101110111;
    rom[41802] = 25'b1111101110011110000001100;
    rom[41803] = 25'b1111101110011101010100010;
    rom[41804] = 25'b1111101110011100100111000;
    rom[41805] = 25'b1111101110011011111010000;
    rom[41806] = 25'b1111101110011011001101010;
    rom[41807] = 25'b1111101110011010100000011;
    rom[41808] = 25'b1111101110011001110011110;
    rom[41809] = 25'b1111101110011001000111010;
    rom[41810] = 25'b1111101110011000011010111;
    rom[41811] = 25'b1111101110010111101110101;
    rom[41812] = 25'b1111101110010111000010011;
    rom[41813] = 25'b1111101110010110010110011;
    rom[41814] = 25'b1111101110010101101010011;
    rom[41815] = 25'b1111101110010100111110100;
    rom[41816] = 25'b1111101110010100010010111;
    rom[41817] = 25'b1111101110010011100111010;
    rom[41818] = 25'b1111101110010010111011110;
    rom[41819] = 25'b1111101110010010010000100;
    rom[41820] = 25'b1111101110010001100101010;
    rom[41821] = 25'b1111101110010000111010001;
    rom[41822] = 25'b1111101110010000001111001;
    rom[41823] = 25'b1111101110001111100100010;
    rom[41824] = 25'b1111101110001110111001100;
    rom[41825] = 25'b1111101110001110001110111;
    rom[41826] = 25'b1111101110001101100100011;
    rom[41827] = 25'b1111101110001100111001111;
    rom[41828] = 25'b1111101110001100001111110;
    rom[41829] = 25'b1111101110001011100101100;
    rom[41830] = 25'b1111101110001010111011100;
    rom[41831] = 25'b1111101110001010010001100;
    rom[41832] = 25'b1111101110001001100111110;
    rom[41833] = 25'b1111101110001000111110000;
    rom[41834] = 25'b1111101110001000010100100;
    rom[41835] = 25'b1111101110000111101011000;
    rom[41836] = 25'b1111101110000111000001110;
    rom[41837] = 25'b1111101110000110011000101;
    rom[41838] = 25'b1111101110000101101111100;
    rom[41839] = 25'b1111101110000101000110100;
    rom[41840] = 25'b1111101110000100011101101;
    rom[41841] = 25'b1111101110000011110100111;
    rom[41842] = 25'b1111101110000011001100010;
    rom[41843] = 25'b1111101110000010100011110;
    rom[41844] = 25'b1111101110000001111011011;
    rom[41845] = 25'b1111101110000001010011001;
    rom[41846] = 25'b1111101110000000101011000;
    rom[41847] = 25'b1111101110000000000011000;
    rom[41848] = 25'b1111101101111111011011001;
    rom[41849] = 25'b1111101101111110110011011;
    rom[41850] = 25'b1111101101111110001011101;
    rom[41851] = 25'b1111101101111101100100000;
    rom[41852] = 25'b1111101101111100111100101;
    rom[41853] = 25'b1111101101111100010101011;
    rom[41854] = 25'b1111101101111011101110010;
    rom[41855] = 25'b1111101101111011000111001;
    rom[41856] = 25'b1111101101111010100000001;
    rom[41857] = 25'b1111101101111001111001010;
    rom[41858] = 25'b1111101101111001010010101;
    rom[41859] = 25'b1111101101111000101100000;
    rom[41860] = 25'b1111101101111000000101101;
    rom[41861] = 25'b1111101101110111011111001;
    rom[41862] = 25'b1111101101110110111000111;
    rom[41863] = 25'b1111101101110110010010110;
    rom[41864] = 25'b1111101101110101101100110;
    rom[41865] = 25'b1111101101110101000111000;
    rom[41866] = 25'b1111101101110100100001001;
    rom[41867] = 25'b1111101101110011111011100;
    rom[41868] = 25'b1111101101110011010110000;
    rom[41869] = 25'b1111101101110010110000101;
    rom[41870] = 25'b1111101101110010001011010;
    rom[41871] = 25'b1111101101110001100110001;
    rom[41872] = 25'b1111101101110001000001001;
    rom[41873] = 25'b1111101101110000011100001;
    rom[41874] = 25'b1111101101101111110111011;
    rom[41875] = 25'b1111101101101111010010101;
    rom[41876] = 25'b1111101101101110101110000;
    rom[41877] = 25'b1111101101101110001001101;
    rom[41878] = 25'b1111101101101101100101010;
    rom[41879] = 25'b1111101101101101000001000;
    rom[41880] = 25'b1111101101101100011100111;
    rom[41881] = 25'b1111101101101011111001000;
    rom[41882] = 25'b1111101101101011010101001;
    rom[41883] = 25'b1111101101101010110001011;
    rom[41884] = 25'b1111101101101010001101110;
    rom[41885] = 25'b1111101101101001101010010;
    rom[41886] = 25'b1111101101101001000110111;
    rom[41887] = 25'b1111101101101000100011100;
    rom[41888] = 25'b1111101101101000000000100;
    rom[41889] = 25'b1111101101100111011101011;
    rom[41890] = 25'b1111101101100110111010100;
    rom[41891] = 25'b1111101101100110010111101;
    rom[41892] = 25'b1111101101100101110101000;
    rom[41893] = 25'b1111101101100101010010100;
    rom[41894] = 25'b1111101101100100110000000;
    rom[41895] = 25'b1111101101100100001101101;
    rom[41896] = 25'b1111101101100011101011100;
    rom[41897] = 25'b1111101101100011001001011;
    rom[41898] = 25'b1111101101100010100111011;
    rom[41899] = 25'b1111101101100010000101101;
    rom[41900] = 25'b1111101101100001100011111;
    rom[41901] = 25'b1111101101100001000010010;
    rom[41902] = 25'b1111101101100000100000110;
    rom[41903] = 25'b1111101101011111111111011;
    rom[41904] = 25'b1111101101011111011110001;
    rom[41905] = 25'b1111101101011110111101000;
    rom[41906] = 25'b1111101101011110011011111;
    rom[41907] = 25'b1111101101011101111011000;
    rom[41908] = 25'b1111101101011101011010010;
    rom[41909] = 25'b1111101101011100111001101;
    rom[41910] = 25'b1111101101011100011001001;
    rom[41911] = 25'b1111101101011011111000101;
    rom[41912] = 25'b1111101101011011011000011;
    rom[41913] = 25'b1111101101011010111000001;
    rom[41914] = 25'b1111101101011010011000001;
    rom[41915] = 25'b1111101101011001111000001;
    rom[41916] = 25'b1111101101011001011000011;
    rom[41917] = 25'b1111101101011000111000101;
    rom[41918] = 25'b1111101101011000011001000;
    rom[41919] = 25'b1111101101010111111001100;
    rom[41920] = 25'b1111101101010111011010001;
    rom[41921] = 25'b1111101101010110111011000;
    rom[41922] = 25'b1111101101010110011011110;
    rom[41923] = 25'b1111101101010101111100110;
    rom[41924] = 25'b1111101101010101011110000;
    rom[41925] = 25'b1111101101010100111111001;
    rom[41926] = 25'b1111101101010100100000100;
    rom[41927] = 25'b1111101101010100000010000;
    rom[41928] = 25'b1111101101010011100011100;
    rom[41929] = 25'b1111101101010011000101010;
    rom[41930] = 25'b1111101101010010100111001;
    rom[41931] = 25'b1111101101010010001001000;
    rom[41932] = 25'b1111101101010001101011001;
    rom[41933] = 25'b1111101101010001001101010;
    rom[41934] = 25'b1111101101010000101111101;
    rom[41935] = 25'b1111101101010000010010000;
    rom[41936] = 25'b1111101101001111110100100;
    rom[41937] = 25'b1111101101001111010111010;
    rom[41938] = 25'b1111101101001110111010000;
    rom[41939] = 25'b1111101101001110011100111;
    rom[41940] = 25'b1111101101001101111111111;
    rom[41941] = 25'b1111101101001101100011000;
    rom[41942] = 25'b1111101101001101000110010;
    rom[41943] = 25'b1111101101001100101001101;
    rom[41944] = 25'b1111101101001100001101000;
    rom[41945] = 25'b1111101101001011110000101;
    rom[41946] = 25'b1111101101001011010100011;
    rom[41947] = 25'b1111101101001010111000010;
    rom[41948] = 25'b1111101101001010011100010;
    rom[41949] = 25'b1111101101001010000000010;
    rom[41950] = 25'b1111101101001001100100100;
    rom[41951] = 25'b1111101101001001001000110;
    rom[41952] = 25'b1111101101001000101101010;
    rom[41953] = 25'b1111101101001000010001110;
    rom[41954] = 25'b1111101101000111110110011;
    rom[41955] = 25'b1111101101000111011011010;
    rom[41956] = 25'b1111101101000111000000000;
    rom[41957] = 25'b1111101101000110100101000;
    rom[41958] = 25'b1111101101000110001010010;
    rom[41959] = 25'b1111101101000101101111011;
    rom[41960] = 25'b1111101101000101010100111;
    rom[41961] = 25'b1111101101000100111010010;
    rom[41962] = 25'b1111101101000100100000000;
    rom[41963] = 25'b1111101101000100000101101;
    rom[41964] = 25'b1111101101000011101011100;
    rom[41965] = 25'b1111101101000011010001011;
    rom[41966] = 25'b1111101101000010110111100;
    rom[41967] = 25'b1111101101000010011101110;
    rom[41968] = 25'b1111101101000010000100000;
    rom[41969] = 25'b1111101101000001101010011;
    rom[41970] = 25'b1111101101000001010001000;
    rom[41971] = 25'b1111101101000000110111110;
    rom[41972] = 25'b1111101101000000011110100;
    rom[41973] = 25'b1111101101000000000101011;
    rom[41974] = 25'b1111101100111111101100011;
    rom[41975] = 25'b1111101100111111010011100;
    rom[41976] = 25'b1111101100111110111010110;
    rom[41977] = 25'b1111101100111110100010001;
    rom[41978] = 25'b1111101100111110001001101;
    rom[41979] = 25'b1111101100111101110001010;
    rom[41980] = 25'b1111101100111101011001000;
    rom[41981] = 25'b1111101100111101000000110;
    rom[41982] = 25'b1111101100111100101000110;
    rom[41983] = 25'b1111101100111100010000110;
    rom[41984] = 25'b1111101100111011111001000;
    rom[41985] = 25'b1111101100111011100001011;
    rom[41986] = 25'b1111101100111011001001110;
    rom[41987] = 25'b1111101100111010110010010;
    rom[41988] = 25'b1111101100111010011011000;
    rom[41989] = 25'b1111101100111010000011110;
    rom[41990] = 25'b1111101100111001101100101;
    rom[41991] = 25'b1111101100111001010101101;
    rom[41992] = 25'b1111101100111000111110110;
    rom[41993] = 25'b1111101100111000101000001;
    rom[41994] = 25'b1111101100111000010001011;
    rom[41995] = 25'b1111101100110111111010111;
    rom[41996] = 25'b1111101100110111100100100;
    rom[41997] = 25'b1111101100110111001110010;
    rom[41998] = 25'b1111101100110110111000000;
    rom[41999] = 25'b1111101100110110100010000;
    rom[42000] = 25'b1111101100110110001100000;
    rom[42001] = 25'b1111101100110101110110010;
    rom[42002] = 25'b1111101100110101100000100;
    rom[42003] = 25'b1111101100110101001010111;
    rom[42004] = 25'b1111101100110100110101100;
    rom[42005] = 25'b1111101100110100100000001;
    rom[42006] = 25'b1111101100110100001011000;
    rom[42007] = 25'b1111101100110011110101111;
    rom[42008] = 25'b1111101100110011100000111;
    rom[42009] = 25'b1111101100110011001011111;
    rom[42010] = 25'b1111101100110010110111010;
    rom[42011] = 25'b1111101100110010100010100;
    rom[42012] = 25'b1111101100110010001110000;
    rom[42013] = 25'b1111101100110001111001100;
    rom[42014] = 25'b1111101100110001100101010;
    rom[42015] = 25'b1111101100110001010001001;
    rom[42016] = 25'b1111101100110000111101000;
    rom[42017] = 25'b1111101100110000101001001;
    rom[42018] = 25'b1111101100110000010101010;
    rom[42019] = 25'b1111101100110000000001100;
    rom[42020] = 25'b1111101100101111101110000;
    rom[42021] = 25'b1111101100101111011010100;
    rom[42022] = 25'b1111101100101111000111010;
    rom[42023] = 25'b1111101100101110110100000;
    rom[42024] = 25'b1111101100101110100000110;
    rom[42025] = 25'b1111101100101110001101110;
    rom[42026] = 25'b1111101100101101111010111;
    rom[42027] = 25'b1111101100101101101000001;
    rom[42028] = 25'b1111101100101101010101100;
    rom[42029] = 25'b1111101100101101000010111;
    rom[42030] = 25'b1111101100101100110000100;
    rom[42031] = 25'b1111101100101100011110001;
    rom[42032] = 25'b1111101100101100001100000;
    rom[42033] = 25'b1111101100101011111001111;
    rom[42034] = 25'b1111101100101011100111111;
    rom[42035] = 25'b1111101100101011010110001;
    rom[42036] = 25'b1111101100101011000100011;
    rom[42037] = 25'b1111101100101010110010101;
    rom[42038] = 25'b1111101100101010100001010;
    rom[42039] = 25'b1111101100101010001111111;
    rom[42040] = 25'b1111101100101001111110100;
    rom[42041] = 25'b1111101100101001101101011;
    rom[42042] = 25'b1111101100101001011100011;
    rom[42043] = 25'b1111101100101001001011100;
    rom[42044] = 25'b1111101100101000111010101;
    rom[42045] = 25'b1111101100101000101010000;
    rom[42046] = 25'b1111101100101000011001011;
    rom[42047] = 25'b1111101100101000001000111;
    rom[42048] = 25'b1111101100100111111000101;
    rom[42049] = 25'b1111101100100111101000011;
    rom[42050] = 25'b1111101100100111011000010;
    rom[42051] = 25'b1111101100100111001000010;
    rom[42052] = 25'b1111101100100110111000011;
    rom[42053] = 25'b1111101100100110101000101;
    rom[42054] = 25'b1111101100100110011001000;
    rom[42055] = 25'b1111101100100110001001011;
    rom[42056] = 25'b1111101100100101111010000;
    rom[42057] = 25'b1111101100100101101010110;
    rom[42058] = 25'b1111101100100101011011101;
    rom[42059] = 25'b1111101100100101001100100;
    rom[42060] = 25'b1111101100100100111101101;
    rom[42061] = 25'b1111101100100100101110110;
    rom[42062] = 25'b1111101100100100100000000;
    rom[42063] = 25'b1111101100100100010001011;
    rom[42064] = 25'b1111101100100100000010111;
    rom[42065] = 25'b1111101100100011110100100;
    rom[42066] = 25'b1111101100100011100110010;
    rom[42067] = 25'b1111101100100011011000001;
    rom[42068] = 25'b1111101100100011001010001;
    rom[42069] = 25'b1111101100100010111100001;
    rom[42070] = 25'b1111101100100010101110011;
    rom[42071] = 25'b1111101100100010100000110;
    rom[42072] = 25'b1111101100100010010011001;
    rom[42073] = 25'b1111101100100010000101101;
    rom[42074] = 25'b1111101100100001111000011;
    rom[42075] = 25'b1111101100100001101011001;
    rom[42076] = 25'b1111101100100001011110000;
    rom[42077] = 25'b1111101100100001010001000;
    rom[42078] = 25'b1111101100100001000100001;
    rom[42079] = 25'b1111101100100000110111011;
    rom[42080] = 25'b1111101100100000101010101;
    rom[42081] = 25'b1111101100100000011110001;
    rom[42082] = 25'b1111101100100000010001110;
    rom[42083] = 25'b1111101100100000000101011;
    rom[42084] = 25'b1111101100011111111001010;
    rom[42085] = 25'b1111101100011111101101010;
    rom[42086] = 25'b1111101100011111100001001;
    rom[42087] = 25'b1111101100011111010101011;
    rom[42088] = 25'b1111101100011111001001101;
    rom[42089] = 25'b1111101100011110111110000;
    rom[42090] = 25'b1111101100011110110010100;
    rom[42091] = 25'b1111101100011110100111001;
    rom[42092] = 25'b1111101100011110011011111;
    rom[42093] = 25'b1111101100011110010000101;
    rom[42094] = 25'b1111101100011110000101101;
    rom[42095] = 25'b1111101100011101111010110;
    rom[42096] = 25'b1111101100011101101111111;
    rom[42097] = 25'b1111101100011101100101001;
    rom[42098] = 25'b1111101100011101011010101;
    rom[42099] = 25'b1111101100011101010000001;
    rom[42100] = 25'b1111101100011101000101110;
    rom[42101] = 25'b1111101100011100111011100;
    rom[42102] = 25'b1111101100011100110001011;
    rom[42103] = 25'b1111101100011100100111011;
    rom[42104] = 25'b1111101100011100011101011;
    rom[42105] = 25'b1111101100011100010011101;
    rom[42106] = 25'b1111101100011100001010000;
    rom[42107] = 25'b1111101100011100000000011;
    rom[42108] = 25'b1111101100011011110111000;
    rom[42109] = 25'b1111101100011011101101101;
    rom[42110] = 25'b1111101100011011100100011;
    rom[42111] = 25'b1111101100011011011011010;
    rom[42112] = 25'b1111101100011011010010011;
    rom[42113] = 25'b1111101100011011001001011;
    rom[42114] = 25'b1111101100011011000000110;
    rom[42115] = 25'b1111101100011010111000000;
    rom[42116] = 25'b1111101100011010101111011;
    rom[42117] = 25'b1111101100011010100111000;
    rom[42118] = 25'b1111101100011010011110110;
    rom[42119] = 25'b1111101100011010010110100;
    rom[42120] = 25'b1111101100011010001110100;
    rom[42121] = 25'b1111101100011010000110011;
    rom[42122] = 25'b1111101100011001111110101;
    rom[42123] = 25'b1111101100011001110110111;
    rom[42124] = 25'b1111101100011001101111001;
    rom[42125] = 25'b1111101100011001100111110;
    rom[42126] = 25'b1111101100011001100000011;
    rom[42127] = 25'b1111101100011001011001000;
    rom[42128] = 25'b1111101100011001010001111;
    rom[42129] = 25'b1111101100011001001010110;
    rom[42130] = 25'b1111101100011001000011110;
    rom[42131] = 25'b1111101100011000111100111;
    rom[42132] = 25'b1111101100011000110110010;
    rom[42133] = 25'b1111101100011000101111101;
    rom[42134] = 25'b1111101100011000101001000;
    rom[42135] = 25'b1111101100011000100010101;
    rom[42136] = 25'b1111101100011000011100011;
    rom[42137] = 25'b1111101100011000010110010;
    rom[42138] = 25'b1111101100011000010000010;
    rom[42139] = 25'b1111101100011000001010010;
    rom[42140] = 25'b1111101100011000000100011;
    rom[42141] = 25'b1111101100010111111110110;
    rom[42142] = 25'b1111101100010111111001001;
    rom[42143] = 25'b1111101100010111110011101;
    rom[42144] = 25'b1111101100010111101110010;
    rom[42145] = 25'b1111101100010111101001000;
    rom[42146] = 25'b1111101100010111100011110;
    rom[42147] = 25'b1111101100010111011110110;
    rom[42148] = 25'b1111101100010111011001111;
    rom[42149] = 25'b1111101100010111010101000;
    rom[42150] = 25'b1111101100010111010000011;
    rom[42151] = 25'b1111101100010111001011101;
    rom[42152] = 25'b1111101100010111000111001;
    rom[42153] = 25'b1111101100010111000010111;
    rom[42154] = 25'b1111101100010110111110101;
    rom[42155] = 25'b1111101100010110111010100;
    rom[42156] = 25'b1111101100010110110110011;
    rom[42157] = 25'b1111101100010110110010011;
    rom[42158] = 25'b1111101100010110101110110;
    rom[42159] = 25'b1111101100010110101011000;
    rom[42160] = 25'b1111101100010110100111011;
    rom[42161] = 25'b1111101100010110100011111;
    rom[42162] = 25'b1111101100010110100000100;
    rom[42163] = 25'b1111101100010110011101010;
    rom[42164] = 25'b1111101100010110011010001;
    rom[42165] = 25'b1111101100010110010111001;
    rom[42166] = 25'b1111101100010110010100001;
    rom[42167] = 25'b1111101100010110010001011;
    rom[42168] = 25'b1111101100010110001110101;
    rom[42169] = 25'b1111101100010110001100000;
    rom[42170] = 25'b1111101100010110001001101;
    rom[42171] = 25'b1111101100010110000111010;
    rom[42172] = 25'b1111101100010110000101000;
    rom[42173] = 25'b1111101100010110000010110;
    rom[42174] = 25'b1111101100010110000000111;
    rom[42175] = 25'b1111101100010101111110111;
    rom[42176] = 25'b1111101100010101111101001;
    rom[42177] = 25'b1111101100010101111011011;
    rom[42178] = 25'b1111101100010101111001110;
    rom[42179] = 25'b1111101100010101111000011;
    rom[42180] = 25'b1111101100010101110111000;
    rom[42181] = 25'b1111101100010101110101101;
    rom[42182] = 25'b1111101100010101110100100;
    rom[42183] = 25'b1111101100010101110011100;
    rom[42184] = 25'b1111101100010101110010100;
    rom[42185] = 25'b1111101100010101110001110;
    rom[42186] = 25'b1111101100010101110001000;
    rom[42187] = 25'b1111101100010101110000100;
    rom[42188] = 25'b1111101100010101110000000;
    rom[42189] = 25'b1111101100010101101111101;
    rom[42190] = 25'b1111101100010101101111011;
    rom[42191] = 25'b1111101100010101101111010;
    rom[42192] = 25'b1111101100010101101111001;
    rom[42193] = 25'b1111101100010101101111010;
    rom[42194] = 25'b1111101100010101101111011;
    rom[42195] = 25'b1111101100010101101111101;
    rom[42196] = 25'b1111101100010101110000000;
    rom[42197] = 25'b1111101100010101110000101;
    rom[42198] = 25'b1111101100010101110001001;
    rom[42199] = 25'b1111101100010101110001111;
    rom[42200] = 25'b1111101100010101110010110;
    rom[42201] = 25'b1111101100010101110011101;
    rom[42202] = 25'b1111101100010101110100110;
    rom[42203] = 25'b1111101100010101110101111;
    rom[42204] = 25'b1111101100010101110111010;
    rom[42205] = 25'b1111101100010101111000101;
    rom[42206] = 25'b1111101100010101111010001;
    rom[42207] = 25'b1111101100010101111011110;
    rom[42208] = 25'b1111101100010101111101011;
    rom[42209] = 25'b1111101100010101111111010;
    rom[42210] = 25'b1111101100010110000001001;
    rom[42211] = 25'b1111101100010110000011001;
    rom[42212] = 25'b1111101100010110000101011;
    rom[42213] = 25'b1111101100010110000111101;
    rom[42214] = 25'b1111101100010110001010000;
    rom[42215] = 25'b1111101100010110001100011;
    rom[42216] = 25'b1111101100010110001111000;
    rom[42217] = 25'b1111101100010110010001110;
    rom[42218] = 25'b1111101100010110010100100;
    rom[42219] = 25'b1111101100010110010111100;
    rom[42220] = 25'b1111101100010110011010011;
    rom[42221] = 25'b1111101100010110011101101;
    rom[42222] = 25'b1111101100010110100000110;
    rom[42223] = 25'b1111101100010110100100001;
    rom[42224] = 25'b1111101100010110100111101;
    rom[42225] = 25'b1111101100010110101011001;
    rom[42226] = 25'b1111101100010110101110110;
    rom[42227] = 25'b1111101100010110110010101;
    rom[42228] = 25'b1111101100010110110110100;
    rom[42229] = 25'b1111101100010110111010100;
    rom[42230] = 25'b1111101100010110111110101;
    rom[42231] = 25'b1111101100010111000010110;
    rom[42232] = 25'b1111101100010111000111001;
    rom[42233] = 25'b1111101100010111001011100;
    rom[42234] = 25'b1111101100010111010000000;
    rom[42235] = 25'b1111101100010111010100110;
    rom[42236] = 25'b1111101100010111011001100;
    rom[42237] = 25'b1111101100010111011110011;
    rom[42238] = 25'b1111101100010111100011010;
    rom[42239] = 25'b1111101100010111101000011;
    rom[42240] = 25'b1111101100010111101101100;
    rom[42241] = 25'b1111101100010111110010111;
    rom[42242] = 25'b1111101100010111111000010;
    rom[42243] = 25'b1111101100010111111101110;
    rom[42244] = 25'b1111101100011000000011010;
    rom[42245] = 25'b1111101100011000001001001;
    rom[42246] = 25'b1111101100011000001110111;
    rom[42247] = 25'b1111101100011000010100110;
    rom[42248] = 25'b1111101100011000011010111;
    rom[42249] = 25'b1111101100011000100001000;
    rom[42250] = 25'b1111101100011000100111010;
    rom[42251] = 25'b1111101100011000101101101;
    rom[42252] = 25'b1111101100011000110100000;
    rom[42253] = 25'b1111101100011000111010101;
    rom[42254] = 25'b1111101100011001000001010;
    rom[42255] = 25'b1111101100011001001000001;
    rom[42256] = 25'b1111101100011001001111000;
    rom[42257] = 25'b1111101100011001010110000;
    rom[42258] = 25'b1111101100011001011101001;
    rom[42259] = 25'b1111101100011001100100011;
    rom[42260] = 25'b1111101100011001101011101;
    rom[42261] = 25'b1111101100011001110011001;
    rom[42262] = 25'b1111101100011001111010101;
    rom[42263] = 25'b1111101100011010000010010;
    rom[42264] = 25'b1111101100011010001010000;
    rom[42265] = 25'b1111101100011010010001110;
    rom[42266] = 25'b1111101100011010011001111;
    rom[42267] = 25'b1111101100011010100001111;
    rom[42268] = 25'b1111101100011010101010000;
    rom[42269] = 25'b1111101100011010110010010;
    rom[42270] = 25'b1111101100011010111010110;
    rom[42271] = 25'b1111101100011011000011010;
    rom[42272] = 25'b1111101100011011001011110;
    rom[42273] = 25'b1111101100011011010100100;
    rom[42274] = 25'b1111101100011011011101010;
    rom[42275] = 25'b1111101100011011100110001;
    rom[42276] = 25'b1111101100011011101111010;
    rom[42277] = 25'b1111101100011011111000011;
    rom[42278] = 25'b1111101100011100000001100;
    rom[42279] = 25'b1111101100011100001010111;
    rom[42280] = 25'b1111101100011100010100010;
    rom[42281] = 25'b1111101100011100011101110;
    rom[42282] = 25'b1111101100011100100111100;
    rom[42283] = 25'b1111101100011100110001010;
    rom[42284] = 25'b1111101100011100111011001;
    rom[42285] = 25'b1111101100011101000101000;
    rom[42286] = 25'b1111101100011101001111001;
    rom[42287] = 25'b1111101100011101011001010;
    rom[42288] = 25'b1111101100011101100011100;
    rom[42289] = 25'b1111101100011101101101111;
    rom[42290] = 25'b1111101100011101111000100;
    rom[42291] = 25'b1111101100011110000011000;
    rom[42292] = 25'b1111101100011110001101101;
    rom[42293] = 25'b1111101100011110011000100;
    rom[42294] = 25'b1111101100011110100011011;
    rom[42295] = 25'b1111101100011110101110100;
    rom[42296] = 25'b1111101100011110111001101;
    rom[42297] = 25'b1111101100011111000100110;
    rom[42298] = 25'b1111101100011111010000001;
    rom[42299] = 25'b1111101100011111011011100;
    rom[42300] = 25'b1111101100011111100111000;
    rom[42301] = 25'b1111101100011111110010101;
    rom[42302] = 25'b1111101100011111111110011;
    rom[42303] = 25'b1111101100100000001010010;
    rom[42304] = 25'b1111101100100000010110010;
    rom[42305] = 25'b1111101100100000100010010;
    rom[42306] = 25'b1111101100100000101110011;
    rom[42307] = 25'b1111101100100000111010101;
    rom[42308] = 25'b1111101100100001000111000;
    rom[42309] = 25'b1111101100100001010011100;
    rom[42310] = 25'b1111101100100001100000000;
    rom[42311] = 25'b1111101100100001101100101;
    rom[42312] = 25'b1111101100100001111001100;
    rom[42313] = 25'b1111101100100010000110010;
    rom[42314] = 25'b1111101100100010010011010;
    rom[42315] = 25'b1111101100100010100000011;
    rom[42316] = 25'b1111101100100010101101101;
    rom[42317] = 25'b1111101100100010111010111;
    rom[42318] = 25'b1111101100100011001000010;
    rom[42319] = 25'b1111101100100011010101110;
    rom[42320] = 25'b1111101100100011100011010;
    rom[42321] = 25'b1111101100100011110001000;
    rom[42322] = 25'b1111101100100011111110111;
    rom[42323] = 25'b1111101100100100001100110;
    rom[42324] = 25'b1111101100100100011010110;
    rom[42325] = 25'b1111101100100100101000111;
    rom[42326] = 25'b1111101100100100110111000;
    rom[42327] = 25'b1111101100100101000101011;
    rom[42328] = 25'b1111101100100101010011110;
    rom[42329] = 25'b1111101100100101100010010;
    rom[42330] = 25'b1111101100100101110000111;
    rom[42331] = 25'b1111101100100101111111101;
    rom[42332] = 25'b1111101100100110001110100;
    rom[42333] = 25'b1111101100100110011101011;
    rom[42334] = 25'b1111101100100110101100011;
    rom[42335] = 25'b1111101100100110111011100;
    rom[42336] = 25'b1111101100100111001010110;
    rom[42337] = 25'b1111101100100111011010001;
    rom[42338] = 25'b1111101100100111101001100;
    rom[42339] = 25'b1111101100100111111001000;
    rom[42340] = 25'b1111101100101000001000110;
    rom[42341] = 25'b1111101100101000011000011;
    rom[42342] = 25'b1111101100101000101000010;
    rom[42343] = 25'b1111101100101000111000001;
    rom[42344] = 25'b1111101100101001001000010;
    rom[42345] = 25'b1111101100101001011000011;
    rom[42346] = 25'b1111101100101001101000101;
    rom[42347] = 25'b1111101100101001111001000;
    rom[42348] = 25'b1111101100101010001001011;
    rom[42349] = 25'b1111101100101010011001111;
    rom[42350] = 25'b1111101100101010101010100;
    rom[42351] = 25'b1111101100101010111011011;
    rom[42352] = 25'b1111101100101011001100001;
    rom[42353] = 25'b1111101100101011011101001;
    rom[42354] = 25'b1111101100101011101110001;
    rom[42355] = 25'b1111101100101011111111011;
    rom[42356] = 25'b1111101100101100010000101;
    rom[42357] = 25'b1111101100101100100001111;
    rom[42358] = 25'b1111101100101100110011011;
    rom[42359] = 25'b1111101100101101000100111;
    rom[42360] = 25'b1111101100101101010110101;
    rom[42361] = 25'b1111101100101101101000010;
    rom[42362] = 25'b1111101100101101111010001;
    rom[42363] = 25'b1111101100101110001100001;
    rom[42364] = 25'b1111101100101110011110010;
    rom[42365] = 25'b1111101100101110110000010;
    rom[42366] = 25'b1111101100101111000010100;
    rom[42367] = 25'b1111101100101111010100111;
    rom[42368] = 25'b1111101100101111100111011;
    rom[42369] = 25'b1111101100101111111001111;
    rom[42370] = 25'b1111101100110000001100101;
    rom[42371] = 25'b1111101100110000011111010;
    rom[42372] = 25'b1111101100110000110010001;
    rom[42373] = 25'b1111101100110001000101001;
    rom[42374] = 25'b1111101100110001011000001;
    rom[42375] = 25'b1111101100110001101011010;
    rom[42376] = 25'b1111101100110001111110100;
    rom[42377] = 25'b1111101100110010010001111;
    rom[42378] = 25'b1111101100110010100101010;
    rom[42379] = 25'b1111101100110010111000110;
    rom[42380] = 25'b1111101100110011001100100;
    rom[42381] = 25'b1111101100110011100000010;
    rom[42382] = 25'b1111101100110011110100000;
    rom[42383] = 25'b1111101100110100001000000;
    rom[42384] = 25'b1111101100110100011100000;
    rom[42385] = 25'b1111101100110100110000001;
    rom[42386] = 25'b1111101100110101000100010;
    rom[42387] = 25'b1111101100110101011000101;
    rom[42388] = 25'b1111101100110101101101001;
    rom[42389] = 25'b1111101100110110000001101;
    rom[42390] = 25'b1111101100110110010110010;
    rom[42391] = 25'b1111101100110110101010111;
    rom[42392] = 25'b1111101100110110111111110;
    rom[42393] = 25'b1111101100110111010100101;
    rom[42394] = 25'b1111101100110111101001110;
    rom[42395] = 25'b1111101100110111111110110;
    rom[42396] = 25'b1111101100111000010100000;
    rom[42397] = 25'b1111101100111000101001010;
    rom[42398] = 25'b1111101100111000111110101;
    rom[42399] = 25'b1111101100111001010100001;
    rom[42400] = 25'b1111101100111001101001110;
    rom[42401] = 25'b1111101100111001111111100;
    rom[42402] = 25'b1111101100111010010101010;
    rom[42403] = 25'b1111101100111010101011001;
    rom[42404] = 25'b1111101100111011000001001;
    rom[42405] = 25'b1111101100111011010111001;
    rom[42406] = 25'b1111101100111011101101010;
    rom[42407] = 25'b1111101100111100000011101;
    rom[42408] = 25'b1111101100111100011010000;
    rom[42409] = 25'b1111101100111100110000100;
    rom[42410] = 25'b1111101100111101000111000;
    rom[42411] = 25'b1111101100111101011101101;
    rom[42412] = 25'b1111101100111101110100100;
    rom[42413] = 25'b1111101100111110001011010;
    rom[42414] = 25'b1111101100111110100010010;
    rom[42415] = 25'b1111101100111110111001010;
    rom[42416] = 25'b1111101100111111010000011;
    rom[42417] = 25'b1111101100111111100111101;
    rom[42418] = 25'b1111101100111111111110111;
    rom[42419] = 25'b1111101101000000010110011;
    rom[42420] = 25'b1111101101000000101101111;
    rom[42421] = 25'b1111101101000001000101100;
    rom[42422] = 25'b1111101101000001011101010;
    rom[42423] = 25'b1111101101000001110101001;
    rom[42424] = 25'b1111101101000010001101000;
    rom[42425] = 25'b1111101101000010100101000;
    rom[42426] = 25'b1111101101000010111101001;
    rom[42427] = 25'b1111101101000011010101010;
    rom[42428] = 25'b1111101101000011101101100;
    rom[42429] = 25'b1111101101000100000101111;
    rom[42430] = 25'b1111101101000100011110011;
    rom[42431] = 25'b1111101101000100110111000;
    rom[42432] = 25'b1111101101000101001111101;
    rom[42433] = 25'b1111101101000101101000011;
    rom[42434] = 25'b1111101101000110000001001;
    rom[42435] = 25'b1111101101000110011010001;
    rom[42436] = 25'b1111101101000110110011001;
    rom[42437] = 25'b1111101101000111001100011;
    rom[42438] = 25'b1111101101000111100101101;
    rom[42439] = 25'b1111101101000111111110111;
    rom[42440] = 25'b1111101101001000011000010;
    rom[42441] = 25'b1111101101001000110001110;
    rom[42442] = 25'b1111101101001001001011100;
    rom[42443] = 25'b1111101101001001100101001;
    rom[42444] = 25'b1111101101001001111110111;
    rom[42445] = 25'b1111101101001010011000110;
    rom[42446] = 25'b1111101101001010110010110;
    rom[42447] = 25'b1111101101001011001100111;
    rom[42448] = 25'b1111101101001011100111000;
    rom[42449] = 25'b1111101101001100000001010;
    rom[42450] = 25'b1111101101001100011011101;
    rom[42451] = 25'b1111101101001100110110001;
    rom[42452] = 25'b1111101101001101010000101;
    rom[42453] = 25'b1111101101001101101011010;
    rom[42454] = 25'b1111101101001110000110000;
    rom[42455] = 25'b1111101101001110100000110;
    rom[42456] = 25'b1111101101001110111011110;
    rom[42457] = 25'b1111101101001111010110110;
    rom[42458] = 25'b1111101101001111110001111;
    rom[42459] = 25'b1111101101010000001101000;
    rom[42460] = 25'b1111101101010000101000010;
    rom[42461] = 25'b1111101101010001000011110;
    rom[42462] = 25'b1111101101010001011111010;
    rom[42463] = 25'b1111101101010001111010110;
    rom[42464] = 25'b1111101101010010010110011;
    rom[42465] = 25'b1111101101010010110010001;
    rom[42466] = 25'b1111101101010011001110000;
    rom[42467] = 25'b1111101101010011101001111;
    rom[42468] = 25'b1111101101010100000101111;
    rom[42469] = 25'b1111101101010100100010000;
    rom[42470] = 25'b1111101101010100111110010;
    rom[42471] = 25'b1111101101010101011010100;
    rom[42472] = 25'b1111101101010101110110111;
    rom[42473] = 25'b1111101101010110010011011;
    rom[42474] = 25'b1111101101010110110000000;
    rom[42475] = 25'b1111101101010111001100101;
    rom[42476] = 25'b1111101101010111101001011;
    rom[42477] = 25'b1111101101011000000110010;
    rom[42478] = 25'b1111101101011000100011010;
    rom[42479] = 25'b1111101101011001000000010;
    rom[42480] = 25'b1111101101011001011101011;
    rom[42481] = 25'b1111101101011001111010101;
    rom[42482] = 25'b1111101101011010010111111;
    rom[42483] = 25'b1111101101011010110101010;
    rom[42484] = 25'b1111101101011011010010110;
    rom[42485] = 25'b1111101101011011110000011;
    rom[42486] = 25'b1111101101011100001110000;
    rom[42487] = 25'b1111101101011100101011110;
    rom[42488] = 25'b1111101101011101001001100;
    rom[42489] = 25'b1111101101011101100111100;
    rom[42490] = 25'b1111101101011110000101100;
    rom[42491] = 25'b1111101101011110100011101;
    rom[42492] = 25'b1111101101011111000001111;
    rom[42493] = 25'b1111101101011111100000001;
    rom[42494] = 25'b1111101101011111111110100;
    rom[42495] = 25'b1111101101100000011101001;
    rom[42496] = 25'b1111101101100000111011101;
    rom[42497] = 25'b1111101101100001011010010;
    rom[42498] = 25'b1111101101100001111001000;
    rom[42499] = 25'b1111101101100010010111111;
    rom[42500] = 25'b1111101101100010110110110;
    rom[42501] = 25'b1111101101100011010101110;
    rom[42502] = 25'b1111101101100011110100111;
    rom[42503] = 25'b1111101101100100010100001;
    rom[42504] = 25'b1111101101100100110011011;
    rom[42505] = 25'b1111101101100101010010110;
    rom[42506] = 25'b1111101101100101110010001;
    rom[42507] = 25'b1111101101100110010001101;
    rom[42508] = 25'b1111101101100110110001011;
    rom[42509] = 25'b1111101101100111010001001;
    rom[42510] = 25'b1111101101100111110000111;
    rom[42511] = 25'b1111101101101000010000110;
    rom[42512] = 25'b1111101101101000110000111;
    rom[42513] = 25'b1111101101101001010000111;
    rom[42514] = 25'b1111101101101001110001000;
    rom[42515] = 25'b1111101101101010010001010;
    rom[42516] = 25'b1111101101101010110001101;
    rom[42517] = 25'b1111101101101011010010000;
    rom[42518] = 25'b1111101101101011110010101;
    rom[42519] = 25'b1111101101101100010011010;
    rom[42520] = 25'b1111101101101100110011111;
    rom[42521] = 25'b1111101101101101010100101;
    rom[42522] = 25'b1111101101101101110101100;
    rom[42523] = 25'b1111101101101110010110100;
    rom[42524] = 25'b1111101101101110110111100;
    rom[42525] = 25'b1111101101101111011000101;
    rom[42526] = 25'b1111101101101111111001111;
    rom[42527] = 25'b1111101101110000011011010;
    rom[42528] = 25'b1111101101110000111100100;
    rom[42529] = 25'b1111101101110001011110000;
    rom[42530] = 25'b1111101101110001111111101;
    rom[42531] = 25'b1111101101110010100001010;
    rom[42532] = 25'b1111101101110011000011000;
    rom[42533] = 25'b1111101101110011100100111;
    rom[42534] = 25'b1111101101110100000110110;
    rom[42535] = 25'b1111101101110100101000110;
    rom[42536] = 25'b1111101101110101001010110;
    rom[42537] = 25'b1111101101110101101101000;
    rom[42538] = 25'b1111101101110110001111010;
    rom[42539] = 25'b1111101101110110110001101;
    rom[42540] = 25'b1111101101110111010100000;
    rom[42541] = 25'b1111101101110111110110100;
    rom[42542] = 25'b1111101101111000011001001;
    rom[42543] = 25'b1111101101111000111011111;
    rom[42544] = 25'b1111101101111001011110101;
    rom[42545] = 25'b1111101101111010000001011;
    rom[42546] = 25'b1111101101111010100100011;
    rom[42547] = 25'b1111101101111011000111100;
    rom[42548] = 25'b1111101101111011101010100;
    rom[42549] = 25'b1111101101111100001101110;
    rom[42550] = 25'b1111101101111100110001000;
    rom[42551] = 25'b1111101101111101010100011;
    rom[42552] = 25'b1111101101111101110111111;
    rom[42553] = 25'b1111101101111110011011011;
    rom[42554] = 25'b1111101101111110111111000;
    rom[42555] = 25'b1111101101111111100010101;
    rom[42556] = 25'b1111101110000000000110100;
    rom[42557] = 25'b1111101110000000101010011;
    rom[42558] = 25'b1111101110000001001110011;
    rom[42559] = 25'b1111101110000001110010011;
    rom[42560] = 25'b1111101110000010010110100;
    rom[42561] = 25'b1111101110000010111010101;
    rom[42562] = 25'b1111101110000011011111000;
    rom[42563] = 25'b1111101110000100000011011;
    rom[42564] = 25'b1111101110000100100111111;
    rom[42565] = 25'b1111101110000101001100100;
    rom[42566] = 25'b1111101110000101110001001;
    rom[42567] = 25'b1111101110000110010101110;
    rom[42568] = 25'b1111101110000110111010101;
    rom[42569] = 25'b1111101110000111011111100;
    rom[42570] = 25'b1111101110001000000100011;
    rom[42571] = 25'b1111101110001000101001100;
    rom[42572] = 25'b1111101110001001001110101;
    rom[42573] = 25'b1111101110001001110011111;
    rom[42574] = 25'b1111101110001010011001001;
    rom[42575] = 25'b1111101110001010111110100;
    rom[42576] = 25'b1111101110001011100100000;
    rom[42577] = 25'b1111101110001100001001100;
    rom[42578] = 25'b1111101110001100101111001;
    rom[42579] = 25'b1111101110001101010100111;
    rom[42580] = 25'b1111101110001101111010101;
    rom[42581] = 25'b1111101110001110100000100;
    rom[42582] = 25'b1111101110001111000110100;
    rom[42583] = 25'b1111101110001111101100101;
    rom[42584] = 25'b1111101110010000010010101;
    rom[42585] = 25'b1111101110010000111000111;
    rom[42586] = 25'b1111101110010001011111001;
    rom[42587] = 25'b1111101110010010000101100;
    rom[42588] = 25'b1111101110010010101100000;
    rom[42589] = 25'b1111101110010011010010101;
    rom[42590] = 25'b1111101110010011111001001;
    rom[42591] = 25'b1111101110010100011111111;
    rom[42592] = 25'b1111101110010101000110101;
    rom[42593] = 25'b1111101110010101101101100;
    rom[42594] = 25'b1111101110010110010100100;
    rom[42595] = 25'b1111101110010110111011100;
    rom[42596] = 25'b1111101110010111100010100;
    rom[42597] = 25'b1111101110011000001001110;
    rom[42598] = 25'b1111101110011000110001001;
    rom[42599] = 25'b1111101110011001011000011;
    rom[42600] = 25'b1111101110011001111111110;
    rom[42601] = 25'b1111101110011010100111010;
    rom[42602] = 25'b1111101110011011001110111;
    rom[42603] = 25'b1111101110011011110110101;
    rom[42604] = 25'b1111101110011100011110010;
    rom[42605] = 25'b1111101110011101000110001;
    rom[42606] = 25'b1111101110011101101110000;
    rom[42607] = 25'b1111101110011110010110001;
    rom[42608] = 25'b1111101110011110111110001;
    rom[42609] = 25'b1111101110011111100110010;
    rom[42610] = 25'b1111101110100000001110100;
    rom[42611] = 25'b1111101110100000110110110;
    rom[42612] = 25'b1111101110100001011111001;
    rom[42613] = 25'b1111101110100010000111101;
    rom[42614] = 25'b1111101110100010110000010;
    rom[42615] = 25'b1111101110100011011000111;
    rom[42616] = 25'b1111101110100100000001100;
    rom[42617] = 25'b1111101110100100101010011;
    rom[42618] = 25'b1111101110100101010011001;
    rom[42619] = 25'b1111101110100101111100001;
    rom[42620] = 25'b1111101110100110100101001;
    rom[42621] = 25'b1111101110100111001110010;
    rom[42622] = 25'b1111101110100111110111011;
    rom[42623] = 25'b1111101110101000100000110;
    rom[42624] = 25'b1111101110101001001010000;
    rom[42625] = 25'b1111101110101001110011100;
    rom[42626] = 25'b1111101110101010011100111;
    rom[42627] = 25'b1111101110101011000110100;
    rom[42628] = 25'b1111101110101011110000001;
    rom[42629] = 25'b1111101110101100011001111;
    rom[42630] = 25'b1111101110101101000011110;
    rom[42631] = 25'b1111101110101101101101100;
    rom[42632] = 25'b1111101110101110010111101;
    rom[42633] = 25'b1111101110101111000001101;
    rom[42634] = 25'b1111101110101111101011110;
    rom[42635] = 25'b1111101110110000010101111;
    rom[42636] = 25'b1111101110110001000000001;
    rom[42637] = 25'b1111101110110001101010100;
    rom[42638] = 25'b1111101110110010010100111;
    rom[42639] = 25'b1111101110110010111111011;
    rom[42640] = 25'b1111101110110011101010000;
    rom[42641] = 25'b1111101110110100010100101;
    rom[42642] = 25'b1111101110110100111111011;
    rom[42643] = 25'b1111101110110101101010010;
    rom[42644] = 25'b1111101110110110010101001;
    rom[42645] = 25'b1111101110110111000000000;
    rom[42646] = 25'b1111101110110111101011001;
    rom[42647] = 25'b1111101110111000010110010;
    rom[42648] = 25'b1111101110111001000001011;
    rom[42649] = 25'b1111101110111001101100101;
    rom[42650] = 25'b1111101110111010011000000;
    rom[42651] = 25'b1111101110111011000011011;
    rom[42652] = 25'b1111101110111011101110111;
    rom[42653] = 25'b1111101110111100011010100;
    rom[42654] = 25'b1111101110111101000110001;
    rom[42655] = 25'b1111101110111101110001111;
    rom[42656] = 25'b1111101110111110011101101;
    rom[42657] = 25'b1111101110111111001001100;
    rom[42658] = 25'b1111101110111111110101100;
    rom[42659] = 25'b1111101111000000100001100;
    rom[42660] = 25'b1111101111000001001101101;
    rom[42661] = 25'b1111101111000001111001111;
    rom[42662] = 25'b1111101111000010100110000;
    rom[42663] = 25'b1111101111000011010010011;
    rom[42664] = 25'b1111101111000011111110110;
    rom[42665] = 25'b1111101111000100101011010;
    rom[42666] = 25'b1111101111000101010111110;
    rom[42667] = 25'b1111101111000110000100100;
    rom[42668] = 25'b1111101111000110110001001;
    rom[42669] = 25'b1111101111000111011101111;
    rom[42670] = 25'b1111101111001000001010110;
    rom[42671] = 25'b1111101111001000110111101;
    rom[42672] = 25'b1111101111001001100100101;
    rom[42673] = 25'b1111101111001010010001101;
    rom[42674] = 25'b1111101111001010111110111;
    rom[42675] = 25'b1111101111001011101100001;
    rom[42676] = 25'b1111101111001100011001011;
    rom[42677] = 25'b1111101111001101000110101;
    rom[42678] = 25'b1111101111001101110100001;
    rom[42679] = 25'b1111101111001110100001101;
    rom[42680] = 25'b1111101111001111001111010;
    rom[42681] = 25'b1111101111001111111100111;
    rom[42682] = 25'b1111101111010000101010101;
    rom[42683] = 25'b1111101111010001011000011;
    rom[42684] = 25'b1111101111010010000110011;
    rom[42685] = 25'b1111101111010010110100010;
    rom[42686] = 25'b1111101111010011100010010;
    rom[42687] = 25'b1111101111010100010000011;
    rom[42688] = 25'b1111101111010100111110100;
    rom[42689] = 25'b1111101111010101101100110;
    rom[42690] = 25'b1111101111010110011011000;
    rom[42691] = 25'b1111101111010111001001100;
    rom[42692] = 25'b1111101111010111110111111;
    rom[42693] = 25'b1111101111011000100110100;
    rom[42694] = 25'b1111101111011001010101001;
    rom[42695] = 25'b1111101111011010000011101;
    rom[42696] = 25'b1111101111011010110010100;
    rom[42697] = 25'b1111101111011011100001010;
    rom[42698] = 25'b1111101111011100010000001;
    rom[42699] = 25'b1111101111011100111111001;
    rom[42700] = 25'b1111101111011101101110001;
    rom[42701] = 25'b1111101111011110011101010;
    rom[42702] = 25'b1111101111011111001100011;
    rom[42703] = 25'b1111101111011111111011101;
    rom[42704] = 25'b1111101111100000101010111;
    rom[42705] = 25'b1111101111100001011010011;
    rom[42706] = 25'b1111101111100010001001110;
    rom[42707] = 25'b1111101111100010111001010;
    rom[42708] = 25'b1111101111100011101000111;
    rom[42709] = 25'b1111101111100100011000101;
    rom[42710] = 25'b1111101111100101001000010;
    rom[42711] = 25'b1111101111100101111000001;
    rom[42712] = 25'b1111101111100110100111111;
    rom[42713] = 25'b1111101111100111010111111;
    rom[42714] = 25'b1111101111101000000111111;
    rom[42715] = 25'b1111101111101000111000000;
    rom[42716] = 25'b1111101111101001101000001;
    rom[42717] = 25'b1111101111101010011000011;
    rom[42718] = 25'b1111101111101011001000101;
    rom[42719] = 25'b1111101111101011111001000;
    rom[42720] = 25'b1111101111101100101001011;
    rom[42721] = 25'b1111101111101101011010000;
    rom[42722] = 25'b1111101111101110001010100;
    rom[42723] = 25'b1111101111101110111011010;
    rom[42724] = 25'b1111101111101111101011111;
    rom[42725] = 25'b1111101111110000011100110;
    rom[42726] = 25'b1111101111110001001101100;
    rom[42727] = 25'b1111101111110001111110011;
    rom[42728] = 25'b1111101111110010101111011;
    rom[42729] = 25'b1111101111110011100000011;
    rom[42730] = 25'b1111101111110100010001100;
    rom[42731] = 25'b1111101111110101000010110;
    rom[42732] = 25'b1111101111110101110100000;
    rom[42733] = 25'b1111101111110110100101011;
    rom[42734] = 25'b1111101111110111010110110;
    rom[42735] = 25'b1111101111111000001000001;
    rom[42736] = 25'b1111101111111000111001101;
    rom[42737] = 25'b1111101111111001101011010;
    rom[42738] = 25'b1111101111111010011101000;
    rom[42739] = 25'b1111101111111011001110110;
    rom[42740] = 25'b1111101111111100000000100;
    rom[42741] = 25'b1111101111111100110010011;
    rom[42742] = 25'b1111101111111101100100011;
    rom[42743] = 25'b1111101111111110010110010;
    rom[42744] = 25'b1111101111111111001000011;
    rom[42745] = 25'b1111101111111111111010100;
    rom[42746] = 25'b1111110000000000101100110;
    rom[42747] = 25'b1111110000000001011111000;
    rom[42748] = 25'b1111110000000010010001011;
    rom[42749] = 25'b1111110000000011000011110;
    rom[42750] = 25'b1111110000000011110110001;
    rom[42751] = 25'b1111110000000100101000110;
    rom[42752] = 25'b1111110000000101011011011;
    rom[42753] = 25'b1111110000000110001101111;
    rom[42754] = 25'b1111110000000111000000110;
    rom[42755] = 25'b1111110000000111110011100;
    rom[42756] = 25'b1111110000001000100110011;
    rom[42757] = 25'b1111110000001001011001011;
    rom[42758] = 25'b1111110000001010001100011;
    rom[42759] = 25'b1111110000001010111111010;
    rom[42760] = 25'b1111110000001011110010100;
    rom[42761] = 25'b1111110000001100100101101;
    rom[42762] = 25'b1111110000001101011000111;
    rom[42763] = 25'b1111110000001110001100010;
    rom[42764] = 25'b1111110000001110111111101;
    rom[42765] = 25'b1111110000001111110011001;
    rom[42766] = 25'b1111110000010000100110101;
    rom[42767] = 25'b1111110000010001011010001;
    rom[42768] = 25'b1111110000010010001101110;
    rom[42769] = 25'b1111110000010011000001100;
    rom[42770] = 25'b1111110000010011110101011;
    rom[42771] = 25'b1111110000010100101001001;
    rom[42772] = 25'b1111110000010101011101000;
    rom[42773] = 25'b1111110000010110010001000;
    rom[42774] = 25'b1111110000010111000101000;
    rom[42775] = 25'b1111110000010111111001001;
    rom[42776] = 25'b1111110000011000101101010;
    rom[42777] = 25'b1111110000011001100001100;
    rom[42778] = 25'b1111110000011010010101110;
    rom[42779] = 25'b1111110000011011001010001;
    rom[42780] = 25'b1111110000011011111110100;
    rom[42781] = 25'b1111110000011100110011000;
    rom[42782] = 25'b1111110000011101100111101;
    rom[42783] = 25'b1111110000011110011100001;
    rom[42784] = 25'b1111110000011111010000111;
    rom[42785] = 25'b1111110000100000000101100;
    rom[42786] = 25'b1111110000100000111010011;
    rom[42787] = 25'b1111110000100001101111010;
    rom[42788] = 25'b1111110000100010100100001;
    rom[42789] = 25'b1111110000100011011001001;
    rom[42790] = 25'b1111110000100100001110001;
    rom[42791] = 25'b1111110000100101000011010;
    rom[42792] = 25'b1111110000100101111000011;
    rom[42793] = 25'b1111110000100110101101101;
    rom[42794] = 25'b1111110000100111100010111;
    rom[42795] = 25'b1111110000101000011000010;
    rom[42796] = 25'b1111110000101001001101101;
    rom[42797] = 25'b1111110000101010000011001;
    rom[42798] = 25'b1111110000101010111000101;
    rom[42799] = 25'b1111110000101011101110010;
    rom[42800] = 25'b1111110000101100100100000;
    rom[42801] = 25'b1111110000101101011001101;
    rom[42802] = 25'b1111110000101110001111100;
    rom[42803] = 25'b1111110000101111000101010;
    rom[42804] = 25'b1111110000101111111011010;
    rom[42805] = 25'b1111110000110000110001001;
    rom[42806] = 25'b1111110000110001100111001;
    rom[42807] = 25'b1111110000110010011101010;
    rom[42808] = 25'b1111110000110011010011011;
    rom[42809] = 25'b1111110000110100001001101;
    rom[42810] = 25'b1111110000110100111111111;
    rom[42811] = 25'b1111110000110101110110001;
    rom[42812] = 25'b1111110000110110101100100;
    rom[42813] = 25'b1111110000110111100011000;
    rom[42814] = 25'b1111110000111000011001100;
    rom[42815] = 25'b1111110000111001010000000;
    rom[42816] = 25'b1111110000111010000110101;
    rom[42817] = 25'b1111110000111010111101011;
    rom[42818] = 25'b1111110000111011110100001;
    rom[42819] = 25'b1111110000111100101011000;
    rom[42820] = 25'b1111110000111101100001111;
    rom[42821] = 25'b1111110000111110011000110;
    rom[42822] = 25'b1111110000111111001111101;
    rom[42823] = 25'b1111110001000000000110110;
    rom[42824] = 25'b1111110001000000111101111;
    rom[42825] = 25'b1111110001000001110101000;
    rom[42826] = 25'b1111110001000010101100010;
    rom[42827] = 25'b1111110001000011100011100;
    rom[42828] = 25'b1111110001000100011010111;
    rom[42829] = 25'b1111110001000101010010010;
    rom[42830] = 25'b1111110001000110001001101;
    rom[42831] = 25'b1111110001000111000001010;
    rom[42832] = 25'b1111110001000111111000111;
    rom[42833] = 25'b1111110001001000110000011;
    rom[42834] = 25'b1111110001001001101000000;
    rom[42835] = 25'b1111110001001010011111110;
    rom[42836] = 25'b1111110001001011010111101;
    rom[42837] = 25'b1111110001001100001111100;
    rom[42838] = 25'b1111110001001101000111011;
    rom[42839] = 25'b1111110001001101111111011;
    rom[42840] = 25'b1111110001001110110111011;
    rom[42841] = 25'b1111110001001111101111100;
    rom[42842] = 25'b1111110001010000100111101;
    rom[42843] = 25'b1111110001010001011111111;
    rom[42844] = 25'b1111110001010010011000001;
    rom[42845] = 25'b1111110001010011010000011;
    rom[42846] = 25'b1111110001010100001000110;
    rom[42847] = 25'b1111110001010101000001010;
    rom[42848] = 25'b1111110001010101111001110;
    rom[42849] = 25'b1111110001010110110010010;
    rom[42850] = 25'b1111110001010111101010110;
    rom[42851] = 25'b1111110001011000100011100;
    rom[42852] = 25'b1111110001011001011100001;
    rom[42853] = 25'b1111110001011010010101000;
    rom[42854] = 25'b1111110001011011001101110;
    rom[42855] = 25'b1111110001011100000110101;
    rom[42856] = 25'b1111110001011100111111101;
    rom[42857] = 25'b1111110001011101111000100;
    rom[42858] = 25'b1111110001011110110001101;
    rom[42859] = 25'b1111110001011111101010101;
    rom[42860] = 25'b1111110001100000100011110;
    rom[42861] = 25'b1111110001100001011101000;
    rom[42862] = 25'b1111110001100010010110010;
    rom[42863] = 25'b1111110001100011001111101;
    rom[42864] = 25'b1111110001100100001001000;
    rom[42865] = 25'b1111110001100101000010011;
    rom[42866] = 25'b1111110001100101111011111;
    rom[42867] = 25'b1111110001100110110101100;
    rom[42868] = 25'b1111110001100111101111001;
    rom[42869] = 25'b1111110001101000101000110;
    rom[42870] = 25'b1111110001101001100010011;
    rom[42871] = 25'b1111110001101010011100001;
    rom[42872] = 25'b1111110001101011010101111;
    rom[42873] = 25'b1111110001101100001111111;
    rom[42874] = 25'b1111110001101101001001110;
    rom[42875] = 25'b1111110001101110000011110;
    rom[42876] = 25'b1111110001101110111101110;
    rom[42877] = 25'b1111110001101111110111110;
    rom[42878] = 25'b1111110001110000110001111;
    rom[42879] = 25'b1111110001110001101100001;
    rom[42880] = 25'b1111110001110010100110011;
    rom[42881] = 25'b1111110001110011100000101;
    rom[42882] = 25'b1111110001110100011011000;
    rom[42883] = 25'b1111110001110101010101011;
    rom[42884] = 25'b1111110001110110001111111;
    rom[42885] = 25'b1111110001110111001010010;
    rom[42886] = 25'b1111110001111000000100111;
    rom[42887] = 25'b1111110001111000111111100;
    rom[42888] = 25'b1111110001111001111010001;
    rom[42889] = 25'b1111110001111010110100111;
    rom[42890] = 25'b1111110001111011101111101;
    rom[42891] = 25'b1111110001111100101010011;
    rom[42892] = 25'b1111110001111101100101010;
    rom[42893] = 25'b1111110001111110100000010;
    rom[42894] = 25'b1111110001111111011011001;
    rom[42895] = 25'b1111110010000000010110001;
    rom[42896] = 25'b1111110010000001010001010;
    rom[42897] = 25'b1111110010000010001100011;
    rom[42898] = 25'b1111110010000011000111100;
    rom[42899] = 25'b1111110010000100000010110;
    rom[42900] = 25'b1111110010000100111110000;
    rom[42901] = 25'b1111110010000101111001011;
    rom[42902] = 25'b1111110010000110110100110;
    rom[42903] = 25'b1111110010000111110000001;
    rom[42904] = 25'b1111110010001000101011101;
    rom[42905] = 25'b1111110010001001100111001;
    rom[42906] = 25'b1111110010001010100010110;
    rom[42907] = 25'b1111110010001011011110011;
    rom[42908] = 25'b1111110010001100011010001;
    rom[42909] = 25'b1111110010001101010101110;
    rom[42910] = 25'b1111110010001110010001101;
    rom[42911] = 25'b1111110010001111001101011;
    rom[42912] = 25'b1111110010010000001001010;
    rom[42913] = 25'b1111110010010001000101010;
    rom[42914] = 25'b1111110010010010000001001;
    rom[42915] = 25'b1111110010010010111101010;
    rom[42916] = 25'b1111110010010011111001011;
    rom[42917] = 25'b1111110010010100110101011;
    rom[42918] = 25'b1111110010010101110001101;
    rom[42919] = 25'b1111110010010110101101111;
    rom[42920] = 25'b1111110010010111101010001;
    rom[42921] = 25'b1111110010011000100110011;
    rom[42922] = 25'b1111110010011001100010111;
    rom[42923] = 25'b1111110010011010011111010;
    rom[42924] = 25'b1111110010011011011011110;
    rom[42925] = 25'b1111110010011100011000010;
    rom[42926] = 25'b1111110010011101010100110;
    rom[42927] = 25'b1111110010011110010001011;
    rom[42928] = 25'b1111110010011111001110000;
    rom[42929] = 25'b1111110010100000001010110;
    rom[42930] = 25'b1111110010100001000111100;
    rom[42931] = 25'b1111110010100010000100011;
    rom[42932] = 25'b1111110010100011000001010;
    rom[42933] = 25'b1111110010100011111110001;
    rom[42934] = 25'b1111110010100100111011001;
    rom[42935] = 25'b1111110010100101111000000;
    rom[42936] = 25'b1111110010100110110101000;
    rom[42937] = 25'b1111110010100111110010010;
    rom[42938] = 25'b1111110010101000101111010;
    rom[42939] = 25'b1111110010101001101100100;
    rom[42940] = 25'b1111110010101010101001110;
    rom[42941] = 25'b1111110010101011100111000;
    rom[42942] = 25'b1111110010101100100100011;
    rom[42943] = 25'b1111110010101101100001101;
    rom[42944] = 25'b1111110010101110011111001;
    rom[42945] = 25'b1111110010101111011100101;
    rom[42946] = 25'b1111110010110000011010001;
    rom[42947] = 25'b1111110010110001010111101;
    rom[42948] = 25'b1111110010110010010101010;
    rom[42949] = 25'b1111110010110011010010111;
    rom[42950] = 25'b1111110010110100010000101;
    rom[42951] = 25'b1111110010110101001110010;
    rom[42952] = 25'b1111110010110110001100001;
    rom[42953] = 25'b1111110010110111001010000;
    rom[42954] = 25'b1111110010111000000111111;
    rom[42955] = 25'b1111110010111001000101110;
    rom[42956] = 25'b1111110010111010000011110;
    rom[42957] = 25'b1111110010111011000001110;
    rom[42958] = 25'b1111110010111011111111110;
    rom[42959] = 25'b1111110010111100111101111;
    rom[42960] = 25'b1111110010111101111100000;
    rom[42961] = 25'b1111110010111110111010010;
    rom[42962] = 25'b1111110010111111111000100;
    rom[42963] = 25'b1111110011000000110110110;
    rom[42964] = 25'b1111110011000001110101001;
    rom[42965] = 25'b1111110011000010110011100;
    rom[42966] = 25'b1111110011000011110001111;
    rom[42967] = 25'b1111110011000100110000011;
    rom[42968] = 25'b1111110011000101101110110;
    rom[42969] = 25'b1111110011000110101101011;
    rom[42970] = 25'b1111110011000111101011111;
    rom[42971] = 25'b1111110011001000101010101;
    rom[42972] = 25'b1111110011001001101001010;
    rom[42973] = 25'b1111110011001010100111111;
    rom[42974] = 25'b1111110011001011100110101;
    rom[42975] = 25'b1111110011001100100101100;
    rom[42976] = 25'b1111110011001101100100011;
    rom[42977] = 25'b1111110011001110100011010;
    rom[42978] = 25'b1111110011001111100010001;
    rom[42979] = 25'b1111110011010000100001010;
    rom[42980] = 25'b1111110011010001100000001;
    rom[42981] = 25'b1111110011010010011111010;
    rom[42982] = 25'b1111110011010011011110010;
    rom[42983] = 25'b1111110011010100011101100;
    rom[42984] = 25'b1111110011010101011100101;
    rom[42985] = 25'b1111110011010110011011111;
    rom[42986] = 25'b1111110011010111011011010;
    rom[42987] = 25'b1111110011011000011010100;
    rom[42988] = 25'b1111110011011001011001111;
    rom[42989] = 25'b1111110011011010011001010;
    rom[42990] = 25'b1111110011011011011000101;
    rom[42991] = 25'b1111110011011100011000001;
    rom[42992] = 25'b1111110011011101010111101;
    rom[42993] = 25'b1111110011011110010111010;
    rom[42994] = 25'b1111110011011111010110111;
    rom[42995] = 25'b1111110011100000010110100;
    rom[42996] = 25'b1111110011100001010110001;
    rom[42997] = 25'b1111110011100010010101111;
    rom[42998] = 25'b1111110011100011010101110;
    rom[42999] = 25'b1111110011100100010101100;
    rom[43000] = 25'b1111110011100101010101011;
    rom[43001] = 25'b1111110011100110010101010;
    rom[43002] = 25'b1111110011100111010101001;
    rom[43003] = 25'b1111110011101000010101001;
    rom[43004] = 25'b1111110011101001010101001;
    rom[43005] = 25'b1111110011101010010101010;
    rom[43006] = 25'b1111110011101011010101010;
    rom[43007] = 25'b1111110011101100010101100;
    rom[43008] = 25'b1111110011101101010101101;
    rom[43009] = 25'b1111110011101110010101110;
    rom[43010] = 25'b1111110011101111010110000;
    rom[43011] = 25'b1111110011110000010110011;
    rom[43012] = 25'b1111110011110001010110101;
    rom[43013] = 25'b1111110011110010010111000;
    rom[43014] = 25'b1111110011110011010111011;
    rom[43015] = 25'b1111110011110100010111111;
    rom[43016] = 25'b1111110011110101011000011;
    rom[43017] = 25'b1111110011110110011000111;
    rom[43018] = 25'b1111110011110111011001011;
    rom[43019] = 25'b1111110011111000011010000;
    rom[43020] = 25'b1111110011111001011010101;
    rom[43021] = 25'b1111110011111010011011011;
    rom[43022] = 25'b1111110011111011011100000;
    rom[43023] = 25'b1111110011111100011100110;
    rom[43024] = 25'b1111110011111101011101101;
    rom[43025] = 25'b1111110011111110011110011;
    rom[43026] = 25'b1111110011111111011111010;
    rom[43027] = 25'b1111110100000000100000001;
    rom[43028] = 25'b1111110100000001100001001;
    rom[43029] = 25'b1111110100000010100010000;
    rom[43030] = 25'b1111110100000011100011001;
    rom[43031] = 25'b1111110100000100100100001;
    rom[43032] = 25'b1111110100000101100101010;
    rom[43033] = 25'b1111110100000110100110011;
    rom[43034] = 25'b1111110100000111100111100;
    rom[43035] = 25'b1111110100001000101000101;
    rom[43036] = 25'b1111110100001001101010000;
    rom[43037] = 25'b1111110100001010101011010;
    rom[43038] = 25'b1111110100001011101100100;
    rom[43039] = 25'b1111110100001100101101111;
    rom[43040] = 25'b1111110100001101101111010;
    rom[43041] = 25'b1111110100001110110000110;
    rom[43042] = 25'b1111110100001111110010001;
    rom[43043] = 25'b1111110100010000110011101;
    rom[43044] = 25'b1111110100010001110101001;
    rom[43045] = 25'b1111110100010010110110101;
    rom[43046] = 25'b1111110100010011111000011;
    rom[43047] = 25'b1111110100010100111010000;
    rom[43048] = 25'b1111110100010101111011101;
    rom[43049] = 25'b1111110100010110111101010;
    rom[43050] = 25'b1111110100010111111111000;
    rom[43051] = 25'b1111110100011001000000111;
    rom[43052] = 25'b1111110100011010000010101;
    rom[43053] = 25'b1111110100011011000100011;
    rom[43054] = 25'b1111110100011100000110011;
    rom[43055] = 25'b1111110100011101001000010;
    rom[43056] = 25'b1111110100011110001010010;
    rom[43057] = 25'b1111110100011111001100001;
    rom[43058] = 25'b1111110100100000001110001;
    rom[43059] = 25'b1111110100100001010000010;
    rom[43060] = 25'b1111110100100010010010011;
    rom[43061] = 25'b1111110100100011010100100;
    rom[43062] = 25'b1111110100100100010110101;
    rom[43063] = 25'b1111110100100101011000110;
    rom[43064] = 25'b1111110100100110011011000;
    rom[43065] = 25'b1111110100100111011101010;
    rom[43066] = 25'b1111110100101000011111100;
    rom[43067] = 25'b1111110100101001100001111;
    rom[43068] = 25'b1111110100101010100100010;
    rom[43069] = 25'b1111110100101011100110101;
    rom[43070] = 25'b1111110100101100101001000;
    rom[43071] = 25'b1111110100101101101011100;
    rom[43072] = 25'b1111110100101110101110000;
    rom[43073] = 25'b1111110100101111110000100;
    rom[43074] = 25'b1111110100110000110011001;
    rom[43075] = 25'b1111110100110001110101101;
    rom[43076] = 25'b1111110100110010111000010;
    rom[43077] = 25'b1111110100110011111010111;
    rom[43078] = 25'b1111110100110100111101101;
    rom[43079] = 25'b1111110100110110000000010;
    rom[43080] = 25'b1111110100110111000011000;
    rom[43081] = 25'b1111110100111000000101110;
    rom[43082] = 25'b1111110100111001001000101;
    rom[43083] = 25'b1111110100111010001011100;
    rom[43084] = 25'b1111110100111011001110011;
    rom[43085] = 25'b1111110100111100010001001;
    rom[43086] = 25'b1111110100111101010100001;
    rom[43087] = 25'b1111110100111110010111001;
    rom[43088] = 25'b1111110100111111011010000;
    rom[43089] = 25'b1111110101000000011101001;
    rom[43090] = 25'b1111110101000001100000001;
    rom[43091] = 25'b1111110101000010100011010;
    rom[43092] = 25'b1111110101000011100110011;
    rom[43093] = 25'b1111110101000100101001100;
    rom[43094] = 25'b1111110101000101101100110;
    rom[43095] = 25'b1111110101000110110000000;
    rom[43096] = 25'b1111110101000111110011010;
    rom[43097] = 25'b1111110101001000110110100;
    rom[43098] = 25'b1111110101001001111001110;
    rom[43099] = 25'b1111110101001010111101001;
    rom[43100] = 25'b1111110101001100000000100;
    rom[43101] = 25'b1111110101001101000011110;
    rom[43102] = 25'b1111110101001110000111010;
    rom[43103] = 25'b1111110101001111001010110;
    rom[43104] = 25'b1111110101010000001110001;
    rom[43105] = 25'b1111110101010001010001101;
    rom[43106] = 25'b1111110101010010010101010;
    rom[43107] = 25'b1111110101010011011000110;
    rom[43108] = 25'b1111110101010100011100011;
    rom[43109] = 25'b1111110101010101100000000;
    rom[43110] = 25'b1111110101010110100011101;
    rom[43111] = 25'b1111110101010111100111011;
    rom[43112] = 25'b1111110101011000101011000;
    rom[43113] = 25'b1111110101011001101110110;
    rom[43114] = 25'b1111110101011010110010100;
    rom[43115] = 25'b1111110101011011110110011;
    rom[43116] = 25'b1111110101011100111010001;
    rom[43117] = 25'b1111110101011101111110000;
    rom[43118] = 25'b1111110101011111000010000;
    rom[43119] = 25'b1111110101100000000101111;
    rom[43120] = 25'b1111110101100001001001110;
    rom[43121] = 25'b1111110101100010001101110;
    rom[43122] = 25'b1111110101100011010001110;
    rom[43123] = 25'b1111110101100100010101110;
    rom[43124] = 25'b1111110101100101011001110;
    rom[43125] = 25'b1111110101100110011101111;
    rom[43126] = 25'b1111110101100111100001111;
    rom[43127] = 25'b1111110101101000100110001;
    rom[43128] = 25'b1111110101101001101010010;
    rom[43129] = 25'b1111110101101010101110011;
    rom[43130] = 25'b1111110101101011110010101;
    rom[43131] = 25'b1111110101101100110110111;
    rom[43132] = 25'b1111110101101101111011001;
    rom[43133] = 25'b1111110101101110111111011;
    rom[43134] = 25'b1111110101110000000011110;
    rom[43135] = 25'b1111110101110001001000000;
    rom[43136] = 25'b1111110101110010001100011;
    rom[43137] = 25'b1111110101110011010000111;
    rom[43138] = 25'b1111110101110100010101010;
    rom[43139] = 25'b1111110101110101011001101;
    rom[43140] = 25'b1111110101110110011110001;
    rom[43141] = 25'b1111110101110111100010101;
    rom[43142] = 25'b1111110101111000100111010;
    rom[43143] = 25'b1111110101111001101011110;
    rom[43144] = 25'b1111110101111010110000010;
    rom[43145] = 25'b1111110101111011110100111;
    rom[43146] = 25'b1111110101111100111001100;
    rom[43147] = 25'b1111110101111101111110001;
    rom[43148] = 25'b1111110101111111000010110;
    rom[43149] = 25'b1111110110000000000111100;
    rom[43150] = 25'b1111110110000001001100010;
    rom[43151] = 25'b1111110110000010010001000;
    rom[43152] = 25'b1111110110000011010101101;
    rom[43153] = 25'b1111110110000100011010100;
    rom[43154] = 25'b1111110110000101011111011;
    rom[43155] = 25'b1111110110000110100100001;
    rom[43156] = 25'b1111110110000111101001000;
    rom[43157] = 25'b1111110110001000101101111;
    rom[43158] = 25'b1111110110001001110010111;
    rom[43159] = 25'b1111110110001010110111110;
    rom[43160] = 25'b1111110110001011111100110;
    rom[43161] = 25'b1111110110001101000001101;
    rom[43162] = 25'b1111110110001110000110110;
    rom[43163] = 25'b1111110110001111001011110;
    rom[43164] = 25'b1111110110010000010000111;
    rom[43165] = 25'b1111110110010001010101111;
    rom[43166] = 25'b1111110110010010011010111;
    rom[43167] = 25'b1111110110010011100000000;
    rom[43168] = 25'b1111110110010100100101010;
    rom[43169] = 25'b1111110110010101101010011;
    rom[43170] = 25'b1111110110010110101111100;
    rom[43171] = 25'b1111110110010111110100110;
    rom[43172] = 25'b1111110110011000111010000;
    rom[43173] = 25'b1111110110011001111111010;
    rom[43174] = 25'b1111110110011011000100100;
    rom[43175] = 25'b1111110110011100001001111;
    rom[43176] = 25'b1111110110011101001111010;
    rom[43177] = 25'b1111110110011110010100100;
    rom[43178] = 25'b1111110110011111011001111;
    rom[43179] = 25'b1111110110100000011111010;
    rom[43180] = 25'b1111110110100001100100101;
    rom[43181] = 25'b1111110110100010101010000;
    rom[43182] = 25'b1111110110100011101111100;
    rom[43183] = 25'b1111110110100100110101000;
    rom[43184] = 25'b1111110110100101111010100;
    rom[43185] = 25'b1111110110100111000000000;
    rom[43186] = 25'b1111110110101000000101100;
    rom[43187] = 25'b1111110110101001001011001;
    rom[43188] = 25'b1111110110101010010000110;
    rom[43189] = 25'b1111110110101011010110010;
    rom[43190] = 25'b1111110110101100011011111;
    rom[43191] = 25'b1111110110101101100001100;
    rom[43192] = 25'b1111110110101110100111001;
    rom[43193] = 25'b1111110110101111101100111;
    rom[43194] = 25'b1111110110110000110010100;
    rom[43195] = 25'b1111110110110001111000010;
    rom[43196] = 25'b1111110110110010111110000;
    rom[43197] = 25'b1111110110110100000011110;
    rom[43198] = 25'b1111110110110101001001100;
    rom[43199] = 25'b1111110110110110001111010;
    rom[43200] = 25'b1111110110110111010101001;
    rom[43201] = 25'b1111110110111000011010111;
    rom[43202] = 25'b1111110110111001100000110;
    rom[43203] = 25'b1111110110111010100110110;
    rom[43204] = 25'b1111110110111011101100101;
    rom[43205] = 25'b1111110110111100110010100;
    rom[43206] = 25'b1111110110111101111000011;
    rom[43207] = 25'b1111110110111110111110011;
    rom[43208] = 25'b1111110111000000000100010;
    rom[43209] = 25'b1111110111000001001010010;
    rom[43210] = 25'b1111110111000010010000010;
    rom[43211] = 25'b1111110111000011010110010;
    rom[43212] = 25'b1111110111000100011100011;
    rom[43213] = 25'b1111110111000101100010011;
    rom[43214] = 25'b1111110111000110101000100;
    rom[43215] = 25'b1111110111000111101110100;
    rom[43216] = 25'b1111110111001000110100101;
    rom[43217] = 25'b1111110111001001111010111;
    rom[43218] = 25'b1111110111001011000001000;
    rom[43219] = 25'b1111110111001100000111001;
    rom[43220] = 25'b1111110111001101001101010;
    rom[43221] = 25'b1111110111001110010011100;
    rom[43222] = 25'b1111110111001111011001101;
    rom[43223] = 25'b1111110111010000011111111;
    rom[43224] = 25'b1111110111010001100110001;
    rom[43225] = 25'b1111110111010010101100011;
    rom[43226] = 25'b1111110111010011110010101;
    rom[43227] = 25'b1111110111010100111001000;
    rom[43228] = 25'b1111110111010101111111011;
    rom[43229] = 25'b1111110111010111000101101;
    rom[43230] = 25'b1111110111011000001100000;
    rom[43231] = 25'b1111110111011001010010010;
    rom[43232] = 25'b1111110111011010011000110;
    rom[43233] = 25'b1111110111011011011111001;
    rom[43234] = 25'b1111110111011100100101100;
    rom[43235] = 25'b1111110111011101101011111;
    rom[43236] = 25'b1111110111011110110010011;
    rom[43237] = 25'b1111110111011111111000110;
    rom[43238] = 25'b1111110111100000111111010;
    rom[43239] = 25'b1111110111100010000101110;
    rom[43240] = 25'b1111110111100011001100010;
    rom[43241] = 25'b1111110111100100010010110;
    rom[43242] = 25'b1111110111100101011001010;
    rom[43243] = 25'b1111110111100110011111110;
    rom[43244] = 25'b1111110111100111100110011;
    rom[43245] = 25'b1111110111101000101100111;
    rom[43246] = 25'b1111110111101001110011100;
    rom[43247] = 25'b1111110111101010111010001;
    rom[43248] = 25'b1111110111101100000000110;
    rom[43249] = 25'b1111110111101101000111011;
    rom[43250] = 25'b1111110111101110001110000;
    rom[43251] = 25'b1111110111101111010100110;
    rom[43252] = 25'b1111110111110000011011011;
    rom[43253] = 25'b1111110111110001100010001;
    rom[43254] = 25'b1111110111110010101000110;
    rom[43255] = 25'b1111110111110011101111100;
    rom[43256] = 25'b1111110111110100110110001;
    rom[43257] = 25'b1111110111110101111101000;
    rom[43258] = 25'b1111110111110111000011101;
    rom[43259] = 25'b1111110111111000001010100;
    rom[43260] = 25'b1111110111111001010001010;
    rom[43261] = 25'b1111110111111010011000000;
    rom[43262] = 25'b1111110111111011011110110;
    rom[43263] = 25'b1111110111111100100101101;
    rom[43264] = 25'b1111110111111101101100100;
    rom[43265] = 25'b1111110111111110110011011;
    rom[43266] = 25'b1111110111111111111010001;
    rom[43267] = 25'b1111111000000001000001000;
    rom[43268] = 25'b1111111000000010000111111;
    rom[43269] = 25'b1111111000000011001110110;
    rom[43270] = 25'b1111111000000100010101101;
    rom[43271] = 25'b1111111000000101011100101;
    rom[43272] = 25'b1111111000000110100011100;
    rom[43273] = 25'b1111111000000111101010100;
    rom[43274] = 25'b1111111000001000110001100;
    rom[43275] = 25'b1111111000001001111000011;
    rom[43276] = 25'b1111111000001010111111011;
    rom[43277] = 25'b1111111000001100000110011;
    rom[43278] = 25'b1111111000001101001101011;
    rom[43279] = 25'b1111111000001110010100011;
    rom[43280] = 25'b1111111000001111011011011;
    rom[43281] = 25'b1111111000010000100010011;
    rom[43282] = 25'b1111111000010001101001100;
    rom[43283] = 25'b1111111000010010110000100;
    rom[43284] = 25'b1111111000010011110111101;
    rom[43285] = 25'b1111111000010100111110101;
    rom[43286] = 25'b1111111000010110000101110;
    rom[43287] = 25'b1111111000010111001100110;
    rom[43288] = 25'b1111111000011000010100000;
    rom[43289] = 25'b1111111000011001011011000;
    rom[43290] = 25'b1111111000011010100010001;
    rom[43291] = 25'b1111111000011011101001010;
    rom[43292] = 25'b1111111000011100110000011;
    rom[43293] = 25'b1111111000011101110111100;
    rom[43294] = 25'b1111111000011110111110110;
    rom[43295] = 25'b1111111000100000000101111;
    rom[43296] = 25'b1111111000100001001101000;
    rom[43297] = 25'b1111111000100010010100010;
    rom[43298] = 25'b1111111000100011011011100;
    rom[43299] = 25'b1111111000100100100010110;
    rom[43300] = 25'b1111111000100101101001111;
    rom[43301] = 25'b1111111000100110110001001;
    rom[43302] = 25'b1111111000100111111000011;
    rom[43303] = 25'b1111111000101000111111100;
    rom[43304] = 25'b1111111000101010000110110;
    rom[43305] = 25'b1111111000101011001110001;
    rom[43306] = 25'b1111111000101100010101011;
    rom[43307] = 25'b1111111000101101011100101;
    rom[43308] = 25'b1111111000101110100011111;
    rom[43309] = 25'b1111111000101111101011010;
    rom[43310] = 25'b1111111000110000110010100;
    rom[43311] = 25'b1111111000110001111001111;
    rom[43312] = 25'b1111111000110011000001001;
    rom[43313] = 25'b1111111000110100001000100;
    rom[43314] = 25'b1111111000110101001111110;
    rom[43315] = 25'b1111111000110110010111001;
    rom[43316] = 25'b1111111000110111011110100;
    rom[43317] = 25'b1111111000111000100101111;
    rom[43318] = 25'b1111111000111001101101010;
    rom[43319] = 25'b1111111000111010110100100;
    rom[43320] = 25'b1111111000111011111011111;
    rom[43321] = 25'b1111111000111101000011011;
    rom[43322] = 25'b1111111000111110001010101;
    rom[43323] = 25'b1111111000111111010010001;
    rom[43324] = 25'b1111111001000000011001100;
    rom[43325] = 25'b1111111001000001100000111;
    rom[43326] = 25'b1111111001000010101000011;
    rom[43327] = 25'b1111111001000011101111110;
    rom[43328] = 25'b1111111001000100110111001;
    rom[43329] = 25'b1111111001000101111110101;
    rom[43330] = 25'b1111111001000111000110000;
    rom[43331] = 25'b1111111001001000001101100;
    rom[43332] = 25'b1111111001001001010100111;
    rom[43333] = 25'b1111111001001010011100011;
    rom[43334] = 25'b1111111001001011100011110;
    rom[43335] = 25'b1111111001001100101011011;
    rom[43336] = 25'b1111111001001101110010110;
    rom[43337] = 25'b1111111001001110111010010;
    rom[43338] = 25'b1111111001010000000001110;
    rom[43339] = 25'b1111111001010001001001001;
    rom[43340] = 25'b1111111001010010010000110;
    rom[43341] = 25'b1111111001010011011000001;
    rom[43342] = 25'b1111111001010100011111110;
    rom[43343] = 25'b1111111001010101100111010;
    rom[43344] = 25'b1111111001010110101110101;
    rom[43345] = 25'b1111111001010111110110010;
    rom[43346] = 25'b1111111001011000111101110;
    rom[43347] = 25'b1111111001011010000101010;
    rom[43348] = 25'b1111111001011011001100110;
    rom[43349] = 25'b1111111001011100010100011;
    rom[43350] = 25'b1111111001011101011011111;
    rom[43351] = 25'b1111111001011110100011011;
    rom[43352] = 25'b1111111001011111101011000;
    rom[43353] = 25'b1111111001100000110010100;
    rom[43354] = 25'b1111111001100001111010000;
    rom[43355] = 25'b1111111001100011000001100;
    rom[43356] = 25'b1111111001100100001001001;
    rom[43357] = 25'b1111111001100101010000110;
    rom[43358] = 25'b1111111001100110011000010;
    rom[43359] = 25'b1111111001100111011111110;
    rom[43360] = 25'b1111111001101000100111011;
    rom[43361] = 25'b1111111001101001101110111;
    rom[43362] = 25'b1111111001101010110110100;
    rom[43363] = 25'b1111111001101011111110001;
    rom[43364] = 25'b1111111001101101000101101;
    rom[43365] = 25'b1111111001101110001101010;
    rom[43366] = 25'b1111111001101111010100110;
    rom[43367] = 25'b1111111001110000011100011;
    rom[43368] = 25'b1111111001110001100100000;
    rom[43369] = 25'b1111111001110010101011101;
    rom[43370] = 25'b1111111001110011110011010;
    rom[43371] = 25'b1111111001110100111010110;
    rom[43372] = 25'b1111111001110110000010011;
    rom[43373] = 25'b1111111001110111001001111;
    rom[43374] = 25'b1111111001111000010001100;
    rom[43375] = 25'b1111111001111001011001001;
    rom[43376] = 25'b1111111001111010100000110;
    rom[43377] = 25'b1111111001111011101000011;
    rom[43378] = 25'b1111111001111100110000000;
    rom[43379] = 25'b1111111001111101110111101;
    rom[43380] = 25'b1111111001111110111111001;
    rom[43381] = 25'b1111111010000000000110110;
    rom[43382] = 25'b1111111010000001001110011;
    rom[43383] = 25'b1111111010000010010110000;
    rom[43384] = 25'b1111111010000011011101100;
    rom[43385] = 25'b1111111010000100100101001;
    rom[43386] = 25'b1111111010000101101100110;
    rom[43387] = 25'b1111111010000110110100011;
    rom[43388] = 25'b1111111010000111111100000;
    rom[43389] = 25'b1111111010001001000011101;
    rom[43390] = 25'b1111111010001010001011010;
    rom[43391] = 25'b1111111010001011010010111;
    rom[43392] = 25'b1111111010001100011010100;
    rom[43393] = 25'b1111111010001101100010000;
    rom[43394] = 25'b1111111010001110101001101;
    rom[43395] = 25'b1111111010001111110001010;
    rom[43396] = 25'b1111111010010000111000111;
    rom[43397] = 25'b1111111010010010000000011;
    rom[43398] = 25'b1111111010010011001000000;
    rom[43399] = 25'b1111111010010100001111101;
    rom[43400] = 25'b1111111010010101010111010;
    rom[43401] = 25'b1111111010010110011110111;
    rom[43402] = 25'b1111111010010111100110100;
    rom[43403] = 25'b1111111010011000101110001;
    rom[43404] = 25'b1111111010011001110101101;
    rom[43405] = 25'b1111111010011010111101010;
    rom[43406] = 25'b1111111010011100000100110;
    rom[43407] = 25'b1111111010011101001100011;
    rom[43408] = 25'b1111111010011110010100000;
    rom[43409] = 25'b1111111010011111011011101;
    rom[43410] = 25'b1111111010100000100011010;
    rom[43411] = 25'b1111111010100001101010110;
    rom[43412] = 25'b1111111010100010110010011;
    rom[43413] = 25'b1111111010100011111001111;
    rom[43414] = 25'b1111111010100101000001100;
    rom[43415] = 25'b1111111010100110001001001;
    rom[43416] = 25'b1111111010100111010000101;
    rom[43417] = 25'b1111111010101000011000010;
    rom[43418] = 25'b1111111010101001011111110;
    rom[43419] = 25'b1111111010101010100111010;
    rom[43420] = 25'b1111111010101011101110111;
    rom[43421] = 25'b1111111010101100110110100;
    rom[43422] = 25'b1111111010101101111110000;
    rom[43423] = 25'b1111111010101111000101100;
    rom[43424] = 25'b1111111010110000001101001;
    rom[43425] = 25'b1111111010110001010100101;
    rom[43426] = 25'b1111111010110010011100001;
    rom[43427] = 25'b1111111010110011100011101;
    rom[43428] = 25'b1111111010110100101011010;
    rom[43429] = 25'b1111111010110101110010110;
    rom[43430] = 25'b1111111010110110111010010;
    rom[43431] = 25'b1111111010111000000001110;
    rom[43432] = 25'b1111111010111001001001011;
    rom[43433] = 25'b1111111010111010010000110;
    rom[43434] = 25'b1111111010111011011000011;
    rom[43435] = 25'b1111111010111100011111111;
    rom[43436] = 25'b1111111010111101100111010;
    rom[43437] = 25'b1111111010111110101110111;
    rom[43438] = 25'b1111111010111111110110010;
    rom[43439] = 25'b1111111011000000111101110;
    rom[43440] = 25'b1111111011000010000101010;
    rom[43441] = 25'b1111111011000011001100101;
    rom[43442] = 25'b1111111011000100010100010;
    rom[43443] = 25'b1111111011000101011011101;
    rom[43444] = 25'b1111111011000110100011001;
    rom[43445] = 25'b1111111011000111101010100;
    rom[43446] = 25'b1111111011001000110010000;
    rom[43447] = 25'b1111111011001001111001011;
    rom[43448] = 25'b1111111011001011000000111;
    rom[43449] = 25'b1111111011001100001000010;
    rom[43450] = 25'b1111111011001101001111110;
    rom[43451] = 25'b1111111011001110010111001;
    rom[43452] = 25'b1111111011001111011110100;
    rom[43453] = 25'b1111111011010000100110000;
    rom[43454] = 25'b1111111011010001101101011;
    rom[43455] = 25'b1111111011010010110100110;
    rom[43456] = 25'b1111111011010011111100001;
    rom[43457] = 25'b1111111011010101000011100;
    rom[43458] = 25'b1111111011010110001010111;
    rom[43459] = 25'b1111111011010111010010010;
    rom[43460] = 25'b1111111011011000011001101;
    rom[43461] = 25'b1111111011011001100001000;
    rom[43462] = 25'b1111111011011010101000010;
    rom[43463] = 25'b1111111011011011101111101;
    rom[43464] = 25'b1111111011011100110111000;
    rom[43465] = 25'b1111111011011101111110010;
    rom[43466] = 25'b1111111011011111000101101;
    rom[43467] = 25'b1111111011100000001100111;
    rom[43468] = 25'b1111111011100001010100010;
    rom[43469] = 25'b1111111011100010011011100;
    rom[43470] = 25'b1111111011100011100010110;
    rom[43471] = 25'b1111111011100100101010000;
    rom[43472] = 25'b1111111011100101110001010;
    rom[43473] = 25'b1111111011100110111000100;
    rom[43474] = 25'b1111111011100111111111110;
    rom[43475] = 25'b1111111011101001000111001;
    rom[43476] = 25'b1111111011101010001110011;
    rom[43477] = 25'b1111111011101011010101101;
    rom[43478] = 25'b1111111011101100011100110;
    rom[43479] = 25'b1111111011101101100100000;
    rom[43480] = 25'b1111111011101110101011001;
    rom[43481] = 25'b1111111011101111110010010;
    rom[43482] = 25'b1111111011110000111001101;
    rom[43483] = 25'b1111111011110010000000110;
    rom[43484] = 25'b1111111011110011000111111;
    rom[43485] = 25'b1111111011110100001111000;
    rom[43486] = 25'b1111111011110101010110010;
    rom[43487] = 25'b1111111011110110011101010;
    rom[43488] = 25'b1111111011110111100100011;
    rom[43489] = 25'b1111111011111000101011100;
    rom[43490] = 25'b1111111011111001110010101;
    rom[43491] = 25'b1111111011111010111001110;
    rom[43492] = 25'b1111111011111100000000110;
    rom[43493] = 25'b1111111011111101000111111;
    rom[43494] = 25'b1111111011111110001110111;
    rom[43495] = 25'b1111111011111111010110000;
    rom[43496] = 25'b1111111100000000011101001;
    rom[43497] = 25'b1111111100000001100100001;
    rom[43498] = 25'b1111111100000010101011001;
    rom[43499] = 25'b1111111100000011110010001;
    rom[43500] = 25'b1111111100000100111001001;
    rom[43501] = 25'b1111111100000110000000001;
    rom[43502] = 25'b1111111100000111000111001;
    rom[43503] = 25'b1111111100001000001110001;
    rom[43504] = 25'b1111111100001001010101000;
    rom[43505] = 25'b1111111100001010011100000;
    rom[43506] = 25'b1111111100001011100011000;
    rom[43507] = 25'b1111111100001100101001111;
    rom[43508] = 25'b1111111100001101110000111;
    rom[43509] = 25'b1111111100001110110111110;
    rom[43510] = 25'b1111111100001111111110101;
    rom[43511] = 25'b1111111100010001000101100;
    rom[43512] = 25'b1111111100010010001100011;
    rom[43513] = 25'b1111111100010011010011010;
    rom[43514] = 25'b1111111100010100011010000;
    rom[43515] = 25'b1111111100010101100000111;
    rom[43516] = 25'b1111111100010110100111110;
    rom[43517] = 25'b1111111100010111101110100;
    rom[43518] = 25'b1111111100011000110101010;
    rom[43519] = 25'b1111111100011001111100001;
    rom[43520] = 25'b1111111100011011000010111;
    rom[43521] = 25'b1111111100011100001001101;
    rom[43522] = 25'b1111111100011101010000011;
    rom[43523] = 25'b1111111100011110010111001;
    rom[43524] = 25'b1111111100011111011101111;
    rom[43525] = 25'b1111111100100000100100100;
    rom[43526] = 25'b1111111100100001101011010;
    rom[43527] = 25'b1111111100100010110001111;
    rom[43528] = 25'b1111111100100011111000101;
    rom[43529] = 25'b1111111100100100111111010;
    rom[43530] = 25'b1111111100100110000101111;
    rom[43531] = 25'b1111111100100111001100100;
    rom[43532] = 25'b1111111100101000010011001;
    rom[43533] = 25'b1111111100101001011001110;
    rom[43534] = 25'b1111111100101010100000010;
    rom[43535] = 25'b1111111100101011100110111;
    rom[43536] = 25'b1111111100101100101101100;
    rom[43537] = 25'b1111111100101101110100000;
    rom[43538] = 25'b1111111100101110111010100;
    rom[43539] = 25'b1111111100110000000001000;
    rom[43540] = 25'b1111111100110001000111100;
    rom[43541] = 25'b1111111100110010001110000;
    rom[43542] = 25'b1111111100110011010100100;
    rom[43543] = 25'b1111111100110100011011000;
    rom[43544] = 25'b1111111100110101100001100;
    rom[43545] = 25'b1111111100110110100111111;
    rom[43546] = 25'b1111111100110111101110010;
    rom[43547] = 25'b1111111100111000110100110;
    rom[43548] = 25'b1111111100111001111011000;
    rom[43549] = 25'b1111111100111011000001011;
    rom[43550] = 25'b1111111100111100000111110;
    rom[43551] = 25'b1111111100111101001110001;
    rom[43552] = 25'b1111111100111110010100011;
    rom[43553] = 25'b1111111100111111011010110;
    rom[43554] = 25'b1111111101000000100001000;
    rom[43555] = 25'b1111111101000001100111011;
    rom[43556] = 25'b1111111101000010101101101;
    rom[43557] = 25'b1111111101000011110011111;
    rom[43558] = 25'b1111111101000100111010000;
    rom[43559] = 25'b1111111101000110000000010;
    rom[43560] = 25'b1111111101000111000110100;
    rom[43561] = 25'b1111111101001000001100101;
    rom[43562] = 25'b1111111101001001010010111;
    rom[43563] = 25'b1111111101001010011001000;
    rom[43564] = 25'b1111111101001011011111001;
    rom[43565] = 25'b1111111101001100100101001;
    rom[43566] = 25'b1111111101001101101011010;
    rom[43567] = 25'b1111111101001110110001011;
    rom[43568] = 25'b1111111101001111110111100;
    rom[43569] = 25'b1111111101010000111101100;
    rom[43570] = 25'b1111111101010010000011100;
    rom[43571] = 25'b1111111101010011001001101;
    rom[43572] = 25'b1111111101010100001111100;
    rom[43573] = 25'b1111111101010101010101100;
    rom[43574] = 25'b1111111101010110011011100;
    rom[43575] = 25'b1111111101010111100001100;
    rom[43576] = 25'b1111111101011000100111011;
    rom[43577] = 25'b1111111101011001101101010;
    rom[43578] = 25'b1111111101011010110011001;
    rom[43579] = 25'b1111111101011011111001001;
    rom[43580] = 25'b1111111101011100111110111;
    rom[43581] = 25'b1111111101011110000100101;
    rom[43582] = 25'b1111111101011111001010100;
    rom[43583] = 25'b1111111101100000010000011;
    rom[43584] = 25'b1111111101100001010110001;
    rom[43585] = 25'b1111111101100010011011111;
    rom[43586] = 25'b1111111101100011100001101;
    rom[43587] = 25'b1111111101100100100111011;
    rom[43588] = 25'b1111111101100101101101001;
    rom[43589] = 25'b1111111101100110110010110;
    rom[43590] = 25'b1111111101100111111000011;
    rom[43591] = 25'b1111111101101000111110001;
    rom[43592] = 25'b1111111101101010000011110;
    rom[43593] = 25'b1111111101101011001001011;
    rom[43594] = 25'b1111111101101100001110111;
    rom[43595] = 25'b1111111101101101010100100;
    rom[43596] = 25'b1111111101101110011010000;
    rom[43597] = 25'b1111111101101111011111101;
    rom[43598] = 25'b1111111101110000100101001;
    rom[43599] = 25'b1111111101110001101010110;
    rom[43600] = 25'b1111111101110010110000001;
    rom[43601] = 25'b1111111101110011110101100;
    rom[43602] = 25'b1111111101110100111011000;
    rom[43603] = 25'b1111111101110110000000011;
    rom[43604] = 25'b1111111101110111000101110;
    rom[43605] = 25'b1111111101111000001011010;
    rom[43606] = 25'b1111111101111001010000101;
    rom[43607] = 25'b1111111101111010010110000;
    rom[43608] = 25'b1111111101111011011011010;
    rom[43609] = 25'b1111111101111100100000100;
    rom[43610] = 25'b1111111101111101100101111;
    rom[43611] = 25'b1111111101111110101011000;
    rom[43612] = 25'b1111111101111111110000011;
    rom[43613] = 25'b1111111110000000110101100;
    rom[43614] = 25'b1111111110000001111010110;
    rom[43615] = 25'b1111111110000011000000000;
    rom[43616] = 25'b1111111110000100000101000;
    rom[43617] = 25'b1111111110000101001010010;
    rom[43618] = 25'b1111111110000110001111011;
    rom[43619] = 25'b1111111110000111010100011;
    rom[43620] = 25'b1111111110001000011001100;
    rom[43621] = 25'b1111111110001001011110100;
    rom[43622] = 25'b1111111110001010100011101;
    rom[43623] = 25'b1111111110001011101000100;
    rom[43624] = 25'b1111111110001100101101100;
    rom[43625] = 25'b1111111110001101110010100;
    rom[43626] = 25'b1111111110001110110111100;
    rom[43627] = 25'b1111111110001111111100011;
    rom[43628] = 25'b1111111110010001000001010;
    rom[43629] = 25'b1111111110010010000110001;
    rom[43630] = 25'b1111111110010011001011000;
    rom[43631] = 25'b1111111110010100001111110;
    rom[43632] = 25'b1111111110010101010100101;
    rom[43633] = 25'b1111111110010110011001011;
    rom[43634] = 25'b1111111110010111011110001;
    rom[43635] = 25'b1111111110011000100010111;
    rom[43636] = 25'b1111111110011001100111101;
    rom[43637] = 25'b1111111110011010101100010;
    rom[43638] = 25'b1111111110011011110001000;
    rom[43639] = 25'b1111111110011100110101101;
    rom[43640] = 25'b1111111110011101111010010;
    rom[43641] = 25'b1111111110011110111110111;
    rom[43642] = 25'b1111111110100000000011100;
    rom[43643] = 25'b1111111110100001001000000;
    rom[43644] = 25'b1111111110100010001100100;
    rom[43645] = 25'b1111111110100011010001000;
    rom[43646] = 25'b1111111110100100010101100;
    rom[43647] = 25'b1111111110100101011010000;
    rom[43648] = 25'b1111111110100110011110011;
    rom[43649] = 25'b1111111110100111100010111;
    rom[43650] = 25'b1111111110101000100111001;
    rom[43651] = 25'b1111111110101001101011100;
    rom[43652] = 25'b1111111110101010101111111;
    rom[43653] = 25'b1111111110101011110100010;
    rom[43654] = 25'b1111111110101100111000100;
    rom[43655] = 25'b1111111110101101111100110;
    rom[43656] = 25'b1111111110101111000001000;
    rom[43657] = 25'b1111111110110000000101010;
    rom[43658] = 25'b1111111110110001001001011;
    rom[43659] = 25'b1111111110110010001101101;
    rom[43660] = 25'b1111111110110011010001110;
    rom[43661] = 25'b1111111110110100010101111;
    rom[43662] = 25'b1111111110110101011010000;
    rom[43663] = 25'b1111111110110110011110001;
    rom[43664] = 25'b1111111110110111100010000;
    rom[43665] = 25'b1111111110111000100110001;
    rom[43666] = 25'b1111111110111001101010001;
    rom[43667] = 25'b1111111110111010101110001;
    rom[43668] = 25'b1111111110111011110010000;
    rom[43669] = 25'b1111111110111100110101111;
    rom[43670] = 25'b1111111110111101111001110;
    rom[43671] = 25'b1111111110111110111101101;
    rom[43672] = 25'b1111111111000000000001101;
    rom[43673] = 25'b1111111111000001000101011;
    rom[43674] = 25'b1111111111000010001001001;
    rom[43675] = 25'b1111111111000011001100111;
    rom[43676] = 25'b1111111111000100010000101;
    rom[43677] = 25'b1111111111000101010100011;
    rom[43678] = 25'b1111111111000110011000001;
    rom[43679] = 25'b1111111111000111011011110;
    rom[43680] = 25'b1111111111001000011111010;
    rom[43681] = 25'b1111111111001001100010111;
    rom[43682] = 25'b1111111111001010100110100;
    rom[43683] = 25'b1111111111001011101010000;
    rom[43684] = 25'b1111111111001100101101101;
    rom[43685] = 25'b1111111111001101110001001;
    rom[43686] = 25'b1111111111001110110100101;
    rom[43687] = 25'b1111111111001111111000000;
    rom[43688] = 25'b1111111111010000111011100;
    rom[43689] = 25'b1111111111010001111110111;
    rom[43690] = 25'b1111111111010011000010010;
    rom[43691] = 25'b1111111111010100000101100;
    rom[43692] = 25'b1111111111010101001000111;
    rom[43693] = 25'b1111111111010110001100001;
    rom[43694] = 25'b1111111111010111001111011;
    rom[43695] = 25'b1111111111011000010010101;
    rom[43696] = 25'b1111111111011001010101111;
    rom[43697] = 25'b1111111111011010011001000;
    rom[43698] = 25'b1111111111011011011100001;
    rom[43699] = 25'b1111111111011100011111010;
    rom[43700] = 25'b1111111111011101100010011;
    rom[43701] = 25'b1111111111011110100101011;
    rom[43702] = 25'b1111111111011111101000011;
    rom[43703] = 25'b1111111111100000101011100;
    rom[43704] = 25'b1111111111100001101110011;
    rom[43705] = 25'b1111111111100010110001011;
    rom[43706] = 25'b1111111111100011110100010;
    rom[43707] = 25'b1111111111100100110111010;
    rom[43708] = 25'b1111111111100101111010001;
    rom[43709] = 25'b1111111111100110111100111;
    rom[43710] = 25'b1111111111100111111111110;
    rom[43711] = 25'b1111111111101001000010100;
    rom[43712] = 25'b1111111111101010000101010;
    rom[43713] = 25'b1111111111101011001000000;
    rom[43714] = 25'b1111111111101100001010101;
    rom[43715] = 25'b1111111111101101001101010;
    rom[43716] = 25'b1111111111101110001111111;
    rom[43717] = 25'b1111111111101111010010101;
    rom[43718] = 25'b1111111111110000010101000;
    rom[43719] = 25'b1111111111110001010111101;
    rom[43720] = 25'b1111111111110010011010001;
    rom[43721] = 25'b1111111111110011011100101;
    rom[43722] = 25'b1111111111110100011111001;
    rom[43723] = 25'b1111111111110101100001100;
    rom[43724] = 25'b1111111111110110100011111;
    rom[43725] = 25'b1111111111110111100110010;
    rom[43726] = 25'b1111111111111000101000101;
    rom[43727] = 25'b1111111111111001101010111;
    rom[43728] = 25'b1111111111111010101101010;
    rom[43729] = 25'b1111111111111011101111011;
    rom[43730] = 25'b1111111111111100110001101;
    rom[43731] = 25'b1111111111111101110011111;
    rom[43732] = 25'b1111111111111110110110000;
    rom[43733] = 25'b1111111111111111111000001;
    rom[43734] = 25'b0000000000000000111010001;
    rom[43735] = 25'b0000000000000001111100001;
    rom[43736] = 25'b0000000000000010111110001;
    rom[43737] = 25'b0000000000000100000000010;
    rom[43738] = 25'b0000000000000101000010001;
    rom[43739] = 25'b0000000000000110000100000;
    rom[43740] = 25'b0000000000000111000110000;
    rom[43741] = 25'b0000000000001000000111111;
    rom[43742] = 25'b0000000000001001001001110;
    rom[43743] = 25'b0000000000001010001011100;
    rom[43744] = 25'b0000000000001011001101011;
    rom[43745] = 25'b0000000000001100001111001;
    rom[43746] = 25'b0000000000001101010000110;
    rom[43747] = 25'b0000000000001110010010100;
    rom[43748] = 25'b0000000000001111010100001;
    rom[43749] = 25'b0000000000010000010101110;
    rom[43750] = 25'b0000000000010001010111011;
    rom[43751] = 25'b0000000000010010011000111;
    rom[43752] = 25'b0000000000010011011010100;
    rom[43753] = 25'b0000000000010100011011111;
    rom[43754] = 25'b0000000000010101011101011;
    rom[43755] = 25'b0000000000010110011110111;
    rom[43756] = 25'b0000000000010111100000010;
    rom[43757] = 25'b0000000000011000100001101;
    rom[43758] = 25'b0000000000011001100010111;
    rom[43759] = 25'b0000000000011010100100010;
    rom[43760] = 25'b0000000000011011100101100;
    rom[43761] = 25'b0000000000011100100110110;
    rom[43762] = 25'b0000000000011101100111111;
    rom[43763] = 25'b0000000000011110101001001;
    rom[43764] = 25'b0000000000011111101010010;
    rom[43765] = 25'b0000000000100000101011011;
    rom[43766] = 25'b0000000000100001101100011;
    rom[43767] = 25'b0000000000100010101101011;
    rom[43768] = 25'b0000000000100011101110011;
    rom[43769] = 25'b0000000000100100101111011;
    rom[43770] = 25'b0000000000100101110000011;
    rom[43771] = 25'b0000000000100110110001010;
    rom[43772] = 25'b0000000000100111110010001;
    rom[43773] = 25'b0000000000101000110011000;
    rom[43774] = 25'b0000000000101001110011110;
    rom[43775] = 25'b0000000000101010110100101;
    rom[43776] = 25'b0000000000101011110101010;
    rom[43777] = 25'b0000000000101100110110000;
    rom[43778] = 25'b0000000000101101110110101;
    rom[43779] = 25'b0000000000101110110111010;
    rom[43780] = 25'b0000000000101111110111111;
    rom[43781] = 25'b0000000000110000111000011;
    rom[43782] = 25'b0000000000110001111000111;
    rom[43783] = 25'b0000000000110010111001100;
    rom[43784] = 25'b0000000000110011111001111;
    rom[43785] = 25'b0000000000110100111010011;
    rom[43786] = 25'b0000000000110101111010110;
    rom[43787] = 25'b0000000000110110111011001;
    rom[43788] = 25'b0000000000110111111011100;
    rom[43789] = 25'b0000000000111000111011110;
    rom[43790] = 25'b0000000000111001111100000;
    rom[43791] = 25'b0000000000111010111100010;
    rom[43792] = 25'b0000000000111011111100011;
    rom[43793] = 25'b0000000000111100111100100;
    rom[43794] = 25'b0000000000111101111100101;
    rom[43795] = 25'b0000000000111110111100110;
    rom[43796] = 25'b0000000000111111111100110;
    rom[43797] = 25'b0000000001000000111100110;
    rom[43798] = 25'b0000000001000001111100110;
    rom[43799] = 25'b0000000001000010111100110;
    rom[43800] = 25'b0000000001000011111100101;
    rom[43801] = 25'b0000000001000100111100100;
    rom[43802] = 25'b0000000001000101111100011;
    rom[43803] = 25'b0000000001000110111100001;
    rom[43804] = 25'b0000000001000111111011111;
    rom[43805] = 25'b0000000001001000111011101;
    rom[43806] = 25'b0000000001001001111011010;
    rom[43807] = 25'b0000000001001010111010111;
    rom[43808] = 25'b0000000001001011111010101;
    rom[43809] = 25'b0000000001001100111010001;
    rom[43810] = 25'b0000000001001101111001101;
    rom[43811] = 25'b0000000001001110111001001;
    rom[43812] = 25'b0000000001001111111000110;
    rom[43813] = 25'b0000000001010000111000001;
    rom[43814] = 25'b0000000001010001110111100;
    rom[43815] = 25'b0000000001010010110110111;
    rom[43816] = 25'b0000000001010011110110001;
    rom[43817] = 25'b0000000001010100110101100;
    rom[43818] = 25'b0000000001010101110100101;
    rom[43819] = 25'b0000000001010110110011111;
    rom[43820] = 25'b0000000001010111110011001;
    rom[43821] = 25'b0000000001011000110010010;
    rom[43822] = 25'b0000000001011001110001010;
    rom[43823] = 25'b0000000001011010110000011;
    rom[43824] = 25'b0000000001011011101111100;
    rom[43825] = 25'b0000000001011100101110011;
    rom[43826] = 25'b0000000001011101101101011;
    rom[43827] = 25'b0000000001011110101100010;
    rom[43828] = 25'b0000000001011111101011001;
    rom[43829] = 25'b0000000001100000101010000;
    rom[43830] = 25'b0000000001100001101000111;
    rom[43831] = 25'b0000000001100010100111101;
    rom[43832] = 25'b0000000001100011100110011;
    rom[43833] = 25'b0000000001100100100101000;
    rom[43834] = 25'b0000000001100101100011101;
    rom[43835] = 25'b0000000001100110100010010;
    rom[43836] = 25'b0000000001100111100000111;
    rom[43837] = 25'b0000000001101000011111011;
    rom[43838] = 25'b0000000001101001011101111;
    rom[43839] = 25'b0000000001101010011100011;
    rom[43840] = 25'b0000000001101011011010110;
    rom[43841] = 25'b0000000001101100011001010;
    rom[43842] = 25'b0000000001101101010111100;
    rom[43843] = 25'b0000000001101110010101110;
    rom[43844] = 25'b0000000001101111010100000;
    rom[43845] = 25'b0000000001110000010010011;
    rom[43846] = 25'b0000000001110001010000100;
    rom[43847] = 25'b0000000001110010001110101;
    rom[43848] = 25'b0000000001110011001100110;
    rom[43849] = 25'b0000000001110100001010111;
    rom[43850] = 25'b0000000001110101001000111;
    rom[43851] = 25'b0000000001110110000110111;
    rom[43852] = 25'b0000000001110111000100110;
    rom[43853] = 25'b0000000001111000000010110;
    rom[43854] = 25'b0000000001111001000000101;
    rom[43855] = 25'b0000000001111001111110100;
    rom[43856] = 25'b0000000001111010111100010;
    rom[43857] = 25'b0000000001111011111010000;
    rom[43858] = 25'b0000000001111100110111110;
    rom[43859] = 25'b0000000001111101110101100;
    rom[43860] = 25'b0000000001111110110011001;
    rom[43861] = 25'b0000000001111111110000101;
    rom[43862] = 25'b0000000010000000101110010;
    rom[43863] = 25'b0000000010000001101011110;
    rom[43864] = 25'b0000000010000010101001010;
    rom[43865] = 25'b0000000010000011100110110;
    rom[43866] = 25'b0000000010000100100100000;
    rom[43867] = 25'b0000000010000101100001011;
    rom[43868] = 25'b0000000010000110011110110;
    rom[43869] = 25'b0000000010000111011100000;
    rom[43870] = 25'b0000000010001000011001010;
    rom[43871] = 25'b0000000010001001010110100;
    rom[43872] = 25'b0000000010001010010011101;
    rom[43873] = 25'b0000000010001011010000110;
    rom[43874] = 25'b0000000010001100001101111;
    rom[43875] = 25'b0000000010001101001010111;
    rom[43876] = 25'b0000000010001110000111111;
    rom[43877] = 25'b0000000010001111000100111;
    rom[43878] = 25'b0000000010010000000001110;
    rom[43879] = 25'b0000000010010000111110101;
    rom[43880] = 25'b0000000010010001111011100;
    rom[43881] = 25'b0000000010010010111000010;
    rom[43882] = 25'b0000000010010011110101000;
    rom[43883] = 25'b0000000010010100110001101;
    rom[43884] = 25'b0000000010010101101110011;
    rom[43885] = 25'b0000000010010110101011000;
    rom[43886] = 25'b0000000010010111100111101;
    rom[43887] = 25'b0000000010011000100100001;
    rom[43888] = 25'b0000000010011001100000101;
    rom[43889] = 25'b0000000010011010011101001;
    rom[43890] = 25'b0000000010011011011001100;
    rom[43891] = 25'b0000000010011100010101111;
    rom[43892] = 25'b0000000010011101010010010;
    rom[43893] = 25'b0000000010011110001110100;
    rom[43894] = 25'b0000000010011111001010110;
    rom[43895] = 25'b0000000010100000000111000;
    rom[43896] = 25'b0000000010100001000011001;
    rom[43897] = 25'b0000000010100001111111010;
    rom[43898] = 25'b0000000010100010111011011;
    rom[43899] = 25'b0000000010100011110111011;
    rom[43900] = 25'b0000000010100100110011100;
    rom[43901] = 25'b0000000010100101101111011;
    rom[43902] = 25'b0000000010100110101011010;
    rom[43903] = 25'b0000000010100111100111010;
    rom[43904] = 25'b0000000010101000100011000;
    rom[43905] = 25'b0000000010101001011110110;
    rom[43906] = 25'b0000000010101010011010100;
    rom[43907] = 25'b0000000010101011010110010;
    rom[43908] = 25'b0000000010101100010001111;
    rom[43909] = 25'b0000000010101101001101100;
    rom[43910] = 25'b0000000010101110001001001;
    rom[43911] = 25'b0000000010101111000100101;
    rom[43912] = 25'b0000000010110000000000001;
    rom[43913] = 25'b0000000010110000111011101;
    rom[43914] = 25'b0000000010110001110111000;
    rom[43915] = 25'b0000000010110010110010010;
    rom[43916] = 25'b0000000010110011101101101;
    rom[43917] = 25'b0000000010110100101000111;
    rom[43918] = 25'b0000000010110101100100001;
    rom[43919] = 25'b0000000010110110011111010;
    rom[43920] = 25'b0000000010110111011010011;
    rom[43921] = 25'b0000000010111000010101100;
    rom[43922] = 25'b0000000010111001010000100;
    rom[43923] = 25'b0000000010111010001011100;
    rom[43924] = 25'b0000000010111011000110101;
    rom[43925] = 25'b0000000010111100000001100;
    rom[43926] = 25'b0000000010111100111100011;
    rom[43927] = 25'b0000000010111101110111001;
    rom[43928] = 25'b0000000010111110110010000;
    rom[43929] = 25'b0000000010111111101100110;
    rom[43930] = 25'b0000000011000000100111011;
    rom[43931] = 25'b0000000011000001100010000;
    rom[43932] = 25'b0000000011000010011100110;
    rom[43933] = 25'b0000000011000011010111010;
    rom[43934] = 25'b0000000011000100010001110;
    rom[43935] = 25'b0000000011000101001100010;
    rom[43936] = 25'b0000000011000110000110110;
    rom[43937] = 25'b0000000011000111000001001;
    rom[43938] = 25'b0000000011000111111011100;
    rom[43939] = 25'b0000000011001000110101110;
    rom[43940] = 25'b0000000011001001110000000;
    rom[43941] = 25'b0000000011001010101010001;
    rom[43942] = 25'b0000000011001011100100011;
    rom[43943] = 25'b0000000011001100011110100;
    rom[43944] = 25'b0000000011001101011000100;
    rom[43945] = 25'b0000000011001110010010101;
    rom[43946] = 25'b0000000011001111001100101;
    rom[43947] = 25'b0000000011010000000110100;
    rom[43948] = 25'b0000000011010001000000011;
    rom[43949] = 25'b0000000011010001111010011;
    rom[43950] = 25'b0000000011010010110100001;
    rom[43951] = 25'b0000000011010011101101111;
    rom[43952] = 25'b0000000011010100100111100;
    rom[43953] = 25'b0000000011010101100001010;
    rom[43954] = 25'b0000000011010110011010111;
    rom[43955] = 25'b0000000011010111010100011;
    rom[43956] = 25'b0000000011011000001101111;
    rom[43957] = 25'b0000000011011001000111100;
    rom[43958] = 25'b0000000011011010000000111;
    rom[43959] = 25'b0000000011011010111010011;
    rom[43960] = 25'b0000000011011011110011101;
    rom[43961] = 25'b0000000011011100101100111;
    rom[43962] = 25'b0000000011011101100110001;
    rom[43963] = 25'b0000000011011110011111011;
    rom[43964] = 25'b0000000011011111011000100;
    rom[43965] = 25'b0000000011100000010001110;
    rom[43966] = 25'b0000000011100001001010110;
    rom[43967] = 25'b0000000011100010000011111;
    rom[43968] = 25'b0000000011100010111100110;
    rom[43969] = 25'b0000000011100011110101101;
    rom[43970] = 25'b0000000011100100101110100;
    rom[43971] = 25'b0000000011100101100111011;
    rom[43972] = 25'b0000000011100110100000010;
    rom[43973] = 25'b0000000011100111011001000;
    rom[43974] = 25'b0000000011101000010001101;
    rom[43975] = 25'b0000000011101001001010011;
    rom[43976] = 25'b0000000011101010000010111;
    rom[43977] = 25'b0000000011101010111011011;
    rom[43978] = 25'b0000000011101011110100000;
    rom[43979] = 25'b0000000011101100101100011;
    rom[43980] = 25'b0000000011101101100100111;
    rom[43981] = 25'b0000000011101110011101010;
    rom[43982] = 25'b0000000011101111010101100;
    rom[43983] = 25'b0000000011110000001101111;
    rom[43984] = 25'b0000000011110001000110001;
    rom[43985] = 25'b0000000011110001111110010;
    rom[43986] = 25'b0000000011110010110110011;
    rom[43987] = 25'b0000000011110011101110100;
    rom[43988] = 25'b0000000011110100100110100;
    rom[43989] = 25'b0000000011110101011110100;
    rom[43990] = 25'b0000000011110110010110100;
    rom[43991] = 25'b0000000011110111001110011;
    rom[43992] = 25'b0000000011111000000110001;
    rom[43993] = 25'b0000000011111000111110000;
    rom[43994] = 25'b0000000011111001110101110;
    rom[43995] = 25'b0000000011111010101101011;
    rom[43996] = 25'b0000000011111011100101001;
    rom[43997] = 25'b0000000011111100011100110;
    rom[43998] = 25'b0000000011111101010100010;
    rom[43999] = 25'b0000000011111110001011110;
    rom[44000] = 25'b0000000011111111000011010;
    rom[44001] = 25'b0000000011111111111010101;
    rom[44002] = 25'b0000000100000000110010000;
    rom[44003] = 25'b0000000100000001101001011;
    rom[44004] = 25'b0000000100000010100000101;
    rom[44005] = 25'b0000000100000011010111111;
    rom[44006] = 25'b0000000100000100001111000;
    rom[44007] = 25'b0000000100000101000110001;
    rom[44008] = 25'b0000000100000101111101010;
    rom[44009] = 25'b0000000100000110110100010;
    rom[44010] = 25'b0000000100000111101011010;
    rom[44011] = 25'b0000000100001000100010001;
    rom[44012] = 25'b0000000100001001011001001;
    rom[44013] = 25'b0000000100001010001111111;
    rom[44014] = 25'b0000000100001011000110101;
    rom[44015] = 25'b0000000100001011111101011;
    rom[44016] = 25'b0000000100001100110100001;
    rom[44017] = 25'b0000000100001101101010110;
    rom[44018] = 25'b0000000100001110100001011;
    rom[44019] = 25'b0000000100001111010111111;
    rom[44020] = 25'b0000000100010000001110011;
    rom[44021] = 25'b0000000100010001000100110;
    rom[44022] = 25'b0000000100010001111011010;
    rom[44023] = 25'b0000000100010010110001100;
    rom[44024] = 25'b0000000100010011100111110;
    rom[44025] = 25'b0000000100010100011110001;
    rom[44026] = 25'b0000000100010101010100010;
    rom[44027] = 25'b0000000100010110001010011;
    rom[44028] = 25'b0000000100010111000000100;
    rom[44029] = 25'b0000000100010111110110100;
    rom[44030] = 25'b0000000100011000101100100;
    rom[44031] = 25'b0000000100011001100010011;
    rom[44032] = 25'b0000000100011010011000011;
    rom[44033] = 25'b0000000100011011001110001;
    rom[44034] = 25'b0000000100011100000100000;
    rom[44035] = 25'b0000000100011100111001110;
    rom[44036] = 25'b0000000100011101101111100;
    rom[44037] = 25'b0000000100011110100101000;
    rom[44038] = 25'b0000000100011111011010101;
    rom[44039] = 25'b0000000100100000010000001;
    rom[44040] = 25'b0000000100100001000101101;
    rom[44041] = 25'b0000000100100001111011001;
    rom[44042] = 25'b0000000100100010110000100;
    rom[44043] = 25'b0000000100100011100101111;
    rom[44044] = 25'b0000000100100100011011001;
    rom[44045] = 25'b0000000100100101010000011;
    rom[44046] = 25'b0000000100100110000101101;
    rom[44047] = 25'b0000000100100110111010110;
    rom[44048] = 25'b0000000100100111101111110;
    rom[44049] = 25'b0000000100101000100100111;
    rom[44050] = 25'b0000000100101001011001110;
    rom[44051] = 25'b0000000100101010001110110;
    rom[44052] = 25'b0000000100101011000011110;
    rom[44053] = 25'b0000000100101011111000100;
    rom[44054] = 25'b0000000100101100101101011;
    rom[44055] = 25'b0000000100101101100010000;
    rom[44056] = 25'b0000000100101110010110101;
    rom[44057] = 25'b0000000100101111001011011;
    rom[44058] = 25'b0000000100101111111111111;
    rom[44059] = 25'b0000000100110000110100011;
    rom[44060] = 25'b0000000100110001101000111;
    rom[44061] = 25'b0000000100110010011101011;
    rom[44062] = 25'b0000000100110011010001110;
    rom[44063] = 25'b0000000100110100000110000;
    rom[44064] = 25'b0000000100110100111010011;
    rom[44065] = 25'b0000000100110101101110100;
    rom[44066] = 25'b0000000100110110100010101;
    rom[44067] = 25'b0000000100110111010110110;
    rom[44068] = 25'b0000000100111000001010111;
    rom[44069] = 25'b0000000100111000111110111;
    rom[44070] = 25'b0000000100111001110010111;
    rom[44071] = 25'b0000000100111010100110110;
    rom[44072] = 25'b0000000100111011011010101;
    rom[44073] = 25'b0000000100111100001110011;
    rom[44074] = 25'b0000000100111101000010001;
    rom[44075] = 25'b0000000100111101110101111;
    rom[44076] = 25'b0000000100111110101001100;
    rom[44077] = 25'b0000000100111111011101001;
    rom[44078] = 25'b0000000101000000010000110;
    rom[44079] = 25'b0000000101000001000100001;
    rom[44080] = 25'b0000000101000001110111101;
    rom[44081] = 25'b0000000101000010101011000;
    rom[44082] = 25'b0000000101000011011110011;
    rom[44083] = 25'b0000000101000100010001101;
    rom[44084] = 25'b0000000101000101000100111;
    rom[44085] = 25'b0000000101000101111000000;
    rom[44086] = 25'b0000000101000110101011001;
    rom[44087] = 25'b0000000101000111011110010;
    rom[44088] = 25'b0000000101001000010001010;
    rom[44089] = 25'b0000000101001001000100010;
    rom[44090] = 25'b0000000101001001110111001;
    rom[44091] = 25'b0000000101001010101010000;
    rom[44092] = 25'b0000000101001011011100110;
    rom[44093] = 25'b0000000101001100001111101;
    rom[44094] = 25'b0000000101001101000010010;
    rom[44095] = 25'b0000000101001101110100111;
    rom[44096] = 25'b0000000101001110100111100;
    rom[44097] = 25'b0000000101001111011010001;
    rom[44098] = 25'b0000000101010000001100101;
    rom[44099] = 25'b0000000101010000111111000;
    rom[44100] = 25'b0000000101010001110001011;
    rom[44101] = 25'b0000000101010010100011101;
    rom[44102] = 25'b0000000101010011010110000;
    rom[44103] = 25'b0000000101010100001000001;
    rom[44104] = 25'b0000000101010100111010011;
    rom[44105] = 25'b0000000101010101101100100;
    rom[44106] = 25'b0000000101010110011110101;
    rom[44107] = 25'b0000000101010111010000101;
    rom[44108] = 25'b0000000101011000000010100;
    rom[44109] = 25'b0000000101011000110100011;
    rom[44110] = 25'b0000000101011001100110010;
    rom[44111] = 25'b0000000101011010011000001;
    rom[44112] = 25'b0000000101011011001001111;
    rom[44113] = 25'b0000000101011011111011100;
    rom[44114] = 25'b0000000101011100101101010;
    rom[44115] = 25'b0000000101011101011110110;
    rom[44116] = 25'b0000000101011110010000010;
    rom[44117] = 25'b0000000101011111000001110;
    rom[44118] = 25'b0000000101011111110011001;
    rom[44119] = 25'b0000000101100000100100101;
    rom[44120] = 25'b0000000101100001010101111;
    rom[44121] = 25'b0000000101100010000111001;
    rom[44122] = 25'b0000000101100010111000011;
    rom[44123] = 25'b0000000101100011101001100;
    rom[44124] = 25'b0000000101100100011010100;
    rom[44125] = 25'b0000000101100101001011101;
    rom[44126] = 25'b0000000101100101111100101;
    rom[44127] = 25'b0000000101100110101101100;
    rom[44128] = 25'b0000000101100111011110011;
    rom[44129] = 25'b0000000101101000001111010;
    rom[44130] = 25'b0000000101101001000000001;
    rom[44131] = 25'b0000000101101001110000110;
    rom[44132] = 25'b0000000101101010100001011;
    rom[44133] = 25'b0000000101101011010010000;
    rom[44134] = 25'b0000000101101100000010101;
    rom[44135] = 25'b0000000101101100110011001;
    rom[44136] = 25'b0000000101101101100011100;
    rom[44137] = 25'b0000000101101110010011111;
    rom[44138] = 25'b0000000101101111000100010;
    rom[44139] = 25'b0000000101101111110100100;
    rom[44140] = 25'b0000000101110000100100110;
    rom[44141] = 25'b0000000101110001010101000;
    rom[44142] = 25'b0000000101110010000101000;
    rom[44143] = 25'b0000000101110010110101001;
    rom[44144] = 25'b0000000101110011100101001;
    rom[44145] = 25'b0000000101110100010101000;
    rom[44146] = 25'b0000000101110101000101000;
    rom[44147] = 25'b0000000101110101110100110;
    rom[44148] = 25'b0000000101110110100100101;
    rom[44149] = 25'b0000000101110111010100010;
    rom[44150] = 25'b0000000101111000000011111;
    rom[44151] = 25'b0000000101111000110011100;
    rom[44152] = 25'b0000000101111001100011001;
    rom[44153] = 25'b0000000101111010010010101;
    rom[44154] = 25'b0000000101111011000010000;
    rom[44155] = 25'b0000000101111011110001100;
    rom[44156] = 25'b0000000101111100100000111;
    rom[44157] = 25'b0000000101111101010000001;
    rom[44158] = 25'b0000000101111101111111011;
    rom[44159] = 25'b0000000101111110101110100;
    rom[44160] = 25'b0000000101111111011101101;
    rom[44161] = 25'b0000000110000000001100110;
    rom[44162] = 25'b0000000110000000111011110;
    rom[44163] = 25'b0000000110000001101010101;
    rom[44164] = 25'b0000000110000010011001101;
    rom[44165] = 25'b0000000110000011001000011;
    rom[44166] = 25'b0000000110000011110111001;
    rom[44167] = 25'b0000000110000100100101111;
    rom[44168] = 25'b0000000110000101010100101;
    rom[44169] = 25'b0000000110000110000011010;
    rom[44170] = 25'b0000000110000110110001110;
    rom[44171] = 25'b0000000110000111100000010;
    rom[44172] = 25'b0000000110001000001110110;
    rom[44173] = 25'b0000000110001000111101000;
    rom[44174] = 25'b0000000110001001101011011;
    rom[44175] = 25'b0000000110001010011001110;
    rom[44176] = 25'b0000000110001011000111111;
    rom[44177] = 25'b0000000110001011110110000;
    rom[44178] = 25'b0000000110001100100100010;
    rom[44179] = 25'b0000000110001101010010010;
    rom[44180] = 25'b0000000110001110000000010;
    rom[44181] = 25'b0000000110001110101110010;
    rom[44182] = 25'b0000000110001111011100001;
    rom[44183] = 25'b0000000110010000001001111;
    rom[44184] = 25'b0000000110010000110111101;
    rom[44185] = 25'b0000000110010001100101011;
    rom[44186] = 25'b0000000110010010010011000;
    rom[44187] = 25'b0000000110010011000000101;
    rom[44188] = 25'b0000000110010011101110001;
    rom[44189] = 25'b0000000110010100011011101;
    rom[44190] = 25'b0000000110010101001001001;
    rom[44191] = 25'b0000000110010101110110100;
    rom[44192] = 25'b0000000110010110100011110;
    rom[44193] = 25'b0000000110010111010001000;
    rom[44194] = 25'b0000000110010111111110010;
    rom[44195] = 25'b0000000110011000101011011;
    rom[44196] = 25'b0000000110011001011000100;
    rom[44197] = 25'b0000000110011010000101100;
    rom[44198] = 25'b0000000110011010110010100;
    rom[44199] = 25'b0000000110011011011111100;
    rom[44200] = 25'b0000000110011100001100010;
    rom[44201] = 25'b0000000110011100111001001;
    rom[44202] = 25'b0000000110011101100101111;
    rom[44203] = 25'b0000000110011110010010100;
    rom[44204] = 25'b0000000110011110111111001;
    rom[44205] = 25'b0000000110011111101011101;
    rom[44206] = 25'b0000000110100000011000010;
    rom[44207] = 25'b0000000110100001000100101;
    rom[44208] = 25'b0000000110100001110001001;
    rom[44209] = 25'b0000000110100010011101100;
    rom[44210] = 25'b0000000110100011001001110;
    rom[44211] = 25'b0000000110100011110101111;
    rom[44212] = 25'b0000000110100100100010001;
    rom[44213] = 25'b0000000110100101001110010;
    rom[44214] = 25'b0000000110100101111010010;
    rom[44215] = 25'b0000000110100110100110010;
    rom[44216] = 25'b0000000110100111010010010;
    rom[44217] = 25'b0000000110100111111110001;
    rom[44218] = 25'b0000000110101000101001111;
    rom[44219] = 25'b0000000110101001010101110;
    rom[44220] = 25'b0000000110101010000001011;
    rom[44221] = 25'b0000000110101010101101000;
    rom[44222] = 25'b0000000110101011011000101;
    rom[44223] = 25'b0000000110101100000100001;
    rom[44224] = 25'b0000000110101100101111101;
    rom[44225] = 25'b0000000110101101011011001;
    rom[44226] = 25'b0000000110101110000110011;
    rom[44227] = 25'b0000000110101110110001110;
    rom[44228] = 25'b0000000110101111011101000;
    rom[44229] = 25'b0000000110110000001000001;
    rom[44230] = 25'b0000000110110000110011010;
    rom[44231] = 25'b0000000110110001011110011;
    rom[44232] = 25'b0000000110110010001001011;
    rom[44233] = 25'b0000000110110010110100011;
    rom[44234] = 25'b0000000110110011011111010;
    rom[44235] = 25'b0000000110110100001010001;
    rom[44236] = 25'b0000000110110100110100111;
    rom[44237] = 25'b0000000110110101011111100;
    rom[44238] = 25'b0000000110110110001010010;
    rom[44239] = 25'b0000000110110110110100110;
    rom[44240] = 25'b0000000110110111011111011;
    rom[44241] = 25'b0000000110111000001001111;
    rom[44242] = 25'b0000000110111000110100010;
    rom[44243] = 25'b0000000110111001011110101;
    rom[44244] = 25'b0000000110111010001001000;
    rom[44245] = 25'b0000000110111010110011001;
    rom[44246] = 25'b0000000110111011011101011;
    rom[44247] = 25'b0000000110111100000111100;
    rom[44248] = 25'b0000000110111100110001101;
    rom[44249] = 25'b0000000110111101011011101;
    rom[44250] = 25'b0000000110111110000101101;
    rom[44251] = 25'b0000000110111110101111100;
    rom[44252] = 25'b0000000110111111011001011;
    rom[44253] = 25'b0000000111000000000011001;
    rom[44254] = 25'b0000000111000000101100111;
    rom[44255] = 25'b0000000111000001010110100;
    rom[44256] = 25'b0000000111000010000000001;
    rom[44257] = 25'b0000000111000010101001101;
    rom[44258] = 25'b0000000111000011010011001;
    rom[44259] = 25'b0000000111000011111100100;
    rom[44260] = 25'b0000000111000100100101111;
    rom[44261] = 25'b0000000111000101001111010;
    rom[44262] = 25'b0000000111000101111000011;
    rom[44263] = 25'b0000000111000110100001101;
    rom[44264] = 25'b0000000111000111001010110;
    rom[44265] = 25'b0000000111000111110011111;
    rom[44266] = 25'b0000000111001000011100111;
    rom[44267] = 25'b0000000111001001000101110;
    rom[44268] = 25'b0000000111001001101110110;
    rom[44269] = 25'b0000000111001010010111101;
    rom[44270] = 25'b0000000111001011000000011;
    rom[44271] = 25'b0000000111001011101001000;
    rom[44272] = 25'b0000000111001100010001101;
    rom[44273] = 25'b0000000111001100111010010;
    rom[44274] = 25'b0000000111001101100010110;
    rom[44275] = 25'b0000000111001110001011011;
    rom[44276] = 25'b0000000111001110110011101;
    rom[44277] = 25'b0000000111001111011100001;
    rom[44278] = 25'b0000000111010000000100011;
    rom[44279] = 25'b0000000111010000101100101;
    rom[44280] = 25'b0000000111010001010100110;
    rom[44281] = 25'b0000000111010001111100111;
    rom[44282] = 25'b0000000111010010100101000;
    rom[44283] = 25'b0000000111010011001101000;
    rom[44284] = 25'b0000000111010011110100111;
    rom[44285] = 25'b0000000111010100011100111;
    rom[44286] = 25'b0000000111010101000100101;
    rom[44287] = 25'b0000000111010101101100011;
    rom[44288] = 25'b0000000111010110010100001;
    rom[44289] = 25'b0000000111010110111011110;
    rom[44290] = 25'b0000000111010111100011010;
    rom[44291] = 25'b0000000111011000001010111;
    rom[44292] = 25'b0000000111011000110010010;
    rom[44293] = 25'b0000000111011001011001101;
    rom[44294] = 25'b0000000111011010000001000;
    rom[44295] = 25'b0000000111011010101000010;
    rom[44296] = 25'b0000000111011011001111100;
    rom[44297] = 25'b0000000111011011110110101;
    rom[44298] = 25'b0000000111011100011101110;
    rom[44299] = 25'b0000000111011101000100111;
    rom[44300] = 25'b0000000111011101101011110;
    rom[44301] = 25'b0000000111011110010010110;
    rom[44302] = 25'b0000000111011110111001100;
    rom[44303] = 25'b0000000111011111100000011;
    rom[44304] = 25'b0000000111100000000111001;
    rom[44305] = 25'b0000000111100000101101111;
    rom[44306] = 25'b0000000111100001010100011;
    rom[44307] = 25'b0000000111100001111011000;
    rom[44308] = 25'b0000000111100010100001011;
    rom[44309] = 25'b0000000111100011000111111;
    rom[44310] = 25'b0000000111100011101110010;
    rom[44311] = 25'b0000000111100100010100101;
    rom[44312] = 25'b0000000111100100111010111;
    rom[44313] = 25'b0000000111100101100001001;
    rom[44314] = 25'b0000000111100110000111001;
    rom[44315] = 25'b0000000111100110101101010;
    rom[44316] = 25'b0000000111100111010011010;
    rom[44317] = 25'b0000000111100111111001010;
    rom[44318] = 25'b0000000111101000011111001;
    rom[44319] = 25'b0000000111101001000100111;
    rom[44320] = 25'b0000000111101001101010101;
    rom[44321] = 25'b0000000111101010010000011;
    rom[44322] = 25'b0000000111101010110110000;
    rom[44323] = 25'b0000000111101011011011101;
    rom[44324] = 25'b0000000111101100000001001;
    rom[44325] = 25'b0000000111101100100110101;
    rom[44326] = 25'b0000000111101101001100000;
    rom[44327] = 25'b0000000111101101110001011;
    rom[44328] = 25'b0000000111101110010110101;
    rom[44329] = 25'b0000000111101110111011111;
    rom[44330] = 25'b0000000111101111100001000;
    rom[44331] = 25'b0000000111110000000110001;
    rom[44332] = 25'b0000000111110000101011010;
    rom[44333] = 25'b0000000111110001010000001;
    rom[44334] = 25'b0000000111110001110101001;
    rom[44335] = 25'b0000000111110010011001111;
    rom[44336] = 25'b0000000111110010111110101;
    rom[44337] = 25'b0000000111110011100011100;
    rom[44338] = 25'b0000000111110100001000000;
    rom[44339] = 25'b0000000111110100101100110;
    rom[44340] = 25'b0000000111110101010001010;
    rom[44341] = 25'b0000000111110101110101110;
    rom[44342] = 25'b0000000111110110011010010;
    rom[44343] = 25'b0000000111110110111110100;
    rom[44344] = 25'b0000000111110111100010111;
    rom[44345] = 25'b0000000111111000000111001;
    rom[44346] = 25'b0000000111111000101011010;
    rom[44347] = 25'b0000000111111001001111011;
    rom[44348] = 25'b0000000111111001110011011;
    rom[44349] = 25'b0000000111111010010111100;
    rom[44350] = 25'b0000000111111010111011011;
    rom[44351] = 25'b0000000111111011011111010;
    rom[44352] = 25'b0000000111111100000011000;
    rom[44353] = 25'b0000000111111100100110111;
    rom[44354] = 25'b0000000111111101001010100;
    rom[44355] = 25'b0000000111111101101110001;
    rom[44356] = 25'b0000000111111110010001101;
    rom[44357] = 25'b0000000111111110110101010;
    rom[44358] = 25'b0000000111111111011000101;
    rom[44359] = 25'b0000000111111111111100000;
    rom[44360] = 25'b0000001000000000011111011;
    rom[44361] = 25'b0000001000000001000010101;
    rom[44362] = 25'b0000001000000001100101111;
    rom[44363] = 25'b0000001000000010001001000;
    rom[44364] = 25'b0000001000000010101100000;
    rom[44365] = 25'b0000001000000011001111000;
    rom[44366] = 25'b0000001000000011110010000;
    rom[44367] = 25'b0000001000000100010100111;
    rom[44368] = 25'b0000001000000100110111101;
    rom[44369] = 25'b0000001000000101011010100;
    rom[44370] = 25'b0000001000000101111101001;
    rom[44371] = 25'b0000001000000110011111110;
    rom[44372] = 25'b0000001000000111000010011;
    rom[44373] = 25'b0000001000000111100100111;
    rom[44374] = 25'b0000001000001000000111011;
    rom[44375] = 25'b0000001000001000101001110;
    rom[44376] = 25'b0000001000001001001100001;
    rom[44377] = 25'b0000001000001001101110011;
    rom[44378] = 25'b0000001000001010010000100;
    rom[44379] = 25'b0000001000001010110010110;
    rom[44380] = 25'b0000001000001011010100111;
    rom[44381] = 25'b0000001000001011110110110;
    rom[44382] = 25'b0000001000001100011000110;
    rom[44383] = 25'b0000001000001100111010110;
    rom[44384] = 25'b0000001000001101011100100;
    rom[44385] = 25'b0000001000001101111110011;
    rom[44386] = 25'b0000001000001110100000000;
    rom[44387] = 25'b0000001000001111000001101;
    rom[44388] = 25'b0000001000001111100011010;
    rom[44389] = 25'b0000001000010000000100110;
    rom[44390] = 25'b0000001000010000100110010;
    rom[44391] = 25'b0000001000010001000111101;
    rom[44392] = 25'b0000001000010001101001000;
    rom[44393] = 25'b0000001000010010001010010;
    rom[44394] = 25'b0000001000010010101011100;
    rom[44395] = 25'b0000001000010011001100101;
    rom[44396] = 25'b0000001000010011101101110;
    rom[44397] = 25'b0000001000010100001110101;
    rom[44398] = 25'b0000001000010100101111101;
    rom[44399] = 25'b0000001000010101010000101;
    rom[44400] = 25'b0000001000010101110001011;
    rom[44401] = 25'b0000001000010110010010001;
    rom[44402] = 25'b0000001000010110110010111;
    rom[44403] = 25'b0000001000010111010011100;
    rom[44404] = 25'b0000001000010111110100001;
    rom[44405] = 25'b0000001000011000010100110;
    rom[44406] = 25'b0000001000011000110101001;
    rom[44407] = 25'b0000001000011001010101100;
    rom[44408] = 25'b0000001000011001110101111;
    rom[44409] = 25'b0000001000011010010110001;
    rom[44410] = 25'b0000001000011010110110011;
    rom[44411] = 25'b0000001000011011010110101;
    rom[44412] = 25'b0000001000011011110110101;
    rom[44413] = 25'b0000001000011100010110101;
    rom[44414] = 25'b0000001000011100110110101;
    rom[44415] = 25'b0000001000011101010110100;
    rom[44416] = 25'b0000001000011101110110011;
    rom[44417] = 25'b0000001000011110010110001;
    rom[44418] = 25'b0000001000011110110101111;
    rom[44419] = 25'b0000001000011111010101100;
    rom[44420] = 25'b0000001000011111110101001;
    rom[44421] = 25'b0000001000100000010100101;
    rom[44422] = 25'b0000001000100000110100001;
    rom[44423] = 25'b0000001000100001010011100;
    rom[44424] = 25'b0000001000100001110010110;
    rom[44425] = 25'b0000001000100010010010001;
    rom[44426] = 25'b0000001000100010110001011;
    rom[44427] = 25'b0000001000100011010000100;
    rom[44428] = 25'b0000001000100011101111100;
    rom[44429] = 25'b0000001000100100001110100;
    rom[44430] = 25'b0000001000100100101101101;
    rom[44431] = 25'b0000001000100101001100100;
    rom[44432] = 25'b0000001000100101101011010;
    rom[44433] = 25'b0000001000100110001010000;
    rom[44434] = 25'b0000001000100110101000110;
    rom[44435] = 25'b0000001000100111000111011;
    rom[44436] = 25'b0000001000100111100110000;
    rom[44437] = 25'b0000001000101000000100100;
    rom[44438] = 25'b0000001000101000100011000;
    rom[44439] = 25'b0000001000101001000001011;
    rom[44440] = 25'b0000001000101001011111110;
    rom[44441] = 25'b0000001000101001111110000;
    rom[44442] = 25'b0000001000101010011100010;
    rom[44443] = 25'b0000001000101010111010011;
    rom[44444] = 25'b0000001000101011011000100;
    rom[44445] = 25'b0000001000101011110110011;
    rom[44446] = 25'b0000001000101100010100011;
    rom[44447] = 25'b0000001000101100110010010;
    rom[44448] = 25'b0000001000101101010000001;
    rom[44449] = 25'b0000001000101101101101111;
    rom[44450] = 25'b0000001000101110001011100;
    rom[44451] = 25'b0000001000101110101001010;
    rom[44452] = 25'b0000001000101111000110110;
    rom[44453] = 25'b0000001000101111100100010;
    rom[44454] = 25'b0000001000110000000001110;
    rom[44455] = 25'b0000001000110000011111010;
    rom[44456] = 25'b0000001000110000111100100;
    rom[44457] = 25'b0000001000110001011001110;
    rom[44458] = 25'b0000001000110001110111000;
    rom[44459] = 25'b0000001000110010010100001;
    rom[44460] = 25'b0000001000110010110001001;
    rom[44461] = 25'b0000001000110011001110001;
    rom[44462] = 25'b0000001000110011101011001;
    rom[44463] = 25'b0000001000110100001000000;
    rom[44464] = 25'b0000001000110100100100110;
    rom[44465] = 25'b0000001000110101000001100;
    rom[44466] = 25'b0000001000110101011110010;
    rom[44467] = 25'b0000001000110101111010111;
    rom[44468] = 25'b0000001000110110010111100;
    rom[44469] = 25'b0000001000110110110100000;
    rom[44470] = 25'b0000001000110111010000011;
    rom[44471] = 25'b0000001000110111101100110;
    rom[44472] = 25'b0000001000111000001001001;
    rom[44473] = 25'b0000001000111000100101010;
    rom[44474] = 25'b0000001000111001000001100;
    rom[44475] = 25'b0000001000111001011101101;
    rom[44476] = 25'b0000001000111001111001110;
    rom[44477] = 25'b0000001000111010010101110;
    rom[44478] = 25'b0000001000111010110001101;
    rom[44479] = 25'b0000001000111011001101100;
    rom[44480] = 25'b0000001000111011101001011;
    rom[44481] = 25'b0000001000111100000101001;
    rom[44482] = 25'b0000001000111100100000110;
    rom[44483] = 25'b0000001000111100111100011;
    rom[44484] = 25'b0000001000111101010111111;
    rom[44485] = 25'b0000001000111101110011011;
    rom[44486] = 25'b0000001000111110001110110;
    rom[44487] = 25'b0000001000111110101010001;
    rom[44488] = 25'b0000001000111111000101100;
    rom[44489] = 25'b0000001000111111100000110;
    rom[44490] = 25'b0000001000111111111011111;
    rom[44491] = 25'b0000001001000000010111000;
    rom[44492] = 25'b0000001001000000110010000;
    rom[44493] = 25'b0000001001000001001101000;
    rom[44494] = 25'b0000001001000001100111111;
    rom[44495] = 25'b0000001001000010000010111;
    rom[44496] = 25'b0000001001000010011101101;
    rom[44497] = 25'b0000001001000010111000011;
    rom[44498] = 25'b0000001001000011010011000;
    rom[44499] = 25'b0000001001000011101101101;
    rom[44500] = 25'b0000001001000100001000001;
    rom[44501] = 25'b0000001001000100100010101;
    rom[44502] = 25'b0000001001000100111101000;
    rom[44503] = 25'b0000001001000101010111011;
    rom[44504] = 25'b0000001001000101110001101;
    rom[44505] = 25'b0000001001000110001011111;
    rom[44506] = 25'b0000001001000110100110000;
    rom[44507] = 25'b0000001001000111000000001;
    rom[44508] = 25'b0000001001000111011010001;
    rom[44509] = 25'b0000001001000111110100001;
    rom[44510] = 25'b0000001001001000001110000;
    rom[44511] = 25'b0000001001001000100111111;
    rom[44512] = 25'b0000001001001001000001101;
    rom[44513] = 25'b0000001001001001011011011;
    rom[44514] = 25'b0000001001001001110101000;
    rom[44515] = 25'b0000001001001010001110100;
    rom[44516] = 25'b0000001001001010101000001;
    rom[44517] = 25'b0000001001001011000001100;
    rom[44518] = 25'b0000001001001011011010111;
    rom[44519] = 25'b0000001001001011110100010;
    rom[44520] = 25'b0000001001001100001101100;
    rom[44521] = 25'b0000001001001100100110110;
    rom[44522] = 25'b0000001001001100111111111;
    rom[44523] = 25'b0000001001001101011001000;
    rom[44524] = 25'b0000001001001101110010000;
    rom[44525] = 25'b0000001001001110001011000;
    rom[44526] = 25'b0000001001001110100011110;
    rom[44527] = 25'b0000001001001110111100101;
    rom[44528] = 25'b0000001001001111010101011;
    rom[44529] = 25'b0000001001001111101110000;
    rom[44530] = 25'b0000001001010000000110110;
    rom[44531] = 25'b0000001001010000011111010;
    rom[44532] = 25'b0000001001010000110111110;
    rom[44533] = 25'b0000001001010001010000010;
    rom[44534] = 25'b0000001001010001101000101;
    rom[44535] = 25'b0000001001010010000000111;
    rom[44536] = 25'b0000001001010010011001001;
    rom[44537] = 25'b0000001001010010110001011;
    rom[44538] = 25'b0000001001010011001001011;
    rom[44539] = 25'b0000001001010011100001100;
    rom[44540] = 25'b0000001001010011111001100;
    rom[44541] = 25'b0000001001010100010001011;
    rom[44542] = 25'b0000001001010100101001011;
    rom[44543] = 25'b0000001001010101000001001;
    rom[44544] = 25'b0000001001010101011000111;
    rom[44545] = 25'b0000001001010101110000100;
    rom[44546] = 25'b0000001001010110001000001;
    rom[44547] = 25'b0000001001010110011111101;
    rom[44548] = 25'b0000001001010110110111001;
    rom[44549] = 25'b0000001001010111001110100;
    rom[44550] = 25'b0000001001010111100101111;
    rom[44551] = 25'b0000001001010111111101010;
    rom[44552] = 25'b0000001001011000010100100;
    rom[44553] = 25'b0000001001011000101011101;
    rom[44554] = 25'b0000001001011001000010110;
    rom[44555] = 25'b0000001001011001011001110;
    rom[44556] = 25'b0000001001011001110000110;
    rom[44557] = 25'b0000001001011010000111101;
    rom[44558] = 25'b0000001001011010011110100;
    rom[44559] = 25'b0000001001011010110101010;
    rom[44560] = 25'b0000001001011011001100000;
    rom[44561] = 25'b0000001001011011100010101;
    rom[44562] = 25'b0000001001011011111001001;
    rom[44563] = 25'b0000001001011100001111110;
    rom[44564] = 25'b0000001001011100100110010;
    rom[44565] = 25'b0000001001011100111100101;
    rom[44566] = 25'b0000001001011101010010111;
    rom[44567] = 25'b0000001001011101101001010;
    rom[44568] = 25'b0000001001011101111111011;
    rom[44569] = 25'b0000001001011110010101100;
    rom[44570] = 25'b0000001001011110101011101;
    rom[44571] = 25'b0000001001011111000001101;
    rom[44572] = 25'b0000001001011111010111101;
    rom[44573] = 25'b0000001001011111101101100;
    rom[44574] = 25'b0000001001100000000011011;
    rom[44575] = 25'b0000001001100000011001001;
    rom[44576] = 25'b0000001001100000101110110;
    rom[44577] = 25'b0000001001100001000100011;
    rom[44578] = 25'b0000001001100001011010000;
    rom[44579] = 25'b0000001001100001101111100;
    rom[44580] = 25'b0000001001100010000101000;
    rom[44581] = 25'b0000001001100010011010011;
    rom[44582] = 25'b0000001001100010101111101;
    rom[44583] = 25'b0000001001100011000100111;
    rom[44584] = 25'b0000001001100011011010000;
    rom[44585] = 25'b0000001001100011101111001;
    rom[44586] = 25'b0000001001100100000100010;
    rom[44587] = 25'b0000001001100100011001010;
    rom[44588] = 25'b0000001001100100101110001;
    rom[44589] = 25'b0000001001100101000011000;
    rom[44590] = 25'b0000001001100101010111111;
    rom[44591] = 25'b0000001001100101101100100;
    rom[44592] = 25'b0000001001100110000001010;
    rom[44593] = 25'b0000001001100110010101111;
    rom[44594] = 25'b0000001001100110101010011;
    rom[44595] = 25'b0000001001100110111110111;
    rom[44596] = 25'b0000001001100111010011010;
    rom[44597] = 25'b0000001001100111100111101;
    rom[44598] = 25'b0000001001100111111100000;
    rom[44599] = 25'b0000001001101000010000001;
    rom[44600] = 25'b0000001001101000100100011;
    rom[44601] = 25'b0000001001101000111000011;
    rom[44602] = 25'b0000001001101001001100100;
    rom[44603] = 25'b0000001001101001100000100;
    rom[44604] = 25'b0000001001101001110100011;
    rom[44605] = 25'b0000001001101010001000010;
    rom[44606] = 25'b0000001001101010011100001;
    rom[44607] = 25'b0000001001101010101111110;
    rom[44608] = 25'b0000001001101011000011011;
    rom[44609] = 25'b0000001001101011010111000;
    rom[44610] = 25'b0000001001101011101010100;
    rom[44611] = 25'b0000001001101011111101111;
    rom[44612] = 25'b0000001001101100010001011;
    rom[44613] = 25'b0000001001101100100100110;
    rom[44614] = 25'b0000001001101100111000000;
    rom[44615] = 25'b0000001001101101001011001;
    rom[44616] = 25'b0000001001101101011110010;
    rom[44617] = 25'b0000001001101101110001100;
    rom[44618] = 25'b0000001001101110000100011;
    rom[44619] = 25'b0000001001101110010111011;
    rom[44620] = 25'b0000001001101110101010011;
    rom[44621] = 25'b0000001001101110111101001;
    rom[44622] = 25'b0000001001101111001111111;
    rom[44623] = 25'b0000001001101111100010100;
    rom[44624] = 25'b0000001001101111110101010;
    rom[44625] = 25'b0000001001110000000111110;
    rom[44626] = 25'b0000001001110000011010010;
    rom[44627] = 25'b0000001001110000101100110;
    rom[44628] = 25'b0000001001110000111111001;
    rom[44629] = 25'b0000001001110001010001100;
    rom[44630] = 25'b0000001001110001100011110;
    rom[44631] = 25'b0000001001110001110101111;
    rom[44632] = 25'b0000001001110010001000000;
    rom[44633] = 25'b0000001001110010011010000;
    rom[44634] = 25'b0000001001110010101100001;
    rom[44635] = 25'b0000001001110010111110000;
    rom[44636] = 25'b0000001001110011001111111;
    rom[44637] = 25'b0000001001110011100001101;
    rom[44638] = 25'b0000001001110011110011011;
    rom[44639] = 25'b0000001001110100000101001;
    rom[44640] = 25'b0000001001110100010110110;
    rom[44641] = 25'b0000001001110100101000010;
    rom[44642] = 25'b0000001001110100111001111;
    rom[44643] = 25'b0000001001110101001011010;
    rom[44644] = 25'b0000001001110101011100101;
    rom[44645] = 25'b0000001001110101101101111;
    rom[44646] = 25'b0000001001110101111111001;
    rom[44647] = 25'b0000001001110110010000010;
    rom[44648] = 25'b0000001001110110100001011;
    rom[44649] = 25'b0000001001110110110010100;
    rom[44650] = 25'b0000001001110111000011011;
    rom[44651] = 25'b0000001001110111010100011;
    rom[44652] = 25'b0000001001110111100101010;
    rom[44653] = 25'b0000001001110111110110000;
    rom[44654] = 25'b0000001001111000000110110;
    rom[44655] = 25'b0000001001111000010111011;
    rom[44656] = 25'b0000001001111000101000000;
    rom[44657] = 25'b0000001001111000111000100;
    rom[44658] = 25'b0000001001111001001001000;
    rom[44659] = 25'b0000001001111001011001011;
    rom[44660] = 25'b0000001001111001101001110;
    rom[44661] = 25'b0000001001111001111010000;
    rom[44662] = 25'b0000001001111010001010010;
    rom[44663] = 25'b0000001001111010011010011;
    rom[44664] = 25'b0000001001111010101010100;
    rom[44665] = 25'b0000001001111010111010100;
    rom[44666] = 25'b0000001001111011001010100;
    rom[44667] = 25'b0000001001111011011010011;
    rom[44668] = 25'b0000001001111011101010010;
    rom[44669] = 25'b0000001001111011111010000;
    rom[44670] = 25'b0000001001111100001001110;
    rom[44671] = 25'b0000001001111100011001011;
    rom[44672] = 25'b0000001001111100101001000;
    rom[44673] = 25'b0000001001111100111000100;
    rom[44674] = 25'b0000001001111101001000000;
    rom[44675] = 25'b0000001001111101010111011;
    rom[44676] = 25'b0000001001111101100110110;
    rom[44677] = 25'b0000001001111101110101111;
    rom[44678] = 25'b0000001001111110000101001;
    rom[44679] = 25'b0000001001111110010100010;
    rom[44680] = 25'b0000001001111110100011011;
    rom[44681] = 25'b0000001001111110110010011;
    rom[44682] = 25'b0000001001111111000001011;
    rom[44683] = 25'b0000001001111111010000010;
    rom[44684] = 25'b0000001001111111011111001;
    rom[44685] = 25'b0000001001111111101101111;
    rom[44686] = 25'b0000001001111111111100100;
    rom[44687] = 25'b0000001010000000001011001;
    rom[44688] = 25'b0000001010000000011001110;
    rom[44689] = 25'b0000001010000000101000010;
    rom[44690] = 25'b0000001010000000110110101;
    rom[44691] = 25'b0000001010000001000101000;
    rom[44692] = 25'b0000001010000001010011011;
    rom[44693] = 25'b0000001010000001100001101;
    rom[44694] = 25'b0000001010000001101111111;
    rom[44695] = 25'b0000001010000001111101111;
    rom[44696] = 25'b0000001010000010001100000;
    rom[44697] = 25'b0000001010000010011010000;
    rom[44698] = 25'b0000001010000010101000000;
    rom[44699] = 25'b0000001010000010110101111;
    rom[44700] = 25'b0000001010000011000011110;
    rom[44701] = 25'b0000001010000011010001011;
    rom[44702] = 25'b0000001010000011011111001;
    rom[44703] = 25'b0000001010000011101100101;
    rom[44704] = 25'b0000001010000011111010011;
    rom[44705] = 25'b0000001010000100000111110;
    rom[44706] = 25'b0000001010000100010101010;
    rom[44707] = 25'b0000001010000100100010101;
    rom[44708] = 25'b0000001010000100101111111;
    rom[44709] = 25'b0000001010000100111101001;
    rom[44710] = 25'b0000001010000101001010011;
    rom[44711] = 25'b0000001010000101010111011;
    rom[44712] = 25'b0000001010000101100100100;
    rom[44713] = 25'b0000001010000101110001100;
    rom[44714] = 25'b0000001010000101111110100;
    rom[44715] = 25'b0000001010000110001011010;
    rom[44716] = 25'b0000001010000110011000001;
    rom[44717] = 25'b0000001010000110100100111;
    rom[44718] = 25'b0000001010000110110001100;
    rom[44719] = 25'b0000001010000110111110001;
    rom[44720] = 25'b0000001010000111001010101;
    rom[44721] = 25'b0000001010000111010111001;
    rom[44722] = 25'b0000001010000111100011101;
    rom[44723] = 25'b0000001010000111110000000;
    rom[44724] = 25'b0000001010000111111100010;
    rom[44725] = 25'b0000001010001000001000100;
    rom[44726] = 25'b0000001010001000010100110;
    rom[44727] = 25'b0000001010001000100000110;
    rom[44728] = 25'b0000001010001000101100111;
    rom[44729] = 25'b0000001010001000111000111;
    rom[44730] = 25'b0000001010001001000100111;
    rom[44731] = 25'b0000001010001001010000101;
    rom[44732] = 25'b0000001010001001011100100;
    rom[44733] = 25'b0000001010001001101000010;
    rom[44734] = 25'b0000001010001001110011111;
    rom[44735] = 25'b0000001010001001111111100;
    rom[44736] = 25'b0000001010001010001011000;
    rom[44737] = 25'b0000001010001010010110100;
    rom[44738] = 25'b0000001010001010100001111;
    rom[44739] = 25'b0000001010001010101101011;
    rom[44740] = 25'b0000001010001010111000101;
    rom[44741] = 25'b0000001010001011000011111;
    rom[44742] = 25'b0000001010001011001111000;
    rom[44743] = 25'b0000001010001011011010001;
    rom[44744] = 25'b0000001010001011100101001;
    rom[44745] = 25'b0000001010001011110000001;
    rom[44746] = 25'b0000001010001011111011000;
    rom[44747] = 25'b0000001010001100000110000;
    rom[44748] = 25'b0000001010001100010000101;
    rom[44749] = 25'b0000001010001100011011011;
    rom[44750] = 25'b0000001010001100100110001;
    rom[44751] = 25'b0000001010001100110000110;
    rom[44752] = 25'b0000001010001100111011010;
    rom[44753] = 25'b0000001010001101000101110;
    rom[44754] = 25'b0000001010001101010000001;
    rom[44755] = 25'b0000001010001101011010100;
    rom[44756] = 25'b0000001010001101100100111;
    rom[44757] = 25'b0000001010001101101111001;
    rom[44758] = 25'b0000001010001101111001010;
    rom[44759] = 25'b0000001010001110000011011;
    rom[44760] = 25'b0000001010001110001101100;
    rom[44761] = 25'b0000001010001110010111011;
    rom[44762] = 25'b0000001010001110100001011;
    rom[44763] = 25'b0000001010001110101011001;
    rom[44764] = 25'b0000001010001110110101000;
    rom[44765] = 25'b0000001010001110111110110;
    rom[44766] = 25'b0000001010001111001000011;
    rom[44767] = 25'b0000001010001111010010000;
    rom[44768] = 25'b0000001010001111011011100;
    rom[44769] = 25'b0000001010001111100101000;
    rom[44770] = 25'b0000001010001111101110100;
    rom[44771] = 25'b0000001010001111110111111;
    rom[44772] = 25'b0000001010010000000001001;
    rom[44773] = 25'b0000001010010000001010011;
    rom[44774] = 25'b0000001010010000010011100;
    rom[44775] = 25'b0000001010010000011100101;
    rom[44776] = 25'b0000001010010000100101101;
    rom[44777] = 25'b0000001010010000101110110;
    rom[44778] = 25'b0000001010010000110111101;
    rom[44779] = 25'b0000001010010001000000100;
    rom[44780] = 25'b0000001010010001001001011;
    rom[44781] = 25'b0000001010010001010010000;
    rom[44782] = 25'b0000001010010001011010110;
    rom[44783] = 25'b0000001010010001100011010;
    rom[44784] = 25'b0000001010010001101011111;
    rom[44785] = 25'b0000001010010001110100011;
    rom[44786] = 25'b0000001010010001111100110;
    rom[44787] = 25'b0000001010010010000101010;
    rom[44788] = 25'b0000001010010010001101100;
    rom[44789] = 25'b0000001010010010010101110;
    rom[44790] = 25'b0000001010010010011110000;
    rom[44791] = 25'b0000001010010010100110001;
    rom[44792] = 25'b0000001010010010101110001;
    rom[44793] = 25'b0000001010010010110110001;
    rom[44794] = 25'b0000001010010010111110001;
    rom[44795] = 25'b0000001010010011000101111;
    rom[44796] = 25'b0000001010010011001101110;
    rom[44797] = 25'b0000001010010011010101100;
    rom[44798] = 25'b0000001010010011011101001;
    rom[44799] = 25'b0000001010010011100100111;
    rom[44800] = 25'b0000001010010011101100011;
    rom[44801] = 25'b0000001010010011110011111;
    rom[44802] = 25'b0000001010010011111011011;
    rom[44803] = 25'b0000001010010100000010110;
    rom[44804] = 25'b0000001010010100001010000;
    rom[44805] = 25'b0000001010010100010001010;
    rom[44806] = 25'b0000001010010100011000100;
    rom[44807] = 25'b0000001010010100011111101;
    rom[44808] = 25'b0000001010010100100110101;
    rom[44809] = 25'b0000001010010100101101101;
    rom[44810] = 25'b0000001010010100110100101;
    rom[44811] = 25'b0000001010010100111011101;
    rom[44812] = 25'b0000001010010101000010011;
    rom[44813] = 25'b0000001010010101001001001;
    rom[44814] = 25'b0000001010010101001111111;
    rom[44815] = 25'b0000001010010101010110100;
    rom[44816] = 25'b0000001010010101011101001;
    rom[44817] = 25'b0000001010010101100011101;
    rom[44818] = 25'b0000001010010101101010001;
    rom[44819] = 25'b0000001010010101110000100;
    rom[44820] = 25'b0000001010010101110110110;
    rom[44821] = 25'b0000001010010101111101000;
    rom[44822] = 25'b0000001010010110000011010;
    rom[44823] = 25'b0000001010010110001001100;
    rom[44824] = 25'b0000001010010110001111100;
    rom[44825] = 25'b0000001010010110010101101;
    rom[44826] = 25'b0000001010010110011011100;
    rom[44827] = 25'b0000001010010110100001100;
    rom[44828] = 25'b0000001010010110100111010;
    rom[44829] = 25'b0000001010010110101101000;
    rom[44830] = 25'b0000001010010110110010111;
    rom[44831] = 25'b0000001010010110111000100;
    rom[44832] = 25'b0000001010010110111110000;
    rom[44833] = 25'b0000001010010111000011101;
    rom[44834] = 25'b0000001010010111001001001;
    rom[44835] = 25'b0000001010010111001110100;
    rom[44836] = 25'b0000001010010111010011111;
    rom[44837] = 25'b0000001010010111011001010;
    rom[44838] = 25'b0000001010010111011110100;
    rom[44839] = 25'b0000001010010111100011101;
    rom[44840] = 25'b0000001010010111101000110;
    rom[44841] = 25'b0000001010010111101101110;
    rom[44842] = 25'b0000001010010111110010110;
    rom[44843] = 25'b0000001010010111110111101;
    rom[44844] = 25'b0000001010010111111100101;
    rom[44845] = 25'b0000001010011000000001011;
    rom[44846] = 25'b0000001010011000000110001;
    rom[44847] = 25'b0000001010011000001010111;
    rom[44848] = 25'b0000001010011000001111100;
    rom[44849] = 25'b0000001010011000010100000;
    rom[44850] = 25'b0000001010011000011000100;
    rom[44851] = 25'b0000001010011000011101000;
    rom[44852] = 25'b0000001010011000100001011;
    rom[44853] = 25'b0000001010011000100101110;
    rom[44854] = 25'b0000001010011000101010000;
    rom[44855] = 25'b0000001010011000101110010;
    rom[44856] = 25'b0000001010011000110010011;
    rom[44857] = 25'b0000001010011000110110011;
    rom[44858] = 25'b0000001010011000111010100;
    rom[44859] = 25'b0000001010011000111110011;
    rom[44860] = 25'b0000001010011001000010010;
    rom[44861] = 25'b0000001010011001000110001;
    rom[44862] = 25'b0000001010011001001010000;
    rom[44863] = 25'b0000001010011001001101101;
    rom[44864] = 25'b0000001010011001010001011;
    rom[44865] = 25'b0000001010011001010100111;
    rom[44866] = 25'b0000001010011001011000011;
    rom[44867] = 25'b0000001010011001011100000;
    rom[44868] = 25'b0000001010011001011111011;
    rom[44869] = 25'b0000001010011001100010110;
    rom[44870] = 25'b0000001010011001100110000;
    rom[44871] = 25'b0000001010011001101001010;
    rom[44872] = 25'b0000001010011001101100011;
    rom[44873] = 25'b0000001010011001101111101;
    rom[44874] = 25'b0000001010011001110010101;
    rom[44875] = 25'b0000001010011001110101101;
    rom[44876] = 25'b0000001010011001111000100;
    rom[44877] = 25'b0000001010011001111011100;
    rom[44878] = 25'b0000001010011001111110010;
    rom[44879] = 25'b0000001010011010000001000;
    rom[44880] = 25'b0000001010011010000011110;
    rom[44881] = 25'b0000001010011010000110011;
    rom[44882] = 25'b0000001010011010001000111;
    rom[44883] = 25'b0000001010011010001011011;
    rom[44884] = 25'b0000001010011010001101111;
    rom[44885] = 25'b0000001010011010010000010;
    rom[44886] = 25'b0000001010011010010010110;
    rom[44887] = 25'b0000001010011010010100111;
    rom[44888] = 25'b0000001010011010010111001;
    rom[44889] = 25'b0000001010011010011001011;
    rom[44890] = 25'b0000001010011010011011011;
    rom[44891] = 25'b0000001010011010011101011;
    rom[44892] = 25'b0000001010011010011111011;
    rom[44893] = 25'b0000001010011010100001011;
    rom[44894] = 25'b0000001010011010100011010;
    rom[44895] = 25'b0000001010011010100101000;
    rom[44896] = 25'b0000001010011010100110110;
    rom[44897] = 25'b0000001010011010101000100;
    rom[44898] = 25'b0000001010011010101010000;
    rom[44899] = 25'b0000001010011010101011101;
    rom[44900] = 25'b0000001010011010101101001;
    rom[44901] = 25'b0000001010011010101110101;
    rom[44902] = 25'b0000001010011010110000000;
    rom[44903] = 25'b0000001010011010110001011;
    rom[44904] = 25'b0000001010011010110010100;
    rom[44905] = 25'b0000001010011010110011110;
    rom[44906] = 25'b0000001010011010110101000;
    rom[44907] = 25'b0000001010011010110110000;
    rom[44908] = 25'b0000001010011010110111000;
    rom[44909] = 25'b0000001010011010111000000;
    rom[44910] = 25'b0000001010011010111001000;
    rom[44911] = 25'b0000001010011010111001111;
    rom[44912] = 25'b0000001010011010111010101;
    rom[44913] = 25'b0000001010011010111011011;
    rom[44914] = 25'b0000001010011010111100000;
    rom[44915] = 25'b0000001010011010111100101;
    rom[44916] = 25'b0000001010011010111101001;
    rom[44917] = 25'b0000001010011010111101101;
    rom[44918] = 25'b0000001010011010111110001;
    rom[44919] = 25'b0000001010011010111110100;
    rom[44920] = 25'b0000001010011010111110111;
    rom[44921] = 25'b0000001010011010111111000;
    rom[44922] = 25'b0000001010011010111111011;
    rom[44923] = 25'b0000001010011010111111011;
    rom[44924] = 25'b0000001010011010111111100;
    rom[44925] = 25'b0000001010011010111111100;
    rom[44926] = 25'b0000001010011010111111100;
    rom[44927] = 25'b0000001010011010111111011;
    rom[44928] = 25'b0000001010011010111111011;
    rom[44929] = 25'b0000001010011010111111000;
    rom[44930] = 25'b0000001010011010111110111;
    rom[44931] = 25'b0000001010011010111110100;
    rom[44932] = 25'b0000001010011010111110001;
    rom[44933] = 25'b0000001010011010111101101;
    rom[44934] = 25'b0000001010011010111101001;
    rom[44935] = 25'b0000001010011010111100101;
    rom[44936] = 25'b0000001010011010111100000;
    rom[44937] = 25'b0000001010011010111011011;
    rom[44938] = 25'b0000001010011010111010101;
    rom[44939] = 25'b0000001010011010111001111;
    rom[44940] = 25'b0000001010011010111001000;
    rom[44941] = 25'b0000001010011010111000000;
    rom[44942] = 25'b0000001010011010110111001;
    rom[44943] = 25'b0000001010011010110110001;
    rom[44944] = 25'b0000001010011010110101000;
    rom[44945] = 25'b0000001010011010110011111;
    rom[44946] = 25'b0000001010011010110010101;
    rom[44947] = 25'b0000001010011010110001011;
    rom[44948] = 25'b0000001010011010110000001;
    rom[44949] = 25'b0000001010011010101110110;
    rom[44950] = 25'b0000001010011010101101010;
    rom[44951] = 25'b0000001010011010101011111;
    rom[44952] = 25'b0000001010011010101010010;
    rom[44953] = 25'b0000001010011010101000101;
    rom[44954] = 25'b0000001010011010100111000;
    rom[44955] = 25'b0000001010011010100101010;
    rom[44956] = 25'b0000001010011010100011011;
    rom[44957] = 25'b0000001010011010100001101;
    rom[44958] = 25'b0000001010011010011111110;
    rom[44959] = 25'b0000001010011010011101110;
    rom[44960] = 25'b0000001010011010011011110;
    rom[44961] = 25'b0000001010011010011001110;
    rom[44962] = 25'b0000001010011010010111100;
    rom[44963] = 25'b0000001010011010010101011;
    rom[44964] = 25'b0000001010011010010011001;
    rom[44965] = 25'b0000001010011010010000111;
    rom[44966] = 25'b0000001010011010001110100;
    rom[44967] = 25'b0000001010011010001100000;
    rom[44968] = 25'b0000001010011010001001101;
    rom[44969] = 25'b0000001010011010000111001;
    rom[44970] = 25'b0000001010011010000100100;
    rom[44971] = 25'b0000001010011010000001111;
    rom[44972] = 25'b0000001010011001111111001;
    rom[44973] = 25'b0000001010011001111100011;
    rom[44974] = 25'b0000001010011001111001101;
    rom[44975] = 25'b0000001010011001110110101;
    rom[44976] = 25'b0000001010011001110011110;
    rom[44977] = 25'b0000001010011001110000110;
    rom[44978] = 25'b0000001010011001101101110;
    rom[44979] = 25'b0000001010011001101010101;
    rom[44980] = 25'b0000001010011001100111100;
    rom[44981] = 25'b0000001010011001100100010;
    rom[44982] = 25'b0000001010011001100001000;
    rom[44983] = 25'b0000001010011001011101101;
    rom[44984] = 25'b0000001010011001011010010;
    rom[44985] = 25'b0000001010011001010110111;
    rom[44986] = 25'b0000001010011001010011010;
    rom[44987] = 25'b0000001010011001001111110;
    rom[44988] = 25'b0000001010011001001100001;
    rom[44989] = 25'b0000001010011001001000100;
    rom[44990] = 25'b0000001010011001000100110;
    rom[44991] = 25'b0000001010011001000001000;
    rom[44992] = 25'b0000001010011000111101001;
    rom[44993] = 25'b0000001010011000111001010;
    rom[44994] = 25'b0000001010011000110101010;
    rom[44995] = 25'b0000001010011000110001010;
    rom[44996] = 25'b0000001010011000101101001;
    rom[44997] = 25'b0000001010011000101001001;
    rom[44998] = 25'b0000001010011000100100111;
    rom[44999] = 25'b0000001010011000100000101;
    rom[45000] = 25'b0000001010011000011100011;
    rom[45001] = 25'b0000001010011000011000000;
    rom[45002] = 25'b0000001010011000010011101;
    rom[45003] = 25'b0000001010011000001111001;
    rom[45004] = 25'b0000001010011000001010101;
    rom[45005] = 25'b0000001010011000000110000;
    rom[45006] = 25'b0000001010011000000001011;
    rom[45007] = 25'b0000001010010111111100110;
    rom[45008] = 25'b0000001010010111111000000;
    rom[45009] = 25'b0000001010010111110011001;
    rom[45010] = 25'b0000001010010111101110010;
    rom[45011] = 25'b0000001010010111101001011;
    rom[45012] = 25'b0000001010010111100100011;
    rom[45013] = 25'b0000001010010111011111011;
    rom[45014] = 25'b0000001010010111011010010;
    rom[45015] = 25'b0000001010010111010101001;
    rom[45016] = 25'b0000001010010111010000000;
    rom[45017] = 25'b0000001010010111001010101;
    rom[45018] = 25'b0000001010010111000101011;
    rom[45019] = 25'b0000001010010111000000000;
    rom[45020] = 25'b0000001010010110111010101;
    rom[45021] = 25'b0000001010010110110101001;
    rom[45022] = 25'b0000001010010110101111101;
    rom[45023] = 25'b0000001010010110101010001;
    rom[45024] = 25'b0000001010010110100100011;
    rom[45025] = 25'b0000001010010110011110101;
    rom[45026] = 25'b0000001010010110011001000;
    rom[45027] = 25'b0000001010010110010011001;
    rom[45028] = 25'b0000001010010110001101010;
    rom[45029] = 25'b0000001010010110000111011;
    rom[45030] = 25'b0000001010010110000001011;
    rom[45031] = 25'b0000001010010101111011011;
    rom[45032] = 25'b0000001010010101110101010;
    rom[45033] = 25'b0000001010010101101111001;
    rom[45034] = 25'b0000001010010101101000111;
    rom[45035] = 25'b0000001010010101100010101;
    rom[45036] = 25'b0000001010010101011100011;
    rom[45037] = 25'b0000001010010101010110000;
    rom[45038] = 25'b0000001010010101001111101;
    rom[45039] = 25'b0000001010010101001001001;
    rom[45040] = 25'b0000001010010101000010101;
    rom[45041] = 25'b0000001010010100111100000;
    rom[45042] = 25'b0000001010010100110101011;
    rom[45043] = 25'b0000001010010100101110110;
    rom[45044] = 25'b0000001010010100100111111;
    rom[45045] = 25'b0000001010010100100001001;
    rom[45046] = 25'b0000001010010100011010010;
    rom[45047] = 25'b0000001010010100010011011;
    rom[45048] = 25'b0000001010010100001100011;
    rom[45049] = 25'b0000001010010100000101011;
    rom[45050] = 25'b0000001010010011111110010;
    rom[45051] = 25'b0000001010010011110111001;
    rom[45052] = 25'b0000001010010011110000000;
    rom[45053] = 25'b0000001010010011101000101;
    rom[45054] = 25'b0000001010010011100001011;
    rom[45055] = 25'b0000001010010011011010001;
    rom[45056] = 25'b0000001010010011010010101;
    rom[45057] = 25'b0000001010010011001011001;
    rom[45058] = 25'b0000001010010011000011101;
    rom[45059] = 25'b0000001010010010111100001;
    rom[45060] = 25'b0000001010010010110100100;
    rom[45061] = 25'b0000001010010010101100110;
    rom[45062] = 25'b0000001010010010100101000;
    rom[45063] = 25'b0000001010010010011101010;
    rom[45064] = 25'b0000001010010010010101100;
    rom[45065] = 25'b0000001010010010001101100;
    rom[45066] = 25'b0000001010010010000101101;
    rom[45067] = 25'b0000001010010001111101101;
    rom[45068] = 25'b0000001010010001110101100;
    rom[45069] = 25'b0000001010010001101101011;
    rom[45070] = 25'b0000001010010001100101010;
    rom[45071] = 25'b0000001010010001011101000;
    rom[45072] = 25'b0000001010010001010100110;
    rom[45073] = 25'b0000001010010001001100011;
    rom[45074] = 25'b0000001010010001000100001;
    rom[45075] = 25'b0000001010010000111011101;
    rom[45076] = 25'b0000001010010000110011001;
    rom[45077] = 25'b0000001010010000101010101;
    rom[45078] = 25'b0000001010010000100010000;
    rom[45079] = 25'b0000001010010000011001011;
    rom[45080] = 25'b0000001010010000010000101;
    rom[45081] = 25'b0000001010010000000111111;
    rom[45082] = 25'b0000001010001111111111001;
    rom[45083] = 25'b0000001010001111110110010;
    rom[45084] = 25'b0000001010001111101101010;
    rom[45085] = 25'b0000001010001111100100010;
    rom[45086] = 25'b0000001010001111011011011;
    rom[45087] = 25'b0000001010001111010010001;
    rom[45088] = 25'b0000001010001111001001001;
    rom[45089] = 25'b0000001010001110111111111;
    rom[45090] = 25'b0000001010001110110110101;
    rom[45091] = 25'b0000001010001110101101011;
    rom[45092] = 25'b0000001010001110100100000;
    rom[45093] = 25'b0000001010001110011010101;
    rom[45094] = 25'b0000001010001110010001001;
    rom[45095] = 25'b0000001010001110000111101;
    rom[45096] = 25'b0000001010001101111110001;
    rom[45097] = 25'b0000001010001101110100100;
    rom[45098] = 25'b0000001010001101101010110;
    rom[45099] = 25'b0000001010001101100001001;
    rom[45100] = 25'b0000001010001101010111011;
    rom[45101] = 25'b0000001010001101001101101;
    rom[45102] = 25'b0000001010001101000011101;
    rom[45103] = 25'b0000001010001100111001101;
    rom[45104] = 25'b0000001010001100101111110;
    rom[45105] = 25'b0000001010001100100101110;
    rom[45106] = 25'b0000001010001100011011101;
    rom[45107] = 25'b0000001010001100010001100;
    rom[45108] = 25'b0000001010001100000111010;
    rom[45109] = 25'b0000001010001011111101001;
    rom[45110] = 25'b0000001010001011110010110;
    rom[45111] = 25'b0000001010001011101000011;
    rom[45112] = 25'b0000001010001011011110000;
    rom[45113] = 25'b0000001010001011010011100;
    rom[45114] = 25'b0000001010001011001001000;
    rom[45115] = 25'b0000001010001010111110100;
    rom[45116] = 25'b0000001010001010110011111;
    rom[45117] = 25'b0000001010001010101001010;
    rom[45118] = 25'b0000001010001010011110100;
    rom[45119] = 25'b0000001010001010010011110;
    rom[45120] = 25'b0000001010001010001000111;
    rom[45121] = 25'b0000001010001001111110001;
    rom[45122] = 25'b0000001010001001110011001;
    rom[45123] = 25'b0000001010001001101000001;
    rom[45124] = 25'b0000001010001001011101001;
    rom[45125] = 25'b0000001010001001010010000;
    rom[45126] = 25'b0000001010001001000110111;
    rom[45127] = 25'b0000001010001000111011101;
    rom[45128] = 25'b0000001010001000110000100;
    rom[45129] = 25'b0000001010001000100101001;
    rom[45130] = 25'b0000001010001000011001111;
    rom[45131] = 25'b0000001010001000001110100;
    rom[45132] = 25'b0000001010001000000011000;
    rom[45133] = 25'b0000001010000111110111100;
    rom[45134] = 25'b0000001010000111101011111;
    rom[45135] = 25'b0000001010000111100000011;
    rom[45136] = 25'b0000001010000111010100110;
    rom[45137] = 25'b0000001010000111001001000;
    rom[45138] = 25'b0000001010000110111101010;
    rom[45139] = 25'b0000001010000110110001100;
    rom[45140] = 25'b0000001010000110100101101;
    rom[45141] = 25'b0000001010000110011001110;
    rom[45142] = 25'b0000001010000110001101110;
    rom[45143] = 25'b0000001010000110000001110;
    rom[45144] = 25'b0000001010000101110101101;
    rom[45145] = 25'b0000001010000101101001100;
    rom[45146] = 25'b0000001010000101011101011;
    rom[45147] = 25'b0000001010000101010001001;
    rom[45148] = 25'b0000001010000101000101000;
    rom[45149] = 25'b0000001010000100111000101;
    rom[45150] = 25'b0000001010000100101100010;
    rom[45151] = 25'b0000001010000100011111111;
    rom[45152] = 25'b0000001010000100010011011;
    rom[45153] = 25'b0000001010000100000110111;
    rom[45154] = 25'b0000001010000011111010010;
    rom[45155] = 25'b0000001010000011101101101;
    rom[45156] = 25'b0000001010000011100001000;
    rom[45157] = 25'b0000001010000011010100010;
    rom[45158] = 25'b0000001010000011000111100;
    rom[45159] = 25'b0000001010000010111010101;
    rom[45160] = 25'b0000001010000010101101111;
    rom[45161] = 25'b0000001010000010100000111;
    rom[45162] = 25'b0000001010000010010011111;
    rom[45163] = 25'b0000001010000010000110111;
    rom[45164] = 25'b0000001010000001111001111;
    rom[45165] = 25'b0000001010000001101100101;
    rom[45166] = 25'b0000001010000001011111100;
    rom[45167] = 25'b0000001010000001010010011;
    rom[45168] = 25'b0000001010000001000101000;
    rom[45169] = 25'b0000001010000000110111110;
    rom[45170] = 25'b0000001010000000101010010;
    rom[45171] = 25'b0000001010000000011100111;
    rom[45172] = 25'b0000001010000000001111011;
    rom[45173] = 25'b0000001010000000000001111;
    rom[45174] = 25'b0000001001111111110100010;
    rom[45175] = 25'b0000001001111111100110101;
    rom[45176] = 25'b0000001001111111011001000;
    rom[45177] = 25'b0000001001111111001011010;
    rom[45178] = 25'b0000001001111110111101100;
    rom[45179] = 25'b0000001001111110101111101;
    rom[45180] = 25'b0000001001111110100001111;
    rom[45181] = 25'b0000001001111110010011111;
    rom[45182] = 25'b0000001001111110000101111;
    rom[45183] = 25'b0000001001111101110111111;
    rom[45184] = 25'b0000001001111101101001110;
    rom[45185] = 25'b0000001001111101011011101;
    rom[45186] = 25'b0000001001111101001101100;
    rom[45187] = 25'b0000001001111100111111010;
    rom[45188] = 25'b0000001001111100110001000;
    rom[45189] = 25'b0000001001111100100010110;
    rom[45190] = 25'b0000001001111100010100011;
    rom[45191] = 25'b0000001001111100000110000;
    rom[45192] = 25'b0000001001111011110111100;
    rom[45193] = 25'b0000001001111011101000111;
    rom[45194] = 25'b0000001001111011011010011;
    rom[45195] = 25'b0000001001111011001011110;
    rom[45196] = 25'b0000001001111010111101001;
    rom[45197] = 25'b0000001001111010101110011;
    rom[45198] = 25'b0000001001111010011111101;
    rom[45199] = 25'b0000001001111010010000111;
    rom[45200] = 25'b0000001001111010000010000;
    rom[45201] = 25'b0000001001111001110011000;
    rom[45202] = 25'b0000001001111001100100001;
    rom[45203] = 25'b0000001001111001010101001;
    rom[45204] = 25'b0000001001111001000110000;
    rom[45205] = 25'b0000001001111000110110111;
    rom[45206] = 25'b0000001001111000100111110;
    rom[45207] = 25'b0000001001111000011000101;
    rom[45208] = 25'b0000001001111000001001011;
    rom[45209] = 25'b0000001001110111111010000;
    rom[45210] = 25'b0000001001110111101010110;
    rom[45211] = 25'b0000001001110111011011010;
    rom[45212] = 25'b0000001001110111001011111;
    rom[45213] = 25'b0000001001110110111100011;
    rom[45214] = 25'b0000001001110110101100111;
    rom[45215] = 25'b0000001001110110011101010;
    rom[45216] = 25'b0000001001110110001101101;
    rom[45217] = 25'b0000001001110101111101111;
    rom[45218] = 25'b0000001001110101101110010;
    rom[45219] = 25'b0000001001110101011110100;
    rom[45220] = 25'b0000001001110101001110101;
    rom[45221] = 25'b0000001001110100111110110;
    rom[45222] = 25'b0000001001110100101110111;
    rom[45223] = 25'b0000001001110100011110111;
    rom[45224] = 25'b0000001001110100001110111;
    rom[45225] = 25'b0000001001110011111110111;
    rom[45226] = 25'b0000001001110011101110101;
    rom[45227] = 25'b0000001001110011011110100;
    rom[45228] = 25'b0000001001110011001110010;
    rom[45229] = 25'b0000001001110010111110000;
    rom[45230] = 25'b0000001001110010101101110;
    rom[45231] = 25'b0000001001110010011101011;
    rom[45232] = 25'b0000001001110010001101000;
    rom[45233] = 25'b0000001001110001111100100;
    rom[45234] = 25'b0000001001110001101100001;
    rom[45235] = 25'b0000001001110001011011100;
    rom[45236] = 25'b0000001001110001001011000;
    rom[45237] = 25'b0000001001110000111010011;
    rom[45238] = 25'b0000001001110000101001101;
    rom[45239] = 25'b0000001001110000011000111;
    rom[45240] = 25'b0000001001110000001000001;
    rom[45241] = 25'b0000001001101111110111010;
    rom[45242] = 25'b0000001001101111100110100;
    rom[45243] = 25'b0000001001101111010101101;
    rom[45244] = 25'b0000001001101111000100101;
    rom[45245] = 25'b0000001001101110110011101;
    rom[45246] = 25'b0000001001101110100010100;
    rom[45247] = 25'b0000001001101110010001011;
    rom[45248] = 25'b0000001001101110000000010;
    rom[45249] = 25'b0000001001101101101111000;
    rom[45250] = 25'b0000001001101101011101111;
    rom[45251] = 25'b0000001001101101001100101;
    rom[45252] = 25'b0000001001101100111011010;
    rom[45253] = 25'b0000001001101100101001111;
    rom[45254] = 25'b0000001001101100011000011;
    rom[45255] = 25'b0000001001101100000110111;
    rom[45256] = 25'b0000001001101011110101011;
    rom[45257] = 25'b0000001001101011100011111;
    rom[45258] = 25'b0000001001101011010010010;
    rom[45259] = 25'b0000001001101011000000101;
    rom[45260] = 25'b0000001001101010101110111;
    rom[45261] = 25'b0000001001101010011101001;
    rom[45262] = 25'b0000001001101010001011011;
    rom[45263] = 25'b0000001001101001111001100;
    rom[45264] = 25'b0000001001101001100111101;
    rom[45265] = 25'b0000001001101001010101101;
    rom[45266] = 25'b0000001001101001000011110;
    rom[45267] = 25'b0000001001101000110001110;
    rom[45268] = 25'b0000001001101000011111101;
    rom[45269] = 25'b0000001001101000001101100;
    rom[45270] = 25'b0000001001100111111011011;
    rom[45271] = 25'b0000001001100111101001001;
    rom[45272] = 25'b0000001001100111010110111;
    rom[45273] = 25'b0000001001100111000100100;
    rom[45274] = 25'b0000001001100110110010010;
    rom[45275] = 25'b0000001001100110011111111;
    rom[45276] = 25'b0000001001100110001101011;
    rom[45277] = 25'b0000001001100101111011000;
    rom[45278] = 25'b0000001001100101101000011;
    rom[45279] = 25'b0000001001100101010101110;
    rom[45280] = 25'b0000001001100101000011001;
    rom[45281] = 25'b0000001001100100110000100;
    rom[45282] = 25'b0000001001100100011101111;
    rom[45283] = 25'b0000001001100100001011000;
    rom[45284] = 25'b0000001001100011111000010;
    rom[45285] = 25'b0000001001100011100101011;
    rom[45286] = 25'b0000001001100011010010100;
    rom[45287] = 25'b0000001001100010111111101;
    rom[45288] = 25'b0000001001100010101100101;
    rom[45289] = 25'b0000001001100010011001101;
    rom[45290] = 25'b0000001001100010000110100;
    rom[45291] = 25'b0000001001100001110011100;
    rom[45292] = 25'b0000001001100001100000011;
    rom[45293] = 25'b0000001001100001001101001;
    rom[45294] = 25'b0000001001100000111001111;
    rom[45295] = 25'b0000001001100000100110100;
    rom[45296] = 25'b0000001001100000010011010;
    rom[45297] = 25'b0000001001011111111111111;
    rom[45298] = 25'b0000001001011111101100100;
    rom[45299] = 25'b0000001001011111011001000;
    rom[45300] = 25'b0000001001011111000101100;
    rom[45301] = 25'b0000001001011110110001111;
    rom[45302] = 25'b0000001001011110011110010;
    rom[45303] = 25'b0000001001011110001010101;
    rom[45304] = 25'b0000001001011101110111000;
    rom[45305] = 25'b0000001001011101100011010;
    rom[45306] = 25'b0000001001011101001111100;
    rom[45307] = 25'b0000001001011100111011101;
    rom[45308] = 25'b0000001001011100100111111;
    rom[45309] = 25'b0000001001011100010011111;
    rom[45310] = 25'b0000001001011100000000000;
    rom[45311] = 25'b0000001001011011101100000;
    rom[45312] = 25'b0000001001011011010111111;
    rom[45313] = 25'b0000001001011011000011111;
    rom[45314] = 25'b0000001001011010101111110;
    rom[45315] = 25'b0000001001011010011011101;
    rom[45316] = 25'b0000001001011010000111011;
    rom[45317] = 25'b0000001001011001110011001;
    rom[45318] = 25'b0000001001011001011110111;
    rom[45319] = 25'b0000001001011001001010100;
    rom[45320] = 25'b0000001001011000110110001;
    rom[45321] = 25'b0000001001011000100001101;
    rom[45322] = 25'b0000001001011000001101010;
    rom[45323] = 25'b0000001001010111111000110;
    rom[45324] = 25'b0000001001010111100100010;
    rom[45325] = 25'b0000001001010111001111100;
    rom[45326] = 25'b0000001001010110111010111;
    rom[45327] = 25'b0000001001010110100110010;
    rom[45328] = 25'b0000001001010110010001100;
    rom[45329] = 25'b0000001001010101111100110;
    rom[45330] = 25'b0000001001010101100111111;
    rom[45331] = 25'b0000001001010101010011001;
    rom[45332] = 25'b0000001001010100111110001;
    rom[45333] = 25'b0000001001010100101001010;
    rom[45334] = 25'b0000001001010100010100010;
    rom[45335] = 25'b0000001001010011111111010;
    rom[45336] = 25'b0000001001010011101010010;
    rom[45337] = 25'b0000001001010011010101001;
    rom[45338] = 25'b0000001001010010111111111;
    rom[45339] = 25'b0000001001010010101010110;
    rom[45340] = 25'b0000001001010010010101100;
    rom[45341] = 25'b0000001001010010000000010;
    rom[45342] = 25'b0000001001010001101010111;
    rom[45343] = 25'b0000001001010001010101100;
    rom[45344] = 25'b0000001001010001000000001;
    rom[45345] = 25'b0000001001010000101010101;
    rom[45346] = 25'b0000001001010000010101001;
    rom[45347] = 25'b0000001001001111111111110;
    rom[45348] = 25'b0000001001001111101010001;
    rom[45349] = 25'b0000001001001111010100100;
    rom[45350] = 25'b0000001001001110111110110;
    rom[45351] = 25'b0000001001001110101001001;
    rom[45352] = 25'b0000001001001110010011011;
    rom[45353] = 25'b0000001001001101111101101;
    rom[45354] = 25'b0000001001001101100111110;
    rom[45355] = 25'b0000001001001101010001111;
    rom[45356] = 25'b0000001001001100111100000;
    rom[45357] = 25'b0000001001001100100110001;
    rom[45358] = 25'b0000001001001100010000001;
    rom[45359] = 25'b0000001001001011111010000;
    rom[45360] = 25'b0000001001001011100100000;
    rom[45361] = 25'b0000001001001011001101111;
    rom[45362] = 25'b0000001001001010110111110;
    rom[45363] = 25'b0000001001001010100001100;
    rom[45364] = 25'b0000001001001010001011010;
    rom[45365] = 25'b0000001001001001110101000;
    rom[45366] = 25'b0000001001001001011110110;
    rom[45367] = 25'b0000001001001001001000011;
    rom[45368] = 25'b0000001001001000110001111;
    rom[45369] = 25'b0000001001001000011011100;
    rom[45370] = 25'b0000001001001000000101001;
    rom[45371] = 25'b0000001001000111101110100;
    rom[45372] = 25'b0000001001000111011000000;
    rom[45373] = 25'b0000001001000111000001011;
    rom[45374] = 25'b0000001001000110101010101;
    rom[45375] = 25'b0000001001000110010100000;
    rom[45376] = 25'b0000001001000101111101010;
    rom[45377] = 25'b0000001001000101100110100;
    rom[45378] = 25'b0000001001000101001111110;
    rom[45379] = 25'b0000001001000100111000111;
    rom[45380] = 25'b0000001001000100100010000;
    rom[45381] = 25'b0000001001000100001011001;
    rom[45382] = 25'b0000001001000011110100001;
    rom[45383] = 25'b0000001001000011011101001;
    rom[45384] = 25'b0000001001000011000110001;
    rom[45385] = 25'b0000001001000010101111000;
    rom[45386] = 25'b0000001001000010010111111;
    rom[45387] = 25'b0000001001000010000000101;
    rom[45388] = 25'b0000001001000001101001100;
    rom[45389] = 25'b0000001001000001010010010;
    rom[45390] = 25'b0000001001000000111011000;
    rom[45391] = 25'b0000001001000000100011101;
    rom[45392] = 25'b0000001001000000001100011;
    rom[45393] = 25'b0000001000111111110100111;
    rom[45394] = 25'b0000001000111111011101100;
    rom[45395] = 25'b0000001000111111000110000;
    rom[45396] = 25'b0000001000111110101110100;
    rom[45397] = 25'b0000001000111110010110111;
    rom[45398] = 25'b0000001000111101111111010;
    rom[45399] = 25'b0000001000111101100111101;
    rom[45400] = 25'b0000001000111101010000000;
    rom[45401] = 25'b0000001000111100111000010;
    rom[45402] = 25'b0000001000111100100000100;
    rom[45403] = 25'b0000001000111100001000110;
    rom[45404] = 25'b0000001000111011110000111;
    rom[45405] = 25'b0000001000111011011001000;
    rom[45406] = 25'b0000001000111011000001001;
    rom[45407] = 25'b0000001000111010101001001;
    rom[45408] = 25'b0000001000111010010001001;
    rom[45409] = 25'b0000001000111001111001001;
    rom[45410] = 25'b0000001000111001100001001;
    rom[45411] = 25'b0000001000111001001001000;
    rom[45412] = 25'b0000001000111000110000110;
    rom[45413] = 25'b0000001000111000011000101;
    rom[45414] = 25'b0000001000111000000000011;
    rom[45415] = 25'b0000001000110111101000001;
    rom[45416] = 25'b0000001000110111001111111;
    rom[45417] = 25'b0000001000110110110111101;
    rom[45418] = 25'b0000001000110110011111010;
    rom[45419] = 25'b0000001000110110000110110;
    rom[45420] = 25'b0000001000110101101110010;
    rom[45421] = 25'b0000001000110101010101110;
    rom[45422] = 25'b0000001000110100111101010;
    rom[45423] = 25'b0000001000110100100100101;
    rom[45424] = 25'b0000001000110100001100001;
    rom[45425] = 25'b0000001000110011110011100;
    rom[45426] = 25'b0000001000110011011010111;
    rom[45427] = 25'b0000001000110011000010001;
    rom[45428] = 25'b0000001000110010101001011;
    rom[45429] = 25'b0000001000110010010000101;
    rom[45430] = 25'b0000001000110001110111110;
    rom[45431] = 25'b0000001000110001011110111;
    rom[45432] = 25'b0000001000110001000110000;
    rom[45433] = 25'b0000001000110000101101000;
    rom[45434] = 25'b0000001000110000010100000;
    rom[45435] = 25'b0000001000101111111011000;
    rom[45436] = 25'b0000001000101111100001111;
    rom[45437] = 25'b0000001000101111001000111;
    rom[45438] = 25'b0000001000101110101111110;
    rom[45439] = 25'b0000001000101110010110101;
    rom[45440] = 25'b0000001000101101111101011;
    rom[45441] = 25'b0000001000101101100100001;
    rom[45442] = 25'b0000001000101101001010111;
    rom[45443] = 25'b0000001000101100110001100;
    rom[45444] = 25'b0000001000101100011000010;
    rom[45445] = 25'b0000001000101011111110111;
    rom[45446] = 25'b0000001000101011100101011;
    rom[45447] = 25'b0000001000101011001011111;
    rom[45448] = 25'b0000001000101010110010011;
    rom[45449] = 25'b0000001000101010011000111;
    rom[45450] = 25'b0000001000101001111111011;
    rom[45451] = 25'b0000001000101001100101110;
    rom[45452] = 25'b0000001000101001001100001;
    rom[45453] = 25'b0000001000101000110010011;
    rom[45454] = 25'b0000001000101000011000110;
    rom[45455] = 25'b0000001000100111111111000;
    rom[45456] = 25'b0000001000100111100101001;
    rom[45457] = 25'b0000001000100111001011010;
    rom[45458] = 25'b0000001000100110110001011;
    rom[45459] = 25'b0000001000100110010111100;
    rom[45460] = 25'b0000001000100101111101110;
    rom[45461] = 25'b0000001000100101100011101;
    rom[45462] = 25'b0000001000100101001001101;
    rom[45463] = 25'b0000001000100100101111101;
    rom[45464] = 25'b0000001000100100010101101;
    rom[45465] = 25'b0000001000100011111011011;
    rom[45466] = 25'b0000001000100011100001010;
    rom[45467] = 25'b0000001000100011000111001;
    rom[45468] = 25'b0000001000100010101100111;
    rom[45469] = 25'b0000001000100010010010101;
    rom[45470] = 25'b0000001000100001111000011;
    rom[45471] = 25'b0000001000100001011110000;
    rom[45472] = 25'b0000001000100001000011101;
    rom[45473] = 25'b0000001000100000101001010;
    rom[45474] = 25'b0000001000100000001110111;
    rom[45475] = 25'b0000001000011111110100011;
    rom[45476] = 25'b0000001000011111011001111;
    rom[45477] = 25'b0000001000011110111111010;
    rom[45478] = 25'b0000001000011110100100110;
    rom[45479] = 25'b0000001000011110001010001;
    rom[45480] = 25'b0000001000011101101111100;
    rom[45481] = 25'b0000001000011101010100111;
    rom[45482] = 25'b0000001000011100111010001;
    rom[45483] = 25'b0000001000011100011111011;
    rom[45484] = 25'b0000001000011100000100101;
    rom[45485] = 25'b0000001000011011101001111;
    rom[45486] = 25'b0000001000011011001110111;
    rom[45487] = 25'b0000001000011010110100000;
    rom[45488] = 25'b0000001000011010011001001;
    rom[45489] = 25'b0000001000011001111110001;
    rom[45490] = 25'b0000001000011001100011001;
    rom[45491] = 25'b0000001000011001001000001;
    rom[45492] = 25'b0000001000011000101101001;
    rom[45493] = 25'b0000001000011000010010000;
    rom[45494] = 25'b0000001000010111110110111;
    rom[45495] = 25'b0000001000010111011011110;
    rom[45496] = 25'b0000001000010111000000101;
    rom[45497] = 25'b0000001000010110100101010;
    rom[45498] = 25'b0000001000010110001010000;
    rom[45499] = 25'b0000001000010101101110110;
    rom[45500] = 25'b0000001000010101010011011;
    rom[45501] = 25'b0000001000010100111000000;
    rom[45502] = 25'b0000001000010100011100101;
    rom[45503] = 25'b0000001000010100000001010;
    rom[45504] = 25'b0000001000010011100101110;
    rom[45505] = 25'b0000001000010011001010010;
    rom[45506] = 25'b0000001000010010101110110;
    rom[45507] = 25'b0000001000010010010011010;
    rom[45508] = 25'b0000001000010001110111101;
    rom[45509] = 25'b0000001000010001011011111;
    rom[45510] = 25'b0000001000010001000000010;
    rom[45511] = 25'b0000001000010000100100100;
    rom[45512] = 25'b0000001000010000001000110;
    rom[45513] = 25'b0000001000001111101101001;
    rom[45514] = 25'b0000001000001111010001011;
    rom[45515] = 25'b0000001000001110110101011;
    rom[45516] = 25'b0000001000001110011001101;
    rom[45517] = 25'b0000001000001101111101101;
    rom[45518] = 25'b0000001000001101100001110;
    rom[45519] = 25'b0000001000001101000101111;
    rom[45520] = 25'b0000001000001100101001110;
    rom[45521] = 25'b0000001000001100001101110;
    rom[45522] = 25'b0000001000001011110001101;
    rom[45523] = 25'b0000001000001011010101101;
    rom[45524] = 25'b0000001000001010111001100;
    rom[45525] = 25'b0000001000001010011101011;
    rom[45526] = 25'b0000001000001010000001001;
    rom[45527] = 25'b0000001000001001100101000;
    rom[45528] = 25'b0000001000001001001000101;
    rom[45529] = 25'b0000001000001000101100011;
    rom[45530] = 25'b0000001000001000010000000;
    rom[45531] = 25'b0000001000000111110011110;
    rom[45532] = 25'b0000001000000111010111011;
    rom[45533] = 25'b0000001000000110111010111;
    rom[45534] = 25'b0000001000000110011110100;
    rom[45535] = 25'b0000001000000110000010000;
    rom[45536] = 25'b0000001000000101100101011;
    rom[45537] = 25'b0000001000000101001001000;
    rom[45538] = 25'b0000001000000100101100011;
    rom[45539] = 25'b0000001000000100001111110;
    rom[45540] = 25'b0000001000000011110011001;
    rom[45541] = 25'b0000001000000011010110100;
    rom[45542] = 25'b0000001000000010111001110;
    rom[45543] = 25'b0000001000000010011101000;
    rom[45544] = 25'b0000001000000010000000010;
    rom[45545] = 25'b0000001000000001100011011;
    rom[45546] = 25'b0000001000000001000110100;
    rom[45547] = 25'b0000001000000000101001110;
    rom[45548] = 25'b0000001000000000001100111;
    rom[45549] = 25'b0000000111111111101111111;
    rom[45550] = 25'b0000000111111111010010111;
    rom[45551] = 25'b0000000111111110110110000;
    rom[45552] = 25'b0000000111111110011001000;
    rom[45553] = 25'b0000000111111101111011111;
    rom[45554] = 25'b0000000111111101011110111;
    rom[45555] = 25'b0000000111111101000001110;
    rom[45556] = 25'b0000000111111100100100101;
    rom[45557] = 25'b0000000111111100000111100;
    rom[45558] = 25'b0000000111111011101010010;
    rom[45559] = 25'b0000000111111011001101000;
    rom[45560] = 25'b0000000111111010101111110;
    rom[45561] = 25'b0000000111111010010010011;
    rom[45562] = 25'b0000000111111001110101001;
    rom[45563] = 25'b0000000111111001010111110;
    rom[45564] = 25'b0000000111111000111010011;
    rom[45565] = 25'b0000000111111000011101000;
    rom[45566] = 25'b0000000111110111111111100;
    rom[45567] = 25'b0000000111110111100010000;
    rom[45568] = 25'b0000000111110111000100100;
    rom[45569] = 25'b0000000111110110100111000;
    rom[45570] = 25'b0000000111110110001001011;
    rom[45571] = 25'b0000000111110101101011110;
    rom[45572] = 25'b0000000111110101001110010;
    rom[45573] = 25'b0000000111110100110000101;
    rom[45574] = 25'b0000000111110100010010111;
    rom[45575] = 25'b0000000111110011110101010;
    rom[45576] = 25'b0000000111110011010111011;
    rom[45577] = 25'b0000000111110010111001101;
    rom[45578] = 25'b0000000111110010011011111;
    rom[45579] = 25'b0000000111110001111110000;
    rom[45580] = 25'b0000000111110001100000001;
    rom[45581] = 25'b0000000111110001000010010;
    rom[45582] = 25'b0000000111110000100100010;
    rom[45583] = 25'b0000000111110000000110011;
    rom[45584] = 25'b0000000111101111101000011;
    rom[45585] = 25'b0000000111101111001010011;
    rom[45586] = 25'b0000000111101110101100011;
    rom[45587] = 25'b0000000111101110001110010;
    rom[45588] = 25'b0000000111101101110000010;
    rom[45589] = 25'b0000000111101101010010001;
    rom[45590] = 25'b0000000111101100110011111;
    rom[45591] = 25'b0000000111101100010101110;
    rom[45592] = 25'b0000000111101011110111100;
    rom[45593] = 25'b0000000111101011011001010;
    rom[45594] = 25'b0000000111101010111011000;
    rom[45595] = 25'b0000000111101010011100110;
    rom[45596] = 25'b0000000111101001111110011;
    rom[45597] = 25'b0000000111101001100000000;
    rom[45598] = 25'b0000000111101001000001101;
    rom[45599] = 25'b0000000111101000100011010;
    rom[45600] = 25'b0000000111101000000100110;
    rom[45601] = 25'b0000000111100111100110011;
    rom[45602] = 25'b0000000111100111000111110;
    rom[45603] = 25'b0000000111100110101001011;
    rom[45604] = 25'b0000000111100110001010110;
    rom[45605] = 25'b0000000111100101101100001;
    rom[45606] = 25'b0000000111100101001101100;
    rom[45607] = 25'b0000000111100100101110111;
    rom[45608] = 25'b0000000111100100010000010;
    rom[45609] = 25'b0000000111100011110001101;
    rom[45610] = 25'b0000000111100011010010111;
    rom[45611] = 25'b0000000111100010110100001;
    rom[45612] = 25'b0000000111100010010101010;
    rom[45613] = 25'b0000000111100001110110100;
    rom[45614] = 25'b0000000111100001010111101;
    rom[45615] = 25'b0000000111100000111000111;
    rom[45616] = 25'b0000000111100000011001111;
    rom[45617] = 25'b0000000111011111111011000;
    rom[45618] = 25'b0000000111011111011100001;
    rom[45619] = 25'b0000000111011110111101001;
    rom[45620] = 25'b0000000111011110011110001;
    rom[45621] = 25'b0000000111011101111111001;
    rom[45622] = 25'b0000000111011101100000001;
    rom[45623] = 25'b0000000111011101000001000;
    rom[45624] = 25'b0000000111011100100001111;
    rom[45625] = 25'b0000000111011100000010110;
    rom[45626] = 25'b0000000111011011100011101;
    rom[45627] = 25'b0000000111011011000100011;
    rom[45628] = 25'b0000000111011010100101010;
    rom[45629] = 25'b0000000111011010000110000;
    rom[45630] = 25'b0000000111011001100110101;
    rom[45631] = 25'b0000000111011001000111011;
    rom[45632] = 25'b0000000111011000101000001;
    rom[45633] = 25'b0000000111011000001000110;
    rom[45634] = 25'b0000000111010111101001011;
    rom[45635] = 25'b0000000111010111001010000;
    rom[45636] = 25'b0000000111010110101010101;
    rom[45637] = 25'b0000000111010110001011001;
    rom[45638] = 25'b0000000111010101101011101;
    rom[45639] = 25'b0000000111010101001100001;
    rom[45640] = 25'b0000000111010100101100101;
    rom[45641] = 25'b0000000111010100001101000;
    rom[45642] = 25'b0000000111010011101101100;
    rom[45643] = 25'b0000000111010011001101110;
    rom[45644] = 25'b0000000111010010101110010;
    rom[45645] = 25'b0000000111010010001110101;
    rom[45646] = 25'b0000000111010001101110111;
    rom[45647] = 25'b0000000111010001001111001;
    rom[45648] = 25'b0000000111010000101111011;
    rom[45649] = 25'b0000000111010000001111101;
    rom[45650] = 25'b0000000111001111101111111;
    rom[45651] = 25'b0000000111001111010000001;
    rom[45652] = 25'b0000000111001110110000010;
    rom[45653] = 25'b0000000111001110010000011;
    rom[45654] = 25'b0000000111001101110000100;
    rom[45655] = 25'b0000000111001101010000100;
    rom[45656] = 25'b0000000111001100110000101;
    rom[45657] = 25'b0000000111001100010000101;
    rom[45658] = 25'b0000000111001011110000110;
    rom[45659] = 25'b0000000111001011010000101;
    rom[45660] = 25'b0000000111001010110000101;
    rom[45661] = 25'b0000000111001010010000100;
    rom[45662] = 25'b0000000111001001110000100;
    rom[45663] = 25'b0000000111001001010000011;
    rom[45664] = 25'b0000000111001000110000010;
    rom[45665] = 25'b0000000111001000010000000;
    rom[45666] = 25'b0000000111000111101111111;
    rom[45667] = 25'b0000000111000111001111101;
    rom[45668] = 25'b0000000111000110101111100;
    rom[45669] = 25'b0000000111000110001111001;
    rom[45670] = 25'b0000000111000101101110111;
    rom[45671] = 25'b0000000111000101001110100;
    rom[45672] = 25'b0000000111000100101110010;
    rom[45673] = 25'b0000000111000100001101111;
    rom[45674] = 25'b0000000111000011101101100;
    rom[45675] = 25'b0000000111000011001101001;
    rom[45676] = 25'b0000000111000010101100101;
    rom[45677] = 25'b0000000111000010001100001;
    rom[45678] = 25'b0000000111000001101011101;
    rom[45679] = 25'b0000000111000001001011001;
    rom[45680] = 25'b0000000111000000101010101;
    rom[45681] = 25'b0000000111000000001010001;
    rom[45682] = 25'b0000000110111111101001101;
    rom[45683] = 25'b0000000110111111001001000;
    rom[45684] = 25'b0000000110111110101000010;
    rom[45685] = 25'b0000000110111110000111110;
    rom[45686] = 25'b0000000110111101100111000;
    rom[45687] = 25'b0000000110111101000110011;
    rom[45688] = 25'b0000000110111100100101100;
    rom[45689] = 25'b0000000110111100000100111;
    rom[45690] = 25'b0000000110111011100100001;
    rom[45691] = 25'b0000000110111011000011011;
    rom[45692] = 25'b0000000110111010100010100;
    rom[45693] = 25'b0000000110111010000001101;
    rom[45694] = 25'b0000000110111001100000110;
    rom[45695] = 25'b0000000110111000111111111;
    rom[45696] = 25'b0000000110111000011111000;
    rom[45697] = 25'b0000000110110111111110001;
    rom[45698] = 25'b0000000110110111011101010;
    rom[45699] = 25'b0000000110110110111100010;
    rom[45700] = 25'b0000000110110110011011010;
    rom[45701] = 25'b0000000110110101111010010;
    rom[45702] = 25'b0000000110110101011001001;
    rom[45703] = 25'b0000000110110100111000001;
    rom[45704] = 25'b0000000110110100010111000;
    rom[45705] = 25'b0000000110110011110101111;
    rom[45706] = 25'b0000000110110011010100111;
    rom[45707] = 25'b0000000110110010110011101;
    rom[45708] = 25'b0000000110110010010010011;
    rom[45709] = 25'b0000000110110001110001010;
    rom[45710] = 25'b0000000110110001010000000;
    rom[45711] = 25'b0000000110110000101110110;
    rom[45712] = 25'b0000000110110000001101100;
    rom[45713] = 25'b0000000110101111101100010;
    rom[45714] = 25'b0000000110101111001011000;
    rom[45715] = 25'b0000000110101110101001101;
    rom[45716] = 25'b0000000110101110001000010;
    rom[45717] = 25'b0000000110101101100111000;
    rom[45718] = 25'b0000000110101101000101100;
    rom[45719] = 25'b0000000110101100100100001;
    rom[45720] = 25'b0000000110101100000010110;
    rom[45721] = 25'b0000000110101011100001010;
    rom[45722] = 25'b0000000110101010111111110;
    rom[45723] = 25'b0000000110101010011110010;
    rom[45724] = 25'b0000000110101001111100110;
    rom[45725] = 25'b0000000110101001011011010;
    rom[45726] = 25'b0000000110101000111001101;
    rom[45727] = 25'b0000000110101000011000000;
    rom[45728] = 25'b0000000110100111110110100;
    rom[45729] = 25'b0000000110100111010100111;
    rom[45730] = 25'b0000000110100110110011010;
    rom[45731] = 25'b0000000110100110010001100;
    rom[45732] = 25'b0000000110100101101111111;
    rom[45733] = 25'b0000000110100101001110001;
    rom[45734] = 25'b0000000110100100101100011;
    rom[45735] = 25'b0000000110100100001010101;
    rom[45736] = 25'b0000000110100011101000111;
    rom[45737] = 25'b0000000110100011000111001;
    rom[45738] = 25'b0000000110100010100101010;
    rom[45739] = 25'b0000000110100010000011011;
    rom[45740] = 25'b0000000110100001100001101;
    rom[45741] = 25'b0000000110100000111111110;
    rom[45742] = 25'b0000000110100000011101110;
    rom[45743] = 25'b0000000110011111111011111;
    rom[45744] = 25'b0000000110011111011001111;
    rom[45745] = 25'b0000000110011110111000000;
    rom[45746] = 25'b0000000110011110010110000;
    rom[45747] = 25'b0000000110011101110100000;
    rom[45748] = 25'b0000000110011101010010000;
    rom[45749] = 25'b0000000110011100110000000;
    rom[45750] = 25'b0000000110011100001110000;
    rom[45751] = 25'b0000000110011011101011111;
    rom[45752] = 25'b0000000110011011001001110;
    rom[45753] = 25'b0000000110011010100111101;
    rom[45754] = 25'b0000000110011010000101100;
    rom[45755] = 25'b0000000110011001100011011;
    rom[45756] = 25'b0000000110011001000001001;
    rom[45757] = 25'b0000000110011000011111000;
    rom[45758] = 25'b0000000110010111111100110;
    rom[45759] = 25'b0000000110010111011010100;
    rom[45760] = 25'b0000000110010110111000010;
    rom[45761] = 25'b0000000110010110010110001;
    rom[45762] = 25'b0000000110010101110011110;
    rom[45763] = 25'b0000000110010101010001011;
    rom[45764] = 25'b0000000110010100101111001;
    rom[45765] = 25'b0000000110010100001100110;
    rom[45766] = 25'b0000000110010011101010011;
    rom[45767] = 25'b0000000110010011001000000;
    rom[45768] = 25'b0000000110010010100101101;
    rom[45769] = 25'b0000000110010010000011001;
    rom[45770] = 25'b0000000110010001100000110;
    rom[45771] = 25'b0000000110010000111110011;
    rom[45772] = 25'b0000000110010000011011111;
    rom[45773] = 25'b0000000110001111111001010;
    rom[45774] = 25'b0000000110001111010110111;
    rom[45775] = 25'b0000000110001110110100010;
    rom[45776] = 25'b0000000110001110010001110;
    rom[45777] = 25'b0000000110001101101111001;
    rom[45778] = 25'b0000000110001101001100100;
    rom[45779] = 25'b0000000110001100101010000;
    rom[45780] = 25'b0000000110001100000111011;
    rom[45781] = 25'b0000000110001011100100110;
    rom[45782] = 25'b0000000110001011000010000;
    rom[45783] = 25'b0000000110001010011111010;
    rom[45784] = 25'b0000000110001001111100101;
    rom[45785] = 25'b0000000110001001011001111;
    rom[45786] = 25'b0000000110001000110111001;
    rom[45787] = 25'b0000000110001000010100100;
    rom[45788] = 25'b0000000110000111110001110;
    rom[45789] = 25'b0000000110000111001110111;
    rom[45790] = 25'b0000000110000110101100001;
    rom[45791] = 25'b0000000110000110001001010;
    rom[45792] = 25'b0000000110000101100110100;
    rom[45793] = 25'b0000000110000101000011101;
    rom[45794] = 25'b0000000110000100100000110;
    rom[45795] = 25'b0000000110000011111101111;
    rom[45796] = 25'b0000000110000011011011000;
    rom[45797] = 25'b0000000110000010111000000;
    rom[45798] = 25'b0000000110000010010101001;
    rom[45799] = 25'b0000000110000001110010001;
    rom[45800] = 25'b0000000110000001001111001;
    rom[45801] = 25'b0000000110000000101100001;
    rom[45802] = 25'b0000000110000000001001001;
    rom[45803] = 25'b0000000101111111100110001;
    rom[45804] = 25'b0000000101111111000011000;
    rom[45805] = 25'b0000000101111110100000000;
    rom[45806] = 25'b0000000101111101111100111;
    rom[45807] = 25'b0000000101111101011001110;
    rom[45808] = 25'b0000000101111100110110110;
    rom[45809] = 25'b0000000101111100010011101;
    rom[45810] = 25'b0000000101111011110000100;
    rom[45811] = 25'b0000000101111011001101010;
    rom[45812] = 25'b0000000101111010101010001;
    rom[45813] = 25'b0000000101111010000111000;
    rom[45814] = 25'b0000000101111001100011110;
    rom[45815] = 25'b0000000101111001000000100;
    rom[45816] = 25'b0000000101111000011101010;
    rom[45817] = 25'b0000000101110111111010000;
    rom[45818] = 25'b0000000101110111010110110;
    rom[45819] = 25'b0000000101110110110011011;
    rom[45820] = 25'b0000000101110110010000001;
    rom[45821] = 25'b0000000101110101101100111;
    rom[45822] = 25'b0000000101110101001001100;
    rom[45823] = 25'b0000000101110100100110001;
    rom[45824] = 25'b0000000101110100000010110;
    rom[45825] = 25'b0000000101110011011111011;
    rom[45826] = 25'b0000000101110010111100000;
    rom[45827] = 25'b0000000101110010011000100;
    rom[45828] = 25'b0000000101110001110101001;
    rom[45829] = 25'b0000000101110001010001101;
    rom[45830] = 25'b0000000101110000101110010;
    rom[45831] = 25'b0000000101110000001010110;
    rom[45832] = 25'b0000000101101111100111010;
    rom[45833] = 25'b0000000101101111000011110;
    rom[45834] = 25'b0000000101101110100000010;
    rom[45835] = 25'b0000000101101101111100110;
    rom[45836] = 25'b0000000101101101011001001;
    rom[45837] = 25'b0000000101101100110101101;
    rom[45838] = 25'b0000000101101100010010000;
    rom[45839] = 25'b0000000101101011101110011;
    rom[45840] = 25'b0000000101101011001010111;
    rom[45841] = 25'b0000000101101010100111001;
    rom[45842] = 25'b0000000101101010000011101;
    rom[45843] = 25'b0000000101101001011111111;
    rom[45844] = 25'b0000000101101000111100010;
    rom[45845] = 25'b0000000101101000011000101;
    rom[45846] = 25'b0000000101100111110100111;
    rom[45847] = 25'b0000000101100111010001001;
    rom[45848] = 25'b0000000101100110101101100;
    rom[45849] = 25'b0000000101100110001001110;
    rom[45850] = 25'b0000000101100101100101111;
    rom[45851] = 25'b0000000101100101000010001;
    rom[45852] = 25'b0000000101100100011110011;
    rom[45853] = 25'b0000000101100011111010101;
    rom[45854] = 25'b0000000101100011010110110;
    rom[45855] = 25'b0000000101100010110011000;
    rom[45856] = 25'b0000000101100010001111001;
    rom[45857] = 25'b0000000101100001101011010;
    rom[45858] = 25'b0000000101100001000111011;
    rom[45859] = 25'b0000000101100000100011100;
    rom[45860] = 25'b0000000101011111111111101;
    rom[45861] = 25'b0000000101011111011011110;
    rom[45862] = 25'b0000000101011110110111110;
    rom[45863] = 25'b0000000101011110010011111;
    rom[45864] = 25'b0000000101011101101111111;
    rom[45865] = 25'b0000000101011101001011111;
    rom[45866] = 25'b0000000101011100101000000;
    rom[45867] = 25'b0000000101011100000100000;
    rom[45868] = 25'b0000000101011011100000000;
    rom[45869] = 25'b0000000101011010111100000;
    rom[45870] = 25'b0000000101011010011000000;
    rom[45871] = 25'b0000000101011001110011111;
    rom[45872] = 25'b0000000101011001001111111;
    rom[45873] = 25'b0000000101011000101011111;
    rom[45874] = 25'b0000000101011000000111110;
    rom[45875] = 25'b0000000101010111100011101;
    rom[45876] = 25'b0000000101010110111111101;
    rom[45877] = 25'b0000000101010110011011100;
    rom[45878] = 25'b0000000101010101110111010;
    rom[45879] = 25'b0000000101010101010011001;
    rom[45880] = 25'b0000000101010100101111000;
    rom[45881] = 25'b0000000101010100001010111;
    rom[45882] = 25'b0000000101010011100110101;
    rom[45883] = 25'b0000000101010011000010100;
    rom[45884] = 25'b0000000101010010011110010;
    rom[45885] = 25'b0000000101010001111010000;
    rom[45886] = 25'b0000000101010001010101110;
    rom[45887] = 25'b0000000101010000110001101;
    rom[45888] = 25'b0000000101010000001101011;
    rom[45889] = 25'b0000000101001111101001001;
    rom[45890] = 25'b0000000101001111000100110;
    rom[45891] = 25'b0000000101001110100000100;
    rom[45892] = 25'b0000000101001101111100010;
    rom[45893] = 25'b0000000101001101010111111;
    rom[45894] = 25'b0000000101001100110011100;
    rom[45895] = 25'b0000000101001100001111010;
    rom[45896] = 25'b0000000101001011101010111;
    rom[45897] = 25'b0000000101001011000110101;
    rom[45898] = 25'b0000000101001010100010001;
    rom[45899] = 25'b0000000101001001111101111;
    rom[45900] = 25'b0000000101001001011001011;
    rom[45901] = 25'b0000000101001000110101000;
    rom[45902] = 25'b0000000101001000010000101;
    rom[45903] = 25'b0000000101000111101100001;
    rom[45904] = 25'b0000000101000111000111110;
    rom[45905] = 25'b0000000101000110100011010;
    rom[45906] = 25'b0000000101000101111110111;
    rom[45907] = 25'b0000000101000101011010011;
    rom[45908] = 25'b0000000101000100110110000;
    rom[45909] = 25'b0000000101000100010001011;
    rom[45910] = 25'b0000000101000011101100111;
    rom[45911] = 25'b0000000101000011001000011;
    rom[45912] = 25'b0000000101000010100011111;
    rom[45913] = 25'b0000000101000001111111011;
    rom[45914] = 25'b0000000101000001011010110;
    rom[45915] = 25'b0000000101000000110110010;
    rom[45916] = 25'b0000000101000000010001101;
    rom[45917] = 25'b0000000100111111101101001;
    rom[45918] = 25'b0000000100111111001000100;
    rom[45919] = 25'b0000000100111110100011111;
    rom[45920] = 25'b0000000100111101111111010;
    rom[45921] = 25'b0000000100111101011010110;
    rom[45922] = 25'b0000000100111100110110001;
    rom[45923] = 25'b0000000100111100010001100;
    rom[45924] = 25'b0000000100111011101100110;
    rom[45925] = 25'b0000000100111011001000001;
    rom[45926] = 25'b0000000100111010100011100;
    rom[45927] = 25'b0000000100111001111110110;
    rom[45928] = 25'b0000000100111001011010001;
    rom[45929] = 25'b0000000100111000110101100;
    rom[45930] = 25'b0000000100111000010000110;
    rom[45931] = 25'b0000000100110111101100000;
    rom[45932] = 25'b0000000100110111000111010;
    rom[45933] = 25'b0000000100110110100010101;
    rom[45934] = 25'b0000000100110101111101110;
    rom[45935] = 25'b0000000100110101011001001;
    rom[45936] = 25'b0000000100110100110100010;
    rom[45937] = 25'b0000000100110100001111100;
    rom[45938] = 25'b0000000100110011101010110;
    rom[45939] = 25'b0000000100110011000110000;
    rom[45940] = 25'b0000000100110010100001010;
    rom[45941] = 25'b0000000100110001111100010;
    rom[45942] = 25'b0000000100110001010111100;
    rom[45943] = 25'b0000000100110000110010110;
    rom[45944] = 25'b0000000100110000001101111;
    rom[45945] = 25'b0000000100101111101001000;
    rom[45946] = 25'b0000000100101111000100001;
    rom[45947] = 25'b0000000100101110011111011;
    rom[45948] = 25'b0000000100101101111010100;
    rom[45949] = 25'b0000000100101101010101101;
    rom[45950] = 25'b0000000100101100110000101;
    rom[45951] = 25'b0000000100101100001011110;
    rom[45952] = 25'b0000000100101011100110111;
    rom[45953] = 25'b0000000100101011000001111;
    rom[45954] = 25'b0000000100101010011101000;
    rom[45955] = 25'b0000000100101001111000001;
    rom[45956] = 25'b0000000100101001010011001;
    rom[45957] = 25'b0000000100101000101110010;
    rom[45958] = 25'b0000000100101000001001010;
    rom[45959] = 25'b0000000100100111100100011;
    rom[45960] = 25'b0000000100100110111111011;
    rom[45961] = 25'b0000000100100110011010011;
    rom[45962] = 25'b0000000100100101110101011;
    rom[45963] = 25'b0000000100100101010000011;
    rom[45964] = 25'b0000000100100100101011011;
    rom[45965] = 25'b0000000100100100000110011;
    rom[45966] = 25'b0000000100100011100001011;
    rom[45967] = 25'b0000000100100010111100011;
    rom[45968] = 25'b0000000100100010010111010;
    rom[45969] = 25'b0000000100100001110010011;
    rom[45970] = 25'b0000000100100001001101010;
    rom[45971] = 25'b0000000100100000101000001;
    rom[45972] = 25'b0000000100100000000011001;
    rom[45973] = 25'b0000000100011111011110000;
    rom[45974] = 25'b0000000100011110111001000;
    rom[45975] = 25'b0000000100011110010011111;
    rom[45976] = 25'b0000000100011101101110110;
    rom[45977] = 25'b0000000100011101001001110;
    rom[45978] = 25'b0000000100011100100100101;
    rom[45979] = 25'b0000000100011011111111100;
    rom[45980] = 25'b0000000100011011011010011;
    rom[45981] = 25'b0000000100011010110101010;
    rom[45982] = 25'b0000000100011010010000001;
    rom[45983] = 25'b0000000100011001101011000;
    rom[45984] = 25'b0000000100011001000101111;
    rom[45985] = 25'b0000000100011000100000101;
    rom[45986] = 25'b0000000100010111111011100;
    rom[45987] = 25'b0000000100010111010110011;
    rom[45988] = 25'b0000000100010110110001001;
    rom[45989] = 25'b0000000100010110001100000;
    rom[45990] = 25'b0000000100010101100110111;
    rom[45991] = 25'b0000000100010101000001101;
    rom[45992] = 25'b0000000100010100011100100;
    rom[45993] = 25'b0000000100010011110111010;
    rom[45994] = 25'b0000000100010011010010000;
    rom[45995] = 25'b0000000100010010101100110;
    rom[45996] = 25'b0000000100010010000111101;
    rom[45997] = 25'b0000000100010001100010011;
    rom[45998] = 25'b0000000100010000111101001;
    rom[45999] = 25'b0000000100010000010111111;
    rom[46000] = 25'b0000000100001111110010101;
    rom[46001] = 25'b0000000100001111001101011;
    rom[46002] = 25'b0000000100001110101000001;
    rom[46003] = 25'b0000000100001110000010111;
    rom[46004] = 25'b0000000100001101011101101;
    rom[46005] = 25'b0000000100001100111000011;
    rom[46006] = 25'b0000000100001100010011001;
    rom[46007] = 25'b0000000100001011101101111;
    rom[46008] = 25'b0000000100001011001000100;
    rom[46009] = 25'b0000000100001010100011010;
    rom[46010] = 25'b0000000100001001111101111;
    rom[46011] = 25'b0000000100001001011000101;
    rom[46012] = 25'b0000000100001000110011011;
    rom[46013] = 25'b0000000100001000001110000;
    rom[46014] = 25'b0000000100000111101000101;
    rom[46015] = 25'b0000000100000111000011011;
    rom[46016] = 25'b0000000100000110011110000;
    rom[46017] = 25'b0000000100000101111000101;
    rom[46018] = 25'b0000000100000101010011010;
    rom[46019] = 25'b0000000100000100101110000;
    rom[46020] = 25'b0000000100000100001000101;
    rom[46021] = 25'b0000000100000011100011011;
    rom[46022] = 25'b0000000100000010111101111;
    rom[46023] = 25'b0000000100000010011000100;
    rom[46024] = 25'b0000000100000001110011001;
    rom[46025] = 25'b0000000100000001001101111;
    rom[46026] = 25'b0000000100000000101000100;
    rom[46027] = 25'b0000000100000000000011001;
    rom[46028] = 25'b0000000011111111011101101;
    rom[46029] = 25'b0000000011111110111000011;
    rom[46030] = 25'b0000000011111110010011000;
    rom[46031] = 25'b0000000011111101101101100;
    rom[46032] = 25'b0000000011111101001000001;
    rom[46033] = 25'b0000000011111100100010110;
    rom[46034] = 25'b0000000011111011111101010;
    rom[46035] = 25'b0000000011111011010111111;
    rom[46036] = 25'b0000000011111010110010100;
    rom[46037] = 25'b0000000011111010001101000;
    rom[46038] = 25'b0000000011111001100111101;
    rom[46039] = 25'b0000000011111001000010010;
    rom[46040] = 25'b0000000011111000011100110;
    rom[46041] = 25'b0000000011110111110111010;
    rom[46042] = 25'b0000000011110111010001111;
    rom[46043] = 25'b0000000011110110101100011;
    rom[46044] = 25'b0000000011110110000111000;
    rom[46045] = 25'b0000000011110101100001100;
    rom[46046] = 25'b0000000011110100111100001;
    rom[46047] = 25'b0000000011110100010110101;
    rom[46048] = 25'b0000000011110011110001001;
    rom[46049] = 25'b0000000011110011001011110;
    rom[46050] = 25'b0000000011110010100110010;
    rom[46051] = 25'b0000000011110010000000111;
    rom[46052] = 25'b0000000011110001011011010;
    rom[46053] = 25'b0000000011110000110101111;
    rom[46054] = 25'b0000000011110000010000011;
    rom[46055] = 25'b0000000011101111101011000;
    rom[46056] = 25'b0000000011101111000101011;
    rom[46057] = 25'b0000000011101110100000000;
    rom[46058] = 25'b0000000011101101111010011;
    rom[46059] = 25'b0000000011101101010101000;
    rom[46060] = 25'b0000000011101100101111011;
    rom[46061] = 25'b0000000011101100001010000;
    rom[46062] = 25'b0000000011101011100100011;
    rom[46063] = 25'b0000000011101010111111000;
    rom[46064] = 25'b0000000011101010011001100;
    rom[46065] = 25'b0000000011101001110100000;
    rom[46066] = 25'b0000000011101001001110100;
    rom[46067] = 25'b0000000011101000101000111;
    rom[46068] = 25'b0000000011101000000011100;
    rom[46069] = 25'b0000000011100111011101111;
    rom[46070] = 25'b0000000011100110111000011;
    rom[46071] = 25'b0000000011100110010010111;
    rom[46072] = 25'b0000000011100101101101011;
    rom[46073] = 25'b0000000011100101000111111;
    rom[46074] = 25'b0000000011100100100010010;
    rom[46075] = 25'b0000000011100011111100110;
    rom[46076] = 25'b0000000011100011010111011;
    rom[46077] = 25'b0000000011100010110001110;
    rom[46078] = 25'b0000000011100010001100010;
    rom[46079] = 25'b0000000011100001100110110;
    rom[46080] = 25'b0000000011100001000001001;
    rom[46081] = 25'b0000000011100000011011101;
    rom[46082] = 25'b0000000011011111110110001;
    rom[46083] = 25'b0000000011011111010000100;
    rom[46084] = 25'b0000000011011110101011000;
    rom[46085] = 25'b0000000011011110000101100;
    rom[46086] = 25'b0000000011011101011111111;
    rom[46087] = 25'b0000000011011100111010011;
    rom[46088] = 25'b0000000011011100010100111;
    rom[46089] = 25'b0000000011011011101111010;
    rom[46090] = 25'b0000000011011011001001110;
    rom[46091] = 25'b0000000011011010100100010;
    rom[46092] = 25'b0000000011011001111110101;
    rom[46093] = 25'b0000000011011001011001001;
    rom[46094] = 25'b0000000011011000110011101;
    rom[46095] = 25'b0000000011011000001110000;
    rom[46096] = 25'b0000000011010111101000100;
    rom[46097] = 25'b0000000011010111000011000;
    rom[46098] = 25'b0000000011010110011101011;
    rom[46099] = 25'b0000000011010101110111111;
    rom[46100] = 25'b0000000011010101010010011;
    rom[46101] = 25'b0000000011010100101100101;
    rom[46102] = 25'b0000000011010100000111001;
    rom[46103] = 25'b0000000011010011100001101;
    rom[46104] = 25'b0000000011010010111100000;
    rom[46105] = 25'b0000000011010010010110100;
    rom[46106] = 25'b0000000011010001110001000;
    rom[46107] = 25'b0000000011010001001011011;
    rom[46108] = 25'b0000000011010000100101111;
    rom[46109] = 25'b0000000011010000000000010;
    rom[46110] = 25'b0000000011001111011010110;
    rom[46111] = 25'b0000000011001110110101001;
    rom[46112] = 25'b0000000011001110001111101;
    rom[46113] = 25'b0000000011001101101010001;
    rom[46114] = 25'b0000000011001101000100100;
    rom[46115] = 25'b0000000011001100011111000;
    rom[46116] = 25'b0000000011001011111001100;
    rom[46117] = 25'b0000000011001011010011111;
    rom[46118] = 25'b0000000011001010101110011;
    rom[46119] = 25'b0000000011001010001000110;
    rom[46120] = 25'b0000000011001001100011010;
    rom[46121] = 25'b0000000011001000111101101;
    rom[46122] = 25'b0000000011001000011000001;
    rom[46123] = 25'b0000000011000111110010101;
    rom[46124] = 25'b0000000011000111001101000;
    rom[46125] = 25'b0000000011000110100111100;
    rom[46126] = 25'b0000000011000110000010000;
    rom[46127] = 25'b0000000011000101011100011;
    rom[46128] = 25'b0000000011000100110110111;
    rom[46129] = 25'b0000000011000100010001011;
    rom[46130] = 25'b0000000011000011101011110;
    rom[46131] = 25'b0000000011000011000110010;
    rom[46132] = 25'b0000000011000010100000110;
    rom[46133] = 25'b0000000011000001111011001;
    rom[46134] = 25'b0000000011000001010101101;
    rom[46135] = 25'b0000000011000000110000001;
    rom[46136] = 25'b0000000011000000001010100;
    rom[46137] = 25'b0000000010111111100101001;
    rom[46138] = 25'b0000000010111110111111100;
    rom[46139] = 25'b0000000010111110011010000;
    rom[46140] = 25'b0000000010111101110100100;
    rom[46141] = 25'b0000000010111101001110111;
    rom[46142] = 25'b0000000010111100101001011;
    rom[46143] = 25'b0000000010111100000011111;
    rom[46144] = 25'b0000000010111011011110011;
    rom[46145] = 25'b0000000010111010111000111;
    rom[46146] = 25'b0000000010111010010011010;
    rom[46147] = 25'b0000000010111001101101111;
    rom[46148] = 25'b0000000010111001001000011;
    rom[46149] = 25'b0000000010111000100010110;
    rom[46150] = 25'b0000000010110111111101011;
    rom[46151] = 25'b0000000010110111010111110;
    rom[46152] = 25'b0000000010110110110010011;
    rom[46153] = 25'b0000000010110110001100110;
    rom[46154] = 25'b0000000010110101100111011;
    rom[46155] = 25'b0000000010110101000001110;
    rom[46156] = 25'b0000000010110100011100011;
    rom[46157] = 25'b0000000010110011110110111;
    rom[46158] = 25'b0000000010110011010001011;
    rom[46159] = 25'b0000000010110010101011111;
    rom[46160] = 25'b0000000010110010000110011;
    rom[46161] = 25'b0000000010110001100000111;
    rom[46162] = 25'b0000000010110000111011011;
    rom[46163] = 25'b0000000010110000010110000;
    rom[46164] = 25'b0000000010101111110000100;
    rom[46165] = 25'b0000000010101111001011000;
    rom[46166] = 25'b0000000010101110100101100;
    rom[46167] = 25'b0000000010101110000000000;
    rom[46168] = 25'b0000000010101101011010101;
    rom[46169] = 25'b0000000010101100110101001;
    rom[46170] = 25'b0000000010101100001111110;
    rom[46171] = 25'b0000000010101011101010010;
    rom[46172] = 25'b0000000010101011000100111;
    rom[46173] = 25'b0000000010101010011111011;
    rom[46174] = 25'b0000000010101001111001111;
    rom[46175] = 25'b0000000010101001010100100;
    rom[46176] = 25'b0000000010101000101111001;
    rom[46177] = 25'b0000000010101000001001101;
    rom[46178] = 25'b0000000010100111100100010;
    rom[46179] = 25'b0000000010100110111110110;
    rom[46180] = 25'b0000000010100110011001011;
    rom[46181] = 25'b0000000010100101110100000;
    rom[46182] = 25'b0000000010100101001110100;
    rom[46183] = 25'b0000000010100100101001001;
    rom[46184] = 25'b0000000010100100000011110;
    rom[46185] = 25'b0000000010100011011110011;
    rom[46186] = 25'b0000000010100010111000111;
    rom[46187] = 25'b0000000010100010010011100;
    rom[46188] = 25'b0000000010100001101110010;
    rom[46189] = 25'b0000000010100001001000110;
    rom[46190] = 25'b0000000010100000100011011;
    rom[46191] = 25'b0000000010011111111110000;
    rom[46192] = 25'b0000000010011111011000110;
    rom[46193] = 25'b0000000010011110110011011;
    rom[46194] = 25'b0000000010011110001110000;
    rom[46195] = 25'b0000000010011101101000101;
    rom[46196] = 25'b0000000010011101000011010;
    rom[46197] = 25'b0000000010011100011101111;
    rom[46198] = 25'b0000000010011011111000101;
    rom[46199] = 25'b0000000010011011010011010;
    rom[46200] = 25'b0000000010011010101101111;
    rom[46201] = 25'b0000000010011010001000100;
    rom[46202] = 25'b0000000010011001100011010;
    rom[46203] = 25'b0000000010011000111101111;
    rom[46204] = 25'b0000000010011000011000101;
    rom[46205] = 25'b0000000010010111110011010;
    rom[46206] = 25'b0000000010010111001110000;
    rom[46207] = 25'b0000000010010110101000101;
    rom[46208] = 25'b0000000010010110000011011;
    rom[46209] = 25'b0000000010010101011110001;
    rom[46210] = 25'b0000000010010100111000110;
    rom[46211] = 25'b0000000010010100010011100;
    rom[46212] = 25'b0000000010010011101110010;
    rom[46213] = 25'b0000000010010011001001000;
    rom[46214] = 25'b0000000010010010100011110;
    rom[46215] = 25'b0000000010010001111110100;
    rom[46216] = 25'b0000000010010001011001010;
    rom[46217] = 25'b0000000010010000110100000;
    rom[46218] = 25'b0000000010010000001110101;
    rom[46219] = 25'b0000000010001111101001100;
    rom[46220] = 25'b0000000010001111000100010;
    rom[46221] = 25'b0000000010001110011111001;
    rom[46222] = 25'b0000000010001101111001111;
    rom[46223] = 25'b0000000010001101010100101;
    rom[46224] = 25'b0000000010001100101111011;
    rom[46225] = 25'b0000000010001100001010010;
    rom[46226] = 25'b0000000010001011100101000;
    rom[46227] = 25'b0000000010001010111111110;
    rom[46228] = 25'b0000000010001010011010101;
    rom[46229] = 25'b0000000010001001110101100;
    rom[46230] = 25'b0000000010001001010000010;
    rom[46231] = 25'b0000000010001000101011001;
    rom[46232] = 25'b0000000010001000000110000;
    rom[46233] = 25'b0000000010000111100000110;
    rom[46234] = 25'b0000000010000110111011110;
    rom[46235] = 25'b0000000010000110010110100;
    rom[46236] = 25'b0000000010000101110001011;
    rom[46237] = 25'b0000000010000101001100010;
    rom[46238] = 25'b0000000010000100100111001;
    rom[46239] = 25'b0000000010000100000010000;
    rom[46240] = 25'b0000000010000011011101000;
    rom[46241] = 25'b0000000010000010110111111;
    rom[46242] = 25'b0000000010000010010010110;
    rom[46243] = 25'b0000000010000001101101101;
    rom[46244] = 25'b0000000010000001001000101;
    rom[46245] = 25'b0000000010000000100011100;
    rom[46246] = 25'b0000000001111111111110100;
    rom[46247] = 25'b0000000001111111011001011;
    rom[46248] = 25'b0000000001111110110100011;
    rom[46249] = 25'b0000000001111110001111011;
    rom[46250] = 25'b0000000001111101101010010;
    rom[46251] = 25'b0000000001111101000101010;
    rom[46252] = 25'b0000000001111100100000001;
    rom[46253] = 25'b0000000001111011111011010;
    rom[46254] = 25'b0000000001111011010110010;
    rom[46255] = 25'b0000000001111010110001001;
    rom[46256] = 25'b0000000001111010001100001;
    rom[46257] = 25'b0000000001111001100111001;
    rom[46258] = 25'b0000000001111001000010010;
    rom[46259] = 25'b0000000001111000011101010;
    rom[46260] = 25'b0000000001110111111000011;
    rom[46261] = 25'b0000000001110111010011011;
    rom[46262] = 25'b0000000001110110101110011;
    rom[46263] = 25'b0000000001110110001001100;
    rom[46264] = 25'b0000000001110101100100100;
    rom[46265] = 25'b0000000001110100111111101;
    rom[46266] = 25'b0000000001110100011010110;
    rom[46267] = 25'b0000000001110011110101110;
    rom[46268] = 25'b0000000001110011010000111;
    rom[46269] = 25'b0000000001110010101100000;
    rom[46270] = 25'b0000000001110010000111001;
    rom[46271] = 25'b0000000001110001100010010;
    rom[46272] = 25'b0000000001110000111101011;
    rom[46273] = 25'b0000000001110000011000100;
    rom[46274] = 25'b0000000001101111110011101;
    rom[46275] = 25'b0000000001101111001110111;
    rom[46276] = 25'b0000000001101110101010000;
    rom[46277] = 25'b0000000001101110000101001;
    rom[46278] = 25'b0000000001101101100000011;
    rom[46279] = 25'b0000000001101100111011100;
    rom[46280] = 25'b0000000001101100010110110;
    rom[46281] = 25'b0000000001101011110010000;
    rom[46282] = 25'b0000000001101011001101001;
    rom[46283] = 25'b0000000001101010101000011;
    rom[46284] = 25'b0000000001101010000011101;
    rom[46285] = 25'b0000000001101001011110111;
    rom[46286] = 25'b0000000001101000111010001;
    rom[46287] = 25'b0000000001101000010101011;
    rom[46288] = 25'b0000000001100111110000110;
    rom[46289] = 25'b0000000001100111001011111;
    rom[46290] = 25'b0000000001100110100111010;
    rom[46291] = 25'b0000000001100110000010100;
    rom[46292] = 25'b0000000001100101011101110;
    rom[46293] = 25'b0000000001100100111001001;
    rom[46294] = 25'b0000000001100100010100100;
    rom[46295] = 25'b0000000001100011101111110;
    rom[46296] = 25'b0000000001100011001011001;
    rom[46297] = 25'b0000000001100010100110100;
    rom[46298] = 25'b0000000001100010000001111;
    rom[46299] = 25'b0000000001100001011101010;
    rom[46300] = 25'b0000000001100000111000100;
    rom[46301] = 25'b0000000001100000010100000;
    rom[46302] = 25'b0000000001011111101111011;
    rom[46303] = 25'b0000000001011111001010111;
    rom[46304] = 25'b0000000001011110100110010;
    rom[46305] = 25'b0000000001011110000001101;
    rom[46306] = 25'b0000000001011101011101001;
    rom[46307] = 25'b0000000001011100111000101;
    rom[46308] = 25'b0000000001011100010100000;
    rom[46309] = 25'b0000000001011011101111100;
    rom[46310] = 25'b0000000001011011001011000;
    rom[46311] = 25'b0000000001011010100110011;
    rom[46312] = 25'b0000000001011010000001111;
    rom[46313] = 25'b0000000001011001011101011;
    rom[46314] = 25'b0000000001011000111001000;
    rom[46315] = 25'b0000000001011000010100100;
    rom[46316] = 25'b0000000001010111110000000;
    rom[46317] = 25'b0000000001010111001011100;
    rom[46318] = 25'b0000000001010110100111001;
    rom[46319] = 25'b0000000001010110000010110;
    rom[46320] = 25'b0000000001010101011110010;
    rom[46321] = 25'b0000000001010100111001111;
    rom[46322] = 25'b0000000001010100010101100;
    rom[46323] = 25'b0000000001010011110001001;
    rom[46324] = 25'b0000000001010011001100101;
    rom[46325] = 25'b0000000001010010101000011;
    rom[46326] = 25'b0000000001010010000100000;
    rom[46327] = 25'b0000000001010001011111110;
    rom[46328] = 25'b0000000001010000111011010;
    rom[46329] = 25'b0000000001010000010111000;
    rom[46330] = 25'b0000000001001111110010110;
    rom[46331] = 25'b0000000001001111001110011;
    rom[46332] = 25'b0000000001001110101010000;
    rom[46333] = 25'b0000000001001110000101111;
    rom[46334] = 25'b0000000001001101100001100;
    rom[46335] = 25'b0000000001001100111101010;
    rom[46336] = 25'b0000000001001100011001000;
    rom[46337] = 25'b0000000001001011110100110;
    rom[46338] = 25'b0000000001001011010000100;
    rom[46339] = 25'b0000000001001010101100011;
    rom[46340] = 25'b0000000001001010001000001;
    rom[46341] = 25'b0000000001001001100100000;
    rom[46342] = 25'b0000000001001000111111110;
    rom[46343] = 25'b0000000001001000011011101;
    rom[46344] = 25'b0000000001000111110111011;
    rom[46345] = 25'b0000000001000111010011010;
    rom[46346] = 25'b0000000001000110101111001;
    rom[46347] = 25'b0000000001000110001011001;
    rom[46348] = 25'b0000000001000101100111000;
    rom[46349] = 25'b0000000001000101000010111;
    rom[46350] = 25'b0000000001000100011110110;
    rom[46351] = 25'b0000000001000011111010110;
    rom[46352] = 25'b0000000001000011010110101;
    rom[46353] = 25'b0000000001000010110010101;
    rom[46354] = 25'b0000000001000010001110101;
    rom[46355] = 25'b0000000001000001101010100;
    rom[46356] = 25'b0000000001000001000110100;
    rom[46357] = 25'b0000000001000000100010100;
    rom[46358] = 25'b0000000000111111111110100;
    rom[46359] = 25'b0000000000111111011010100;
    rom[46360] = 25'b0000000000111110110110101;
    rom[46361] = 25'b0000000000111110010010101;
    rom[46362] = 25'b0000000000111101101110101;
    rom[46363] = 25'b0000000000111101001010111;
    rom[46364] = 25'b0000000000111100100110111;
    rom[46365] = 25'b0000000000111100000010111;
    rom[46366] = 25'b0000000000111011011111000;
    rom[46367] = 25'b0000000000111010111011001;
    rom[46368] = 25'b0000000000111010010111011;
    rom[46369] = 25'b0000000000111001110011100;
    rom[46370] = 25'b0000000000111001001111101;
    rom[46371] = 25'b0000000000111000101011111;
    rom[46372] = 25'b0000000000111000001000000;
    rom[46373] = 25'b0000000000110111100100010;
    rom[46374] = 25'b0000000000110111000000011;
    rom[46375] = 25'b0000000000110110011100101;
    rom[46376] = 25'b0000000000110101111000111;
    rom[46377] = 25'b0000000000110101010101001;
    rom[46378] = 25'b0000000000110100110001011;
    rom[46379] = 25'b0000000000110100001101101;
    rom[46380] = 25'b0000000000110011101001111;
    rom[46381] = 25'b0000000000110011000110010;
    rom[46382] = 25'b0000000000110010100010100;
    rom[46383] = 25'b0000000000110001111110111;
    rom[46384] = 25'b0000000000110001011011010;
    rom[46385] = 25'b0000000000110000110111100;
    rom[46386] = 25'b0000000000110000010011111;
    rom[46387] = 25'b0000000000101111110000010;
    rom[46388] = 25'b0000000000101111001100110;
    rom[46389] = 25'b0000000000101110101001001;
    rom[46390] = 25'b0000000000101110000101101;
    rom[46391] = 25'b0000000000101101100010000;
    rom[46392] = 25'b0000000000101100111110011;
    rom[46393] = 25'b0000000000101100011010111;
    rom[46394] = 25'b0000000000101011110111011;
    rom[46395] = 25'b0000000000101011010011111;
    rom[46396] = 25'b0000000000101010110000011;
    rom[46397] = 25'b0000000000101010001100111;
    rom[46398] = 25'b0000000000101001101001011;
    rom[46399] = 25'b0000000000101001000101111;
    rom[46400] = 25'b0000000000101000100010100;
    rom[46401] = 25'b0000000000100111111111001;
    rom[46402] = 25'b0000000000100111011011101;
    rom[46403] = 25'b0000000000100110111000010;
    rom[46404] = 25'b0000000000100110010100111;
    rom[46405] = 25'b0000000000100101110001100;
    rom[46406] = 25'b0000000000100101001110001;
    rom[46407] = 25'b0000000000100100101010111;
    rom[46408] = 25'b0000000000100100000111100;
    rom[46409] = 25'b0000000000100011100100001;
    rom[46410] = 25'b0000000000100011000000111;
    rom[46411] = 25'b0000000000100010011101100;
    rom[46412] = 25'b0000000000100001111010011;
    rom[46413] = 25'b0000000000100001010111000;
    rom[46414] = 25'b0000000000100000110011111;
    rom[46415] = 25'b0000000000100000010000101;
    rom[46416] = 25'b0000000000011111101101011;
    rom[46417] = 25'b0000000000011111001010010;
    rom[46418] = 25'b0000000000011110100111000;
    rom[46419] = 25'b0000000000011110000011110;
    rom[46420] = 25'b0000000000011101100000110;
    rom[46421] = 25'b0000000000011100111101101;
    rom[46422] = 25'b0000000000011100011010100;
    rom[46423] = 25'b0000000000011011110111011;
    rom[46424] = 25'b0000000000011011010100010;
    rom[46425] = 25'b0000000000011010110001001;
    rom[46426] = 25'b0000000000011010001110001;
    rom[46427] = 25'b0000000000011001101011001;
    rom[46428] = 25'b0000000000011001001000000;
    rom[46429] = 25'b0000000000011000100101000;
    rom[46430] = 25'b0000000000011000000010000;
    rom[46431] = 25'b0000000000010111011111000;
    rom[46432] = 25'b0000000000010110111100001;
    rom[46433] = 25'b0000000000010110011001000;
    rom[46434] = 25'b0000000000010101110110001;
    rom[46435] = 25'b0000000000010101010011010;
    rom[46436] = 25'b0000000000010100110000010;
    rom[46437] = 25'b0000000000010100001101100;
    rom[46438] = 25'b0000000000010011101010100;
    rom[46439] = 25'b0000000000010011000111101;
    rom[46440] = 25'b0000000000010010100100111;
    rom[46441] = 25'b0000000000010010000010000;
    rom[46442] = 25'b0000000000010001011111001;
    rom[46443] = 25'b0000000000010000111100011;
    rom[46444] = 25'b0000000000010000011001101;
    rom[46445] = 25'b0000000000001111110110110;
    rom[46446] = 25'b0000000000001111010100000;
    rom[46447] = 25'b0000000000001110110001010;
    rom[46448] = 25'b0000000000001110001110100;
    rom[46449] = 25'b0000000000001101101011111;
    rom[46450] = 25'b0000000000001101001001001;
    rom[46451] = 25'b0000000000001100100110100;
    rom[46452] = 25'b0000000000001100000011111;
    rom[46453] = 25'b0000000000001011100001010;
    rom[46454] = 25'b0000000000001010111110101;
    rom[46455] = 25'b0000000000001010011100000;
    rom[46456] = 25'b0000000000001001111001011;
    rom[46457] = 25'b0000000000001001010110111;
    rom[46458] = 25'b0000000000001000110100010;
    rom[46459] = 25'b0000000000001000010001110;
    rom[46460] = 25'b0000000000000111101111001;
    rom[46461] = 25'b0000000000000111001100110;
    rom[46462] = 25'b0000000000000110101010001;
    rom[46463] = 25'b0000000000000110000111110;
    rom[46464] = 25'b0000000000000101100101010;
    rom[46465] = 25'b0000000000000101000010110;
    rom[46466] = 25'b0000000000000100100000011;
    rom[46467] = 25'b0000000000000011111110000;
    rom[46468] = 25'b0000000000000011011011101;
    rom[46469] = 25'b0000000000000010111001010;
    rom[46470] = 25'b0000000000000010010110111;
    rom[46471] = 25'b0000000000000001110100100;
    rom[46472] = 25'b0000000000000001010010010;
    rom[46473] = 25'b0000000000000000101111111;
    rom[46474] = 25'b0000000000000000001101101;
    rom[46475] = 25'b1111111111111111101011011;
    rom[46476] = 25'b1111111111111111001001001;
    rom[46477] = 25'b1111111111111110100110111;
    rom[46478] = 25'b1111111111111110000100101;
    rom[46479] = 25'b1111111111111101100010100;
    rom[46480] = 25'b1111111111111101000000010;
    rom[46481] = 25'b1111111111111100011110001;
    rom[46482] = 25'b1111111111111011111100000;
    rom[46483] = 25'b1111111111111011011001110;
    rom[46484] = 25'b1111111111111010110111101;
    rom[46485] = 25'b1111111111111010010101101;
    rom[46486] = 25'b1111111111111001110011100;
    rom[46487] = 25'b1111111111111001010001011;
    rom[46488] = 25'b1111111111111000101111011;
    rom[46489] = 25'b1111111111111000001101011;
    rom[46490] = 25'b1111111111110111101011011;
    rom[46491] = 25'b1111111111110111001001011;
    rom[46492] = 25'b1111111111110110100111011;
    rom[46493] = 25'b1111111111110110000101011;
    rom[46494] = 25'b1111111111110101100011100;
    rom[46495] = 25'b1111111111110101000001100;
    rom[46496] = 25'b1111111111110100011111101;
    rom[46497] = 25'b1111111111110011111101101;
    rom[46498] = 25'b1111111111110011011011111;
    rom[46499] = 25'b1111111111110010111010000;
    rom[46500] = 25'b1111111111110010011000001;
    rom[46501] = 25'b1111111111110001110110011;
    rom[46502] = 25'b1111111111110001010100100;
    rom[46503] = 25'b1111111111110000110010110;
    rom[46504] = 25'b1111111111110000010001000;
    rom[46505] = 25'b1111111111101111101111010;
    rom[46506] = 25'b1111111111101111001101100;
    rom[46507] = 25'b1111111111101110101011110;
    rom[46508] = 25'b1111111111101110001010001;
    rom[46509] = 25'b1111111111101101101000100;
    rom[46510] = 25'b1111111111101101000110110;
    rom[46511] = 25'b1111111111101100100101001;
    rom[46512] = 25'b1111111111101100000011100;
    rom[46513] = 25'b1111111111101011100001111;
    rom[46514] = 25'b1111111111101011000000011;
    rom[46515] = 25'b1111111111101010011110110;
    rom[46516] = 25'b1111111111101001111101010;
    rom[46517] = 25'b1111111111101001011011110;
    rom[46518] = 25'b1111111111101000111010001;
    rom[46519] = 25'b1111111111101000011000110;
    rom[46520] = 25'b1111111111100111110111010;
    rom[46521] = 25'b1111111111100111010101110;
    rom[46522] = 25'b1111111111100110110100011;
    rom[46523] = 25'b1111111111100110010010111;
    rom[46524] = 25'b1111111111100101110001101;
    rom[46525] = 25'b1111111111100101010000001;
    rom[46526] = 25'b1111111111100100101110111;
    rom[46527] = 25'b1111111111100100001101100;
    rom[46528] = 25'b1111111111100011101100010;
    rom[46529] = 25'b1111111111100011001010111;
    rom[46530] = 25'b1111111111100010101001101;
    rom[46531] = 25'b1111111111100010001000011;
    rom[46532] = 25'b1111111111100001100111001;
    rom[46533] = 25'b1111111111100001000101111;
    rom[46534] = 25'b1111111111100000100100101;
    rom[46535] = 25'b1111111111100000000011100;
    rom[46536] = 25'b1111111111011111100010011;
    rom[46537] = 25'b1111111111011111000001010;
    rom[46538] = 25'b1111111111011110100000000;
    rom[46539] = 25'b1111111111011101111111000;
    rom[46540] = 25'b1111111111011101011101111;
    rom[46541] = 25'b1111111111011100111100110;
    rom[46542] = 25'b1111111111011100011011111;
    rom[46543] = 25'b1111111111011011111010110;
    rom[46544] = 25'b1111111111011011011001110;
    rom[46545] = 25'b1111111111011010111000110;
    rom[46546] = 25'b1111111111011010010111110;
    rom[46547] = 25'b1111111111011001110110110;
    rom[46548] = 25'b1111111111011001010101111;
    rom[46549] = 25'b1111111111011000110101000;
    rom[46550] = 25'b1111111111011000010100001;
    rom[46551] = 25'b1111111111010111110011010;
    rom[46552] = 25'b1111111111010111010010011;
    rom[46553] = 25'b1111111111010110110001101;
    rom[46554] = 25'b1111111111010110010000110;
    rom[46555] = 25'b1111111111010101110000000;
    rom[46556] = 25'b1111111111010101001111010;
    rom[46557] = 25'b1111111111010100101110100;
    rom[46558] = 25'b1111111111010100001101101;
    rom[46559] = 25'b1111111111010011101101000;
    rom[46560] = 25'b1111111111010011001100010;
    rom[46561] = 25'b1111111111010010101011101;
    rom[46562] = 25'b1111111111010010001011000;
    rom[46563] = 25'b1111111111010001101010011;
    rom[46564] = 25'b1111111111010001001001110;
    rom[46565] = 25'b1111111111010000101001001;
    rom[46566] = 25'b1111111111010000001000101;
    rom[46567] = 25'b1111111111001111101000001;
    rom[46568] = 25'b1111111111001111000111101;
    rom[46569] = 25'b1111111111001110100111001;
    rom[46570] = 25'b1111111111001110000110101;
    rom[46571] = 25'b1111111111001101100110001;
    rom[46572] = 25'b1111111111001101000101101;
    rom[46573] = 25'b1111111111001100100101010;
    rom[46574] = 25'b1111111111001100000100111;
    rom[46575] = 25'b1111111111001011100100100;
    rom[46576] = 25'b1111111111001011000100001;
    rom[46577] = 25'b1111111111001010100011110;
    rom[46578] = 25'b1111111111001010000011011;
    rom[46579] = 25'b1111111111001001100011001;
    rom[46580] = 25'b1111111111001001000010111;
    rom[46581] = 25'b1111111111001000100010101;
    rom[46582] = 25'b1111111111001000000010011;
    rom[46583] = 25'b1111111111000111100010001;
    rom[46584] = 25'b1111111111000111000010000;
    rom[46585] = 25'b1111111111000110100001110;
    rom[46586] = 25'b1111111111000110000001101;
    rom[46587] = 25'b1111111111000101100001100;
    rom[46588] = 25'b1111111111000101000001011;
    rom[46589] = 25'b1111111111000100100001010;
    rom[46590] = 25'b1111111111000100000001010;
    rom[46591] = 25'b1111111111000011100001010;
    rom[46592] = 25'b1111111111000011000001010;
    rom[46593] = 25'b1111111111000010100001001;
    rom[46594] = 25'b1111111111000010000001010;
    rom[46595] = 25'b1111111111000001100001010;
    rom[46596] = 25'b1111111111000001000001011;
    rom[46597] = 25'b1111111111000000100001011;
    rom[46598] = 25'b1111111111000000000001100;
    rom[46599] = 25'b1111111110111111100001101;
    rom[46600] = 25'b1111111110111111000001110;
    rom[46601] = 25'b1111111110111110100010000;
    rom[46602] = 25'b1111111110111110000010010;
    rom[46603] = 25'b1111111110111101100010011;
    rom[46604] = 25'b1111111110111101000010101;
    rom[46605] = 25'b1111111110111100100010111;
    rom[46606] = 25'b1111111110111100000011001;
    rom[46607] = 25'b1111111110111011100011011;
    rom[46608] = 25'b1111111110111011000011110;
    rom[46609] = 25'b1111111110111010100100001;
    rom[46610] = 25'b1111111110111010000100100;
    rom[46611] = 25'b1111111110111001100100111;
    rom[46612] = 25'b1111111110111001000101011;
    rom[46613] = 25'b1111111110111000100101110;
    rom[46614] = 25'b1111111110111000000110010;
    rom[46615] = 25'b1111111110110111100110101;
    rom[46616] = 25'b1111111110110111000111001;
    rom[46617] = 25'b1111111110110110100111110;
    rom[46618] = 25'b1111111110110110001000010;
    rom[46619] = 25'b1111111110110101101000111;
    rom[46620] = 25'b1111111110110101001001011;
    rom[46621] = 25'b1111111110110100101010000;
    rom[46622] = 25'b1111111110110100001010101;
    rom[46623] = 25'b1111111110110011101011011;
    rom[46624] = 25'b1111111110110011001100000;
    rom[46625] = 25'b1111111110110010101100101;
    rom[46626] = 25'b1111111110110010001101011;
    rom[46627] = 25'b1111111110110001101110001;
    rom[46628] = 25'b1111111110110001001110111;
    rom[46629] = 25'b1111111110110000101111110;
    rom[46630] = 25'b1111111110110000010000100;
    rom[46631] = 25'b1111111110101111110001011;
    rom[46632] = 25'b1111111110101111010010010;
    rom[46633] = 25'b1111111110101110110011000;
    rom[46634] = 25'b1111111110101110010100000;
    rom[46635] = 25'b1111111110101101110101000;
    rom[46636] = 25'b1111111110101101010101111;
    rom[46637] = 25'b1111111110101100110110111;
    rom[46638] = 25'b1111111110101100010111111;
    rom[46639] = 25'b1111111110101011111000111;
    rom[46640] = 25'b1111111110101011011001111;
    rom[46641] = 25'b1111111110101010111011000;
    rom[46642] = 25'b1111111110101010011100001;
    rom[46643] = 25'b1111111110101001111101001;
    rom[46644] = 25'b1111111110101001011110010;
    rom[46645] = 25'b1111111110101000111111100;
    rom[46646] = 25'b1111111110101000100000101;
    rom[46647] = 25'b1111111110101000000001111;
    rom[46648] = 25'b1111111110100111100011001;
    rom[46649] = 25'b1111111110100111000100010;
    rom[46650] = 25'b1111111110100110100101100;
    rom[46651] = 25'b1111111110100110000110111;
    rom[46652] = 25'b1111111110100101101000010;
    rom[46653] = 25'b1111111110100101001001101;
    rom[46654] = 25'b1111111110100100101010111;
    rom[46655] = 25'b1111111110100100001100010;
    rom[46656] = 25'b1111111110100011101101101;
    rom[46657] = 25'b1111111110100011001111001;
    rom[46658] = 25'b1111111110100010110000101;
    rom[46659] = 25'b1111111110100010010010001;
    rom[46660] = 25'b1111111110100001110011101;
    rom[46661] = 25'b1111111110100001010101001;
    rom[46662] = 25'b1111111110100000110110101;
    rom[46663] = 25'b1111111110100000011000010;
    rom[46664] = 25'b1111111110011111111001111;
    rom[46665] = 25'b1111111110011111011011100;
    rom[46666] = 25'b1111111110011110111101001;
    rom[46667] = 25'b1111111110011110011110110;
    rom[46668] = 25'b1111111110011110000000100;
    rom[46669] = 25'b1111111110011101100010001;
    rom[46670] = 25'b1111111110011101000011111;
    rom[46671] = 25'b1111111110011100100101110;
    rom[46672] = 25'b1111111110011100000111100;
    rom[46673] = 25'b1111111110011011101001011;
    rom[46674] = 25'b1111111110011011001011001;
    rom[46675] = 25'b1111111110011010101101000;
    rom[46676] = 25'b1111111110011010001111000;
    rom[46677] = 25'b1111111110011001110000111;
    rom[46678] = 25'b1111111110011001010010110;
    rom[46679] = 25'b1111111110011000110100110;
    rom[46680] = 25'b1111111110011000010110110;
    rom[46681] = 25'b1111111110010111111000110;
    rom[46682] = 25'b1111111110010111011010110;
    rom[46683] = 25'b1111111110010110111100111;
    rom[46684] = 25'b1111111110010110011110111;
    rom[46685] = 25'b1111111110010110000001000;
    rom[46686] = 25'b1111111110010101100011001;
    rom[46687] = 25'b1111111110010101000101010;
    rom[46688] = 25'b1111111110010100100111100;
    rom[46689] = 25'b1111111110010100001001110;
    rom[46690] = 25'b1111111110010011101011111;
    rom[46691] = 25'b1111111110010011001110001;
    rom[46692] = 25'b1111111110010010110000011;
    rom[46693] = 25'b1111111110010010010010110;
    rom[46694] = 25'b1111111110010001110101000;
    rom[46695] = 25'b1111111110010001010111011;
    rom[46696] = 25'b1111111110010000111001111;
    rom[46697] = 25'b1111111110010000011100010;
    rom[46698] = 25'b1111111110001111111110101;
    rom[46699] = 25'b1111111110001111100001001;
    rom[46700] = 25'b1111111110001111000011100;
    rom[46701] = 25'b1111111110001110100110001;
    rom[46702] = 25'b1111111110001110001000101;
    rom[46703] = 25'b1111111110001101101011001;
    rom[46704] = 25'b1111111110001101001101101;
    rom[46705] = 25'b1111111110001100110000011;
    rom[46706] = 25'b1111111110001100010010111;
    rom[46707] = 25'b1111111110001011110101101;
    rom[46708] = 25'b1111111110001011011000010;
    rom[46709] = 25'b1111111110001010111010111;
    rom[46710] = 25'b1111111110001010011101101;
    rom[46711] = 25'b1111111110001010000000011;
    rom[46712] = 25'b1111111110001001100011001;
    rom[46713] = 25'b1111111110001001000101111;
    rom[46714] = 25'b1111111110001000101000110;
    rom[46715] = 25'b1111111110001000001011101;
    rom[46716] = 25'b1111111110000111101110100;
    rom[46717] = 25'b1111111110000111010001011;
    rom[46718] = 25'b1111111110000110110100011;
    rom[46719] = 25'b1111111110000110010111010;
    rom[46720] = 25'b1111111110000101111010010;
    rom[46721] = 25'b1111111110000101011101010;
    rom[46722] = 25'b1111111110000101000000010;
    rom[46723] = 25'b1111111110000100100011010;
    rom[46724] = 25'b1111111110000100000110100;
    rom[46725] = 25'b1111111110000011101001100;
    rom[46726] = 25'b1111111110000011001100101;
    rom[46727] = 25'b1111111110000010101111110;
    rom[46728] = 25'b1111111110000010010011000;
    rom[46729] = 25'b1111111110000001110110001;
    rom[46730] = 25'b1111111110000001011001011;
    rom[46731] = 25'b1111111110000000111100101;
    rom[46732] = 25'b1111111110000000100000000;
    rom[46733] = 25'b1111111110000000000011010;
    rom[46734] = 25'b1111111101111111100110101;
    rom[46735] = 25'b1111111101111111001010000;
    rom[46736] = 25'b1111111101111110101101010;
    rom[46737] = 25'b1111111101111110010000110;
    rom[46738] = 25'b1111111101111101110100001;
    rom[46739] = 25'b1111111101111101010111101;
    rom[46740] = 25'b1111111101111100111011001;
    rom[46741] = 25'b1111111101111100011110101;
    rom[46742] = 25'b1111111101111100000010010;
    rom[46743] = 25'b1111111101111011100101110;
    rom[46744] = 25'b1111111101111011001001011;
    rom[46745] = 25'b1111111101111010101101000;
    rom[46746] = 25'b1111111101111010010000101;
    rom[46747] = 25'b1111111101111001110100010;
    rom[46748] = 25'b1111111101111001011000000;
    rom[46749] = 25'b1111111101111000111011101;
    rom[46750] = 25'b1111111101111000011111100;
    rom[46751] = 25'b1111111101111000000011001;
    rom[46752] = 25'b1111111101110111100111000;
    rom[46753] = 25'b1111111101110111001010111;
    rom[46754] = 25'b1111111101110110101110101;
    rom[46755] = 25'b1111111101110110010010100;
    rom[46756] = 25'b1111111101110101110110011;
    rom[46757] = 25'b1111111101110101011010011;
    rom[46758] = 25'b1111111101110100111110011;
    rom[46759] = 25'b1111111101110100100010011;
    rom[46760] = 25'b1111111101110100000110011;
    rom[46761] = 25'b1111111101110011101010011;
    rom[46762] = 25'b1111111101110011001110011;
    rom[46763] = 25'b1111111101110010110010100;
    rom[46764] = 25'b1111111101110010010110101;
    rom[46765] = 25'b1111111101110001111010111;
    rom[46766] = 25'b1111111101110001011111000;
    rom[46767] = 25'b1111111101110001000011001;
    rom[46768] = 25'b1111111101110000100111011;
    rom[46769] = 25'b1111111101110000001011101;
    rom[46770] = 25'b1111111101101111101111111;
    rom[46771] = 25'b1111111101101111010100010;
    rom[46772] = 25'b1111111101101110111000100;
    rom[46773] = 25'b1111111101101110011100111;
    rom[46774] = 25'b1111111101101110000001011;
    rom[46775] = 25'b1111111101101101100101101;
    rom[46776] = 25'b1111111101101101001010001;
    rom[46777] = 25'b1111111101101100101110101;
    rom[46778] = 25'b1111111101101100010011001;
    rom[46779] = 25'b1111111101101011110111101;
    rom[46780] = 25'b1111111101101011011100001;
    rom[46781] = 25'b1111111101101011000000110;
    rom[46782] = 25'b1111111101101010100101010;
    rom[46783] = 25'b1111111101101010001001111;
    rom[46784] = 25'b1111111101101001101110101;
    rom[46785] = 25'b1111111101101001010011010;
    rom[46786] = 25'b1111111101101000110111111;
    rom[46787] = 25'b1111111101101000011100101;
    rom[46788] = 25'b1111111101101000000001100;
    rom[46789] = 25'b1111111101100111100110010;
    rom[46790] = 25'b1111111101100111001011000;
    rom[46791] = 25'b1111111101100110101111111;
    rom[46792] = 25'b1111111101100110010100110;
    rom[46793] = 25'b1111111101100101111001110;
    rom[46794] = 25'b1111111101100101011110101;
    rom[46795] = 25'b1111111101100101000011100;
    rom[46796] = 25'b1111111101100100101000100;
    rom[46797] = 25'b1111111101100100001101101;
    rom[46798] = 25'b1111111101100011110010101;
    rom[46799] = 25'b1111111101100011010111101;
    rom[46800] = 25'b1111111101100010111100110;
    rom[46801] = 25'b1111111101100010100001110;
    rom[46802] = 25'b1111111101100010000111000;
    rom[46803] = 25'b1111111101100001101100001;
    rom[46804] = 25'b1111111101100001010001010;
    rom[46805] = 25'b1111111101100000110110101;
    rom[46806] = 25'b1111111101100000011011110;
    rom[46807] = 25'b1111111101100000000001001;
    rom[46808] = 25'b1111111101011111100110011;
    rom[46809] = 25'b1111111101011111001011110;
    rom[46810] = 25'b1111111101011110110001001;
    rom[46811] = 25'b1111111101011110010110100;
    rom[46812] = 25'b1111111101011101111011111;
    rom[46813] = 25'b1111111101011101100001011;
    rom[46814] = 25'b1111111101011101000110111;
    rom[46815] = 25'b1111111101011100101100011;
    rom[46816] = 25'b1111111101011100010001111;
    rom[46817] = 25'b1111111101011011110111011;
    rom[46818] = 25'b1111111101011011011101000;
    rom[46819] = 25'b1111111101011011000010101;
    rom[46820] = 25'b1111111101011010101000010;
    rom[46821] = 25'b1111111101011010001110000;
    rom[46822] = 25'b1111111101011001110011101;
    rom[46823] = 25'b1111111101011001011001011;
    rom[46824] = 25'b1111111101011000111111001;
    rom[46825] = 25'b1111111101011000100100111;
    rom[46826] = 25'b1111111101011000001010101;
    rom[46827] = 25'b1111111101010111110000100;
    rom[46828] = 25'b1111111101010111010110011;
    rom[46829] = 25'b1111111101010110111100010;
    rom[46830] = 25'b1111111101010110100010001;
    rom[46831] = 25'b1111111101010110001000001;
    rom[46832] = 25'b1111111101010101101110001;
    rom[46833] = 25'b1111111101010101010100001;
    rom[46834] = 25'b1111111101010100111010001;
    rom[46835] = 25'b1111111101010100100000010;
    rom[46836] = 25'b1111111101010100000110010;
    rom[46837] = 25'b1111111101010011101100011;
    rom[46838] = 25'b1111111101010011010010100;
    rom[46839] = 25'b1111111101010010111000110;
    rom[46840] = 25'b1111111101010010011110111;
    rom[46841] = 25'b1111111101010010000101001;
    rom[46842] = 25'b1111111101010001101011100;
    rom[46843] = 25'b1111111101010001010001101;
    rom[46844] = 25'b1111111101010000111000000;
    rom[46845] = 25'b1111111101010000011110011;
    rom[46846] = 25'b1111111101010000000100110;
    rom[46847] = 25'b1111111101001111101011001;
    rom[46848] = 25'b1111111101001111010001100;
    rom[46849] = 25'b1111111101001110111000000;
    rom[46850] = 25'b1111111101001110011110101;
    rom[46851] = 25'b1111111101001110000101001;
    rom[46852] = 25'b1111111101001101101011101;
    rom[46853] = 25'b1111111101001101010010001;
    rom[46854] = 25'b1111111101001100111000110;
    rom[46855] = 25'b1111111101001100011111011;
    rom[46856] = 25'b1111111101001100000110001;
    rom[46857] = 25'b1111111101001011101100110;
    rom[46858] = 25'b1111111101001011010011100;
    rom[46859] = 25'b1111111101001010111010010;
    rom[46860] = 25'b1111111101001010100001000;
    rom[46861] = 25'b1111111101001010000111110;
    rom[46862] = 25'b1111111101001001101110101;
    rom[46863] = 25'b1111111101001001010101100;
    rom[46864] = 25'b1111111101001000111100011;
    rom[46865] = 25'b1111111101001000100011011;
    rom[46866] = 25'b1111111101001000001010010;
    rom[46867] = 25'b1111111101000111110001001;
    rom[46868] = 25'b1111111101000111011000010;
    rom[46869] = 25'b1111111101000110111111010;
    rom[46870] = 25'b1111111101000110100110010;
    rom[46871] = 25'b1111111101000110001101011;
    rom[46872] = 25'b1111111101000101110100100;
    rom[46873] = 25'b1111111101000101011011101;
    rom[46874] = 25'b1111111101000101000010111;
    rom[46875] = 25'b1111111101000100101010001;
    rom[46876] = 25'b1111111101000100010001011;
    rom[46877] = 25'b1111111101000011111000101;
    rom[46878] = 25'b1111111101000011011111111;
    rom[46879] = 25'b1111111101000011000111001;
    rom[46880] = 25'b1111111101000010101110100;
    rom[46881] = 25'b1111111101000010010101111;
    rom[46882] = 25'b1111111101000001111101010;
    rom[46883] = 25'b1111111101000001100100110;
    rom[46884] = 25'b1111111101000001001100001;
    rom[46885] = 25'b1111111101000000110011110;
    rom[46886] = 25'b1111111101000000011011010;
    rom[46887] = 25'b1111111101000000000010110;
    rom[46888] = 25'b1111111100111111101010011;
    rom[46889] = 25'b1111111100111111010010000;
    rom[46890] = 25'b1111111100111110111001101;
    rom[46891] = 25'b1111111100111110100001011;
    rom[46892] = 25'b1111111100111110001001000;
    rom[46893] = 25'b1111111100111101110000111;
    rom[46894] = 25'b1111111100111101011000100;
    rom[46895] = 25'b1111111100111101000000011;
    rom[46896] = 25'b1111111100111100101000001;
    rom[46897] = 25'b1111111100111100010000000;
    rom[46898] = 25'b1111111100111011110111111;
    rom[46899] = 25'b1111111100111011011111110;
    rom[46900] = 25'b1111111100111011000111110;
    rom[46901] = 25'b1111111100111010101111110;
    rom[46902] = 25'b1111111100111010010111110;
    rom[46903] = 25'b1111111100111001111111110;
    rom[46904] = 25'b1111111100111001100111110;
    rom[46905] = 25'b1111111100111001001111111;
    rom[46906] = 25'b1111111100111000111000000;
    rom[46907] = 25'b1111111100111000100000001;
    rom[46908] = 25'b1111111100111000001000011;
    rom[46909] = 25'b1111111100110111110000100;
    rom[46910] = 25'b1111111100110111011000110;
    rom[46911] = 25'b1111111100110111000001000;
    rom[46912] = 25'b1111111100110110101001011;
    rom[46913] = 25'b1111111100110110010001101;
    rom[46914] = 25'b1111111100110101111010000;
    rom[46915] = 25'b1111111100110101100010011;
    rom[46916] = 25'b1111111100110101001010110;
    rom[46917] = 25'b1111111100110100110011010;
    rom[46918] = 25'b1111111100110100011011110;
    rom[46919] = 25'b1111111100110100000100010;
    rom[46920] = 25'b1111111100110011101100110;
    rom[46921] = 25'b1111111100110011010101010;
    rom[46922] = 25'b1111111100110010111110000;
    rom[46923] = 25'b1111111100110010100110101;
    rom[46924] = 25'b1111111100110010001111010;
    rom[46925] = 25'b1111111100110001110111111;
    rom[46926] = 25'b1111111100110001100000101;
    rom[46927] = 25'b1111111100110001001001011;
    rom[46928] = 25'b1111111100110000110010001;
    rom[46929] = 25'b1111111100110000011010111;
    rom[46930] = 25'b1111111100110000000011110;
    rom[46931] = 25'b1111111100101111101100101;
    rom[46932] = 25'b1111111100101111010101100;
    rom[46933] = 25'b1111111100101110111110011;
    rom[46934] = 25'b1111111100101110100111011;
    rom[46935] = 25'b1111111100101110010000011;
    rom[46936] = 25'b1111111100101101111001011;
    rom[46937] = 25'b1111111100101101100010100;
    rom[46938] = 25'b1111111100101101001011101;
    rom[46939] = 25'b1111111100101100110100101;
    rom[46940] = 25'b1111111100101100011101110;
    rom[46941] = 25'b1111111100101100000110111;
    rom[46942] = 25'b1111111100101011110000001;
    rom[46943] = 25'b1111111100101011011001011;
    rom[46944] = 25'b1111111100101011000010101;
    rom[46945] = 25'b1111111100101010101011111;
    rom[46946] = 25'b1111111100101010010101010;
    rom[46947] = 25'b1111111100101001111110101;
    rom[46948] = 25'b1111111100101001101000000;
    rom[46949] = 25'b1111111100101001010001011;
    rom[46950] = 25'b1111111100101000111010110;
    rom[46951] = 25'b1111111100101000100100010;
    rom[46952] = 25'b1111111100101000001101110;
    rom[46953] = 25'b1111111100100111110111011;
    rom[46954] = 25'b1111111100100111100000111;
    rom[46955] = 25'b1111111100100111001010100;
    rom[46956] = 25'b1111111100100110110100001;
    rom[46957] = 25'b1111111100100110011101110;
    rom[46958] = 25'b1111111100100110000111011;
    rom[46959] = 25'b1111111100100101110001001;
    rom[46960] = 25'b1111111100100101011010111;
    rom[46961] = 25'b1111111100100101000100110;
    rom[46962] = 25'b1111111100100100101110100;
    rom[46963] = 25'b1111111100100100011000011;
    rom[46964] = 25'b1111111100100100000010010;
    rom[46965] = 25'b1111111100100011101100001;
    rom[46966] = 25'b1111111100100011010110000;
    rom[46967] = 25'b1111111100100011000000000;
    rom[46968] = 25'b1111111100100010101010000;
    rom[46969] = 25'b1111111100100010010100000;
    rom[46970] = 25'b1111111100100001111110001;
    rom[46971] = 25'b1111111100100001101000001;
    rom[46972] = 25'b1111111100100001010010010;
    rom[46973] = 25'b1111111100100000111100011;
    rom[46974] = 25'b1111111100100000100110101;
    rom[46975] = 25'b1111111100100000010000110;
    rom[46976] = 25'b1111111100011111111011000;
    rom[46977] = 25'b1111111100011111100101010;
    rom[46978] = 25'b1111111100011111001111100;
    rom[46979] = 25'b1111111100011110111001111;
    rom[46980] = 25'b1111111100011110100100010;
    rom[46981] = 25'b1111111100011110001110101;
    rom[46982] = 25'b1111111100011101111001000;
    rom[46983] = 25'b1111111100011101100011100;
    rom[46984] = 25'b1111111100011101001110000;
    rom[46985] = 25'b1111111100011100111000100;
    rom[46986] = 25'b1111111100011100100011000;
    rom[46987] = 25'b1111111100011100001101101;
    rom[46988] = 25'b1111111100011011111000010;
    rom[46989] = 25'b1111111100011011100010111;
    rom[46990] = 25'b1111111100011011001101101;
    rom[46991] = 25'b1111111100011010111000010;
    rom[46992] = 25'b1111111100011010100011000;
    rom[46993] = 25'b1111111100011010001101110;
    rom[46994] = 25'b1111111100011001111000100;
    rom[46995] = 25'b1111111100011001100011011;
    rom[46996] = 25'b1111111100011001001110010;
    rom[46997] = 25'b1111111100011000111001001;
    rom[46998] = 25'b1111111100011000100100000;
    rom[46999] = 25'b1111111100011000001111000;
    rom[47000] = 25'b1111111100010111111010000;
    rom[47001] = 25'b1111111100010111100101000;
    rom[47002] = 25'b1111111100010111010000000;
    rom[47003] = 25'b1111111100010110111011001;
    rom[47004] = 25'b1111111100010110100110010;
    rom[47005] = 25'b1111111100010110010001011;
    rom[47006] = 25'b1111111100010101111100100;
    rom[47007] = 25'b1111111100010101100111110;
    rom[47008] = 25'b1111111100010101010010111;
    rom[47009] = 25'b1111111100010100111110001;
    rom[47010] = 25'b1111111100010100101001100;
    rom[47011] = 25'b1111111100010100010100111;
    rom[47012] = 25'b1111111100010100000000001;
    rom[47013] = 25'b1111111100010011101011100;
    rom[47014] = 25'b1111111100010011010111000;
    rom[47015] = 25'b1111111100010011000010100;
    rom[47016] = 25'b1111111100010010101101111;
    rom[47017] = 25'b1111111100010010011001100;
    rom[47018] = 25'b1111111100010010000101000;
    rom[47019] = 25'b1111111100010001110000100;
    rom[47020] = 25'b1111111100010001011100001;
    rom[47021] = 25'b1111111100010001000111111;
    rom[47022] = 25'b1111111100010000110011100;
    rom[47023] = 25'b1111111100010000011111010;
    rom[47024] = 25'b1111111100010000001011000;
    rom[47025] = 25'b1111111100001111110110101;
    rom[47026] = 25'b1111111100001111100010100;
    rom[47027] = 25'b1111111100001111001110011;
    rom[47028] = 25'b1111111100001110111010001;
    rom[47029] = 25'b1111111100001110100110001;
    rom[47030] = 25'b1111111100001110010010000;
    rom[47031] = 25'b1111111100001101111101111;
    rom[47032] = 25'b1111111100001101101010000;
    rom[47033] = 25'b1111111100001101010110000;
    rom[47034] = 25'b1111111100001101000010000;
    rom[47035] = 25'b1111111100001100101110001;
    rom[47036] = 25'b1111111100001100011010010;
    rom[47037] = 25'b1111111100001100000110010;
    rom[47038] = 25'b1111111100001011110010100;
    rom[47039] = 25'b1111111100001011011110110;
    rom[47040] = 25'b1111111100001011001010111;
    rom[47041] = 25'b1111111100001010110111010;
    rom[47042] = 25'b1111111100001010100011100;
    rom[47043] = 25'b1111111100001010001111111;
    rom[47044] = 25'b1111111100001001111100001;
    rom[47045] = 25'b1111111100001001101000101;
    rom[47046] = 25'b1111111100001001010101000;
    rom[47047] = 25'b1111111100001001000001100;
    rom[47048] = 25'b1111111100001000101110000;
    rom[47049] = 25'b1111111100001000011010100;
    rom[47050] = 25'b1111111100001000000111001;
    rom[47051] = 25'b1111111100000111110011101;
    rom[47052] = 25'b1111111100000111100000011;
    rom[47053] = 25'b1111111100000111001101000;
    rom[47054] = 25'b1111111100000110111001101;
    rom[47055] = 25'b1111111100000110100110011;
    rom[47056] = 25'b1111111100000110010011001;
    rom[47057] = 25'b1111111100000101111111111;
    rom[47058] = 25'b1111111100000101101100110;
    rom[47059] = 25'b1111111100000101011001100;
    rom[47060] = 25'b1111111100000101000110011;
    rom[47061] = 25'b1111111100000100110011010;
    rom[47062] = 25'b1111111100000100100000010;
    rom[47063] = 25'b1111111100000100001101010;
    rom[47064] = 25'b1111111100000011111010010;
    rom[47065] = 25'b1111111100000011100111010;
    rom[47066] = 25'b1111111100000011010100010;
    rom[47067] = 25'b1111111100000011000001011;
    rom[47068] = 25'b1111111100000010101110101;
    rom[47069] = 25'b1111111100000010011011110;
    rom[47070] = 25'b1111111100000010001000111;
    rom[47071] = 25'b1111111100000001110110001;
    rom[47072] = 25'b1111111100000001100011011;
    rom[47073] = 25'b1111111100000001010000110;
    rom[47074] = 25'b1111111100000000111110000;
    rom[47075] = 25'b1111111100000000101011011;
    rom[47076] = 25'b1111111100000000011000110;
    rom[47077] = 25'b1111111100000000000110010;
    rom[47078] = 25'b1111111011111111110011101;
    rom[47079] = 25'b1111111011111111100001001;
    rom[47080] = 25'b1111111011111111001110101;
    rom[47081] = 25'b1111111011111110111100001;
    rom[47082] = 25'b1111111011111110101001110;
    rom[47083] = 25'b1111111011111110010111011;
    rom[47084] = 25'b1111111011111110000101000;
    rom[47085] = 25'b1111111011111101110010110;
    rom[47086] = 25'b1111111011111101100000011;
    rom[47087] = 25'b1111111011111101001110001;
    rom[47088] = 25'b1111111011111100111011111;
    rom[47089] = 25'b1111111011111100101001110;
    rom[47090] = 25'b1111111011111100010111101;
    rom[47091] = 25'b1111111011111100000101100;
    rom[47092] = 25'b1111111011111011110011011;
    rom[47093] = 25'b1111111011111011100001010;
    rom[47094] = 25'b1111111011111011001111010;
    rom[47095] = 25'b1111111011111010111101001;
    rom[47096] = 25'b1111111011111010101011010;
    rom[47097] = 25'b1111111011111010011001011;
    rom[47098] = 25'b1111111011111010000111011;
    rom[47099] = 25'b1111111011111001110101100;
    rom[47100] = 25'b1111111011111001100011110;
    rom[47101] = 25'b1111111011111001010001111;
    rom[47102] = 25'b1111111011111001000000001;
    rom[47103] = 25'b1111111011111000101110011;
    rom[47104] = 25'b1111111011111000011100101;
    rom[47105] = 25'b1111111011111000001011000;
    rom[47106] = 25'b1111111011110111111001011;
    rom[47107] = 25'b1111111011110111100111110;
    rom[47108] = 25'b1111111011110111010110001;
    rom[47109] = 25'b1111111011110111000100101;
    rom[47110] = 25'b1111111011110110110011001;
    rom[47111] = 25'b1111111011110110100001101;
    rom[47112] = 25'b1111111011110110010000001;
    rom[47113] = 25'b1111111011110101111110110;
    rom[47114] = 25'b1111111011110101101101011;
    rom[47115] = 25'b1111111011110101011100000;
    rom[47116] = 25'b1111111011110101001010101;
    rom[47117] = 25'b1111111011110100111001011;
    rom[47118] = 25'b1111111011110100101000001;
    rom[47119] = 25'b1111111011110100010110111;
    rom[47120] = 25'b1111111011110100000101110;
    rom[47121] = 25'b1111111011110011110100100;
    rom[47122] = 25'b1111111011110011100011011;
    rom[47123] = 25'b1111111011110011010010011;
    rom[47124] = 25'b1111111011110011000001010;
    rom[47125] = 25'b1111111011110010110000010;
    rom[47126] = 25'b1111111011110010011111010;
    rom[47127] = 25'b1111111011110010001110010;
    rom[47128] = 25'b1111111011110001111101011;
    rom[47129] = 25'b1111111011110001101100100;
    rom[47130] = 25'b1111111011110001011011100;
    rom[47131] = 25'b1111111011110001001010110;
    rom[47132] = 25'b1111111011110000111001111;
    rom[47133] = 25'b1111111011110000101001001;
    rom[47134] = 25'b1111111011110000011000011;
    rom[47135] = 25'b1111111011110000000111110;
    rom[47136] = 25'b1111111011101111110111001;
    rom[47137] = 25'b1111111011101111100110100;
    rom[47138] = 25'b1111111011101111010101111;
    rom[47139] = 25'b1111111011101111000101010;
    rom[47140] = 25'b1111111011101110110100101;
    rom[47141] = 25'b1111111011101110100100010;
    rom[47142] = 25'b1111111011101110010011110;
    rom[47143] = 25'b1111111011101110000011010;
    rom[47144] = 25'b1111111011101101110010111;
    rom[47145] = 25'b1111111011101101100010100;
    rom[47146] = 25'b1111111011101101010010001;
    rom[47147] = 25'b1111111011101101000001110;
    rom[47148] = 25'b1111111011101100110001100;
    rom[47149] = 25'b1111111011101100100001010;
    rom[47150] = 25'b1111111011101100010001000;
    rom[47151] = 25'b1111111011101100000000111;
    rom[47152] = 25'b1111111011101011110000110;
    rom[47153] = 25'b1111111011101011100000101;
    rom[47154] = 25'b1111111011101011010000100;
    rom[47155] = 25'b1111111011101011000000100;
    rom[47156] = 25'b1111111011101010110000100;
    rom[47157] = 25'b1111111011101010100000100;
    rom[47158] = 25'b1111111011101010010000100;
    rom[47159] = 25'b1111111011101010000000101;
    rom[47160] = 25'b1111111011101001110000110;
    rom[47161] = 25'b1111111011101001100000111;
    rom[47162] = 25'b1111111011101001010001000;
    rom[47163] = 25'b1111111011101001000001010;
    rom[47164] = 25'b1111111011101000110001100;
    rom[47165] = 25'b1111111011101000100001110;
    rom[47166] = 25'b1111111011101000010010001;
    rom[47167] = 25'b1111111011101000000010011;
    rom[47168] = 25'b1111111011100111110010111;
    rom[47169] = 25'b1111111011100111100011010;
    rom[47170] = 25'b1111111011100111010011101;
    rom[47171] = 25'b1111111011100111000100001;
    rom[47172] = 25'b1111111011100110110100101;
    rom[47173] = 25'b1111111011100110100101010;
    rom[47174] = 25'b1111111011100110010101110;
    rom[47175] = 25'b1111111011100110000110011;
    rom[47176] = 25'b1111111011100101110111000;
    rom[47177] = 25'b1111111011100101100111101;
    rom[47178] = 25'b1111111011100101011000011;
    rom[47179] = 25'b1111111011100101001001001;
    rom[47180] = 25'b1111111011100100111001111;
    rom[47181] = 25'b1111111011100100101010110;
    rom[47182] = 25'b1111111011100100011011100;
    rom[47183] = 25'b1111111011100100001100011;
    rom[47184] = 25'b1111111011100011111101011;
    rom[47185] = 25'b1111111011100011101110001;
    rom[47186] = 25'b1111111011100011011111001;
    rom[47187] = 25'b1111111011100011010000010;
    rom[47188] = 25'b1111111011100011000001001;
    rom[47189] = 25'b1111111011100010110010010;
    rom[47190] = 25'b1111111011100010100011011;
    rom[47191] = 25'b1111111011100010010100100;
    rom[47192] = 25'b1111111011100010000101101;
    rom[47193] = 25'b1111111011100001110110111;
    rom[47194] = 25'b1111111011100001101000001;
    rom[47195] = 25'b1111111011100001011001011;
    rom[47196] = 25'b1111111011100001001010101;
    rom[47197] = 25'b1111111011100000111100000;
    rom[47198] = 25'b1111111011100000101101011;
    rom[47199] = 25'b1111111011100000011110101;
    rom[47200] = 25'b1111111011100000010000001;
    rom[47201] = 25'b1111111011100000000001101;
    rom[47202] = 25'b1111111011011111110011001;
    rom[47203] = 25'b1111111011011111100100101;
    rom[47204] = 25'b1111111011011111010110010;
    rom[47205] = 25'b1111111011011111000111110;
    rom[47206] = 25'b1111111011011110111001011;
    rom[47207] = 25'b1111111011011110101011001;
    rom[47208] = 25'b1111111011011110011100110;
    rom[47209] = 25'b1111111011011110001110100;
    rom[47210] = 25'b1111111011011110000000010;
    rom[47211] = 25'b1111111011011101110010000;
    rom[47212] = 25'b1111111011011101100011110;
    rom[47213] = 25'b1111111011011101010101110;
    rom[47214] = 25'b1111111011011101000111101;
    rom[47215] = 25'b1111111011011100111001100;
    rom[47216] = 25'b1111111011011100101011011;
    rom[47217] = 25'b1111111011011100011101011;
    rom[47218] = 25'b1111111011011100001111100;
    rom[47219] = 25'b1111111011011100000001100;
    rom[47220] = 25'b1111111011011011110011100;
    rom[47221] = 25'b1111111011011011100101110;
    rom[47222] = 25'b1111111011011011010111111;
    rom[47223] = 25'b1111111011011011001010000;
    rom[47224] = 25'b1111111011011010111100010;
    rom[47225] = 25'b1111111011011010101110100;
    rom[47226] = 25'b1111111011011010100000111;
    rom[47227] = 25'b1111111011011010010011001;
    rom[47228] = 25'b1111111011011010000101100;
    rom[47229] = 25'b1111111011011001110111111;
    rom[47230] = 25'b1111111011011001101010010;
    rom[47231] = 25'b1111111011011001011100110;
    rom[47232] = 25'b1111111011011001001111010;
    rom[47233] = 25'b1111111011011001000001101;
    rom[47234] = 25'b1111111011011000110100010;
    rom[47235] = 25'b1111111011011000100110111;
    rom[47236] = 25'b1111111011011000011001011;
    rom[47237] = 25'b1111111011011000001100000;
    rom[47238] = 25'b1111111011010111111110110;
    rom[47239] = 25'b1111111011010111110001100;
    rom[47240] = 25'b1111111011010111100100010;
    rom[47241] = 25'b1111111011010111010111000;
    rom[47242] = 25'b1111111011010111001001111;
    rom[47243] = 25'b1111111011010110111100101;
    rom[47244] = 25'b1111111011010110101111100;
    rom[47245] = 25'b1111111011010110100010011;
    rom[47246] = 25'b1111111011010110010101011;
    rom[47247] = 25'b1111111011010110001000011;
    rom[47248] = 25'b1111111011010101111011011;
    rom[47249] = 25'b1111111011010101101110011;
    rom[47250] = 25'b1111111011010101100001100;
    rom[47251] = 25'b1111111011010101010100101;
    rom[47252] = 25'b1111111011010101000111110;
    rom[47253] = 25'b1111111011010100111011000;
    rom[47254] = 25'b1111111011010100101110001;
    rom[47255] = 25'b1111111011010100100001011;
    rom[47256] = 25'b1111111011010100010100101;
    rom[47257] = 25'b1111111011010100001000000;
    rom[47258] = 25'b1111111011010011111011010;
    rom[47259] = 25'b1111111011010011101110101;
    rom[47260] = 25'b1111111011010011100010000;
    rom[47261] = 25'b1111111011010011010101100;
    rom[47262] = 25'b1111111011010011001001000;
    rom[47263] = 25'b1111111011010010111100100;
    rom[47264] = 25'b1111111011010010110000000;
    rom[47265] = 25'b1111111011010010100011101;
    rom[47266] = 25'b1111111011010010010111010;
    rom[47267] = 25'b1111111011010010001010111;
    rom[47268] = 25'b1111111011010001111110100;
    rom[47269] = 25'b1111111011010001110010010;
    rom[47270] = 25'b1111111011010001100110000;
    rom[47271] = 25'b1111111011010001011001110;
    rom[47272] = 25'b1111111011010001001101101;
    rom[47273] = 25'b1111111011010001000001011;
    rom[47274] = 25'b1111111011010000110101010;
    rom[47275] = 25'b1111111011010000101001001;
    rom[47276] = 25'b1111111011010000011101001;
    rom[47277] = 25'b1111111011010000010001000;
    rom[47278] = 25'b1111111011010000000101001;
    rom[47279] = 25'b1111111011001111111001000;
    rom[47280] = 25'b1111111011001111101101010;
    rom[47281] = 25'b1111111011001111100001010;
    rom[47282] = 25'b1111111011001111010101011;
    rom[47283] = 25'b1111111011001111001001101;
    rom[47284] = 25'b1111111011001110111101110;
    rom[47285] = 25'b1111111011001110110010000;
    rom[47286] = 25'b1111111011001110100110011;
    rom[47287] = 25'b1111111011001110011010100;
    rom[47288] = 25'b1111111011001110001110111;
    rom[47289] = 25'b1111111011001110000011010;
    rom[47290] = 25'b1111111011001101110111110;
    rom[47291] = 25'b1111111011001101101100001;
    rom[47292] = 25'b1111111011001101100000100;
    rom[47293] = 25'b1111111011001101010101001;
    rom[47294] = 25'b1111111011001101001001101;
    rom[47295] = 25'b1111111011001100111110010;
    rom[47296] = 25'b1111111011001100110010110;
    rom[47297] = 25'b1111111011001100100111011;
    rom[47298] = 25'b1111111011001100011100001;
    rom[47299] = 25'b1111111011001100010000110;
    rom[47300] = 25'b1111111011001100000101100;
    rom[47301] = 25'b1111111011001011111010010;
    rom[47302] = 25'b1111111011001011101111001;
    rom[47303] = 25'b1111111011001011100011111;
    rom[47304] = 25'b1111111011001011011000110;
    rom[47305] = 25'b1111111011001011001101101;
    rom[47306] = 25'b1111111011001011000010100;
    rom[47307] = 25'b1111111011001010110111100;
    rom[47308] = 25'b1111111011001010101100100;
    rom[47309] = 25'b1111111011001010100001101;
    rom[47310] = 25'b1111111011001010010110100;
    rom[47311] = 25'b1111111011001010001011110;
    rom[47312] = 25'b1111111011001010000000110;
    rom[47313] = 25'b1111111011001001110110000;
    rom[47314] = 25'b1111111011001001101011001;
    rom[47315] = 25'b1111111011001001100000011;
    rom[47316] = 25'b1111111011001001010101101;
    rom[47317] = 25'b1111111011001001001010111;
    rom[47318] = 25'b1111111011001001000000010;
    rom[47319] = 25'b1111111011001000110101101;
    rom[47320] = 25'b1111111011001000101011001;
    rom[47321] = 25'b1111111011001000100000011;
    rom[47322] = 25'b1111111011001000010101111;
    rom[47323] = 25'b1111111011001000001011011;
    rom[47324] = 25'b1111111011001000000001000;
    rom[47325] = 25'b1111111011000111110110100;
    rom[47326] = 25'b1111111011000111101100000;
    rom[47327] = 25'b1111111011000111100001101;
    rom[47328] = 25'b1111111011000111010111010;
    rom[47329] = 25'b1111111011000111001101000;
    rom[47330] = 25'b1111111011000111000010110;
    rom[47331] = 25'b1111111011000110111000100;
    rom[47332] = 25'b1111111011000110101110010;
    rom[47333] = 25'b1111111011000110100100001;
    rom[47334] = 25'b1111111011000110011010000;
    rom[47335] = 25'b1111111011000110001111111;
    rom[47336] = 25'b1111111011000110000101110;
    rom[47337] = 25'b1111111011000101111011110;
    rom[47338] = 25'b1111111011000101110001110;
    rom[47339] = 25'b1111111011000101100111110;
    rom[47340] = 25'b1111111011000101011101110;
    rom[47341] = 25'b1111111011000101010011111;
    rom[47342] = 25'b1111111011000101001010000;
    rom[47343] = 25'b1111111011000101000000001;
    rom[47344] = 25'b1111111011000100110110010;
    rom[47345] = 25'b1111111011000100101100100;
    rom[47346] = 25'b1111111011000100100010110;
    rom[47347] = 25'b1111111011000100011001001;
    rom[47348] = 25'b1111111011000100001111011;
    rom[47349] = 25'b1111111011000100000101110;
    rom[47350] = 25'b1111111011000011111100001;
    rom[47351] = 25'b1111111011000011110010100;
    rom[47352] = 25'b1111111011000011101001000;
    rom[47353] = 25'b1111111011000011011111100;
    rom[47354] = 25'b1111111011000011010101111;
    rom[47355] = 25'b1111111011000011001100100;
    rom[47356] = 25'b1111111011000011000011001;
    rom[47357] = 25'b1111111011000010111001110;
    rom[47358] = 25'b1111111011000010110000011;
    rom[47359] = 25'b1111111011000010100111000;
    rom[47360] = 25'b1111111011000010011101110;
    rom[47361] = 25'b1111111011000010010100100;
    rom[47362] = 25'b1111111011000010001011010;
    rom[47363] = 25'b1111111011000010000010001;
    rom[47364] = 25'b1111111011000001111000111;
    rom[47365] = 25'b1111111011000001101111110;
    rom[47366] = 25'b1111111011000001100110110;
    rom[47367] = 25'b1111111011000001011101101;
    rom[47368] = 25'b1111111011000001010100101;
    rom[47369] = 25'b1111111011000001001011101;
    rom[47370] = 25'b1111111011000001000010101;
    rom[47371] = 25'b1111111011000000111001110;
    rom[47372] = 25'b1111111011000000110000111;
    rom[47373] = 25'b1111111011000000101000000;
    rom[47374] = 25'b1111111011000000011111001;
    rom[47375] = 25'b1111111011000000010110011;
    rom[47376] = 25'b1111111011000000001101101;
    rom[47377] = 25'b1111111011000000000100111;
    rom[47378] = 25'b1111111010111111111100001;
    rom[47379] = 25'b1111111010111111110011100;
    rom[47380] = 25'b1111111010111111101010111;
    rom[47381] = 25'b1111111010111111100010010;
    rom[47382] = 25'b1111111010111111011001110;
    rom[47383] = 25'b1111111010111111010001010;
    rom[47384] = 25'b1111111010111111001000110;
    rom[47385] = 25'b1111111010111111000000010;
    rom[47386] = 25'b1111111010111110110111110;
    rom[47387] = 25'b1111111010111110101111011;
    rom[47388] = 25'b1111111010111110100111000;
    rom[47389] = 25'b1111111010111110011110101;
    rom[47390] = 25'b1111111010111110010110011;
    rom[47391] = 25'b1111111010111110001110000;
    rom[47392] = 25'b1111111010111110000101111;
    rom[47393] = 25'b1111111010111101111101101;
    rom[47394] = 25'b1111111010111101110101100;
    rom[47395] = 25'b1111111010111101101101011;
    rom[47396] = 25'b1111111010111101100101010;
    rom[47397] = 25'b1111111010111101011101001;
    rom[47398] = 25'b1111111010111101010101001;
    rom[47399] = 25'b1111111010111101001101000;
    rom[47400] = 25'b1111111010111101000101001;
    rom[47401] = 25'b1111111010111100111101001;
    rom[47402] = 25'b1111111010111100110101010;
    rom[47403] = 25'b1111111010111100101101011;
    rom[47404] = 25'b1111111010111100100101100;
    rom[47405] = 25'b1111111010111100011101110;
    rom[47406] = 25'b1111111010111100010110000;
    rom[47407] = 25'b1111111010111100001110010;
    rom[47408] = 25'b1111111010111100000110100;
    rom[47409] = 25'b1111111010111011111110110;
    rom[47410] = 25'b1111111010111011110111001;
    rom[47411] = 25'b1111111010111011101111101;
    rom[47412] = 25'b1111111010111011101000000;
    rom[47413] = 25'b1111111010111011100000100;
    rom[47414] = 25'b1111111010111011011000111;
    rom[47415] = 25'b1111111010111011010001011;
    rom[47416] = 25'b1111111010111011001001111;
    rom[47417] = 25'b1111111010111011000010100;
    rom[47418] = 25'b1111111010111010111011001;
    rom[47419] = 25'b1111111010111010110011110;
    rom[47420] = 25'b1111111010111010101100100;
    rom[47421] = 25'b1111111010111010100101001;
    rom[47422] = 25'b1111111010111010011110000;
    rom[47423] = 25'b1111111010111010010110101;
    rom[47424] = 25'b1111111010111010001111100;
    rom[47425] = 25'b1111111010111010001000011;
    rom[47426] = 25'b1111111010111010000001001;
    rom[47427] = 25'b1111111010111001111010001;
    rom[47428] = 25'b1111111010111001110011001;
    rom[47429] = 25'b1111111010111001101100001;
    rom[47430] = 25'b1111111010111001100101001;
    rom[47431] = 25'b1111111010111001011110001;
    rom[47432] = 25'b1111111010111001010111001;
    rom[47433] = 25'b1111111010111001010000010;
    rom[47434] = 25'b1111111010111001001001011;
    rom[47435] = 25'b1111111010111001000010100;
    rom[47436] = 25'b1111111010111000111011110;
    rom[47437] = 25'b1111111010111000110101000;
    rom[47438] = 25'b1111111010111000101110010;
    rom[47439] = 25'b1111111010111000100111100;
    rom[47440] = 25'b1111111010111000100000111;
    rom[47441] = 25'b1111111010111000011010010;
    rom[47442] = 25'b1111111010111000010011101;
    rom[47443] = 25'b1111111010111000001101000;
    rom[47444] = 25'b1111111010111000000110100;
    rom[47445] = 25'b1111111010111000000000000;
    rom[47446] = 25'b1111111010110111111001100;
    rom[47447] = 25'b1111111010110111110011000;
    rom[47448] = 25'b1111111010110111101100110;
    rom[47449] = 25'b1111111010110111100110010;
    rom[47450] = 25'b1111111010110111011111111;
    rom[47451] = 25'b1111111010110111011001101;
    rom[47452] = 25'b1111111010110111010011011;
    rom[47453] = 25'b1111111010110111001101001;
    rom[47454] = 25'b1111111010110111000110111;
    rom[47455] = 25'b1111111010110111000000110;
    rom[47456] = 25'b1111111010110110111010100;
    rom[47457] = 25'b1111111010110110110100011;
    rom[47458] = 25'b1111111010110110101110011;
    rom[47459] = 25'b1111111010110110101000010;
    rom[47460] = 25'b1111111010110110100010010;
    rom[47461] = 25'b1111111010110110011100010;
    rom[47462] = 25'b1111111010110110010110011;
    rom[47463] = 25'b1111111010110110010000011;
    rom[47464] = 25'b1111111010110110001010100;
    rom[47465] = 25'b1111111010110110000100101;
    rom[47466] = 25'b1111111010110101111110110;
    rom[47467] = 25'b1111111010110101111001000;
    rom[47468] = 25'b1111111010110101110011010;
    rom[47469] = 25'b1111111010110101101101100;
    rom[47470] = 25'b1111111010110101100111110;
    rom[47471] = 25'b1111111010110101100010001;
    rom[47472] = 25'b1111111010110101011100100;
    rom[47473] = 25'b1111111010110101010110111;
    rom[47474] = 25'b1111111010110101010001010;
    rom[47475] = 25'b1111111010110101001011110;
    rom[47476] = 25'b1111111010110101000110010;
    rom[47477] = 25'b1111111010110101000000111;
    rom[47478] = 25'b1111111010110100111011011;
    rom[47479] = 25'b1111111010110100110110000;
    rom[47480] = 25'b1111111010110100110000101;
    rom[47481] = 25'b1111111010110100101011010;
    rom[47482] = 25'b1111111010110100100110000;
    rom[47483] = 25'b1111111010110100100000101;
    rom[47484] = 25'b1111111010110100011011011;
    rom[47485] = 25'b1111111010110100010110010;
    rom[47486] = 25'b1111111010110100010001000;
    rom[47487] = 25'b1111111010110100001011111;
    rom[47488] = 25'b1111111010110100000110101;
    rom[47489] = 25'b1111111010110100000001101;
    rom[47490] = 25'b1111111010110011111100101;
    rom[47491] = 25'b1111111010110011110111100;
    rom[47492] = 25'b1111111010110011110010101;
    rom[47493] = 25'b1111111010110011101101101;
    rom[47494] = 25'b1111111010110011101000110;
    rom[47495] = 25'b1111111010110011100011110;
    rom[47496] = 25'b1111111010110011011110111;
    rom[47497] = 25'b1111111010110011011010000;
    rom[47498] = 25'b1111111010110011010101010;
    rom[47499] = 25'b1111111010110011010000100;
    rom[47500] = 25'b1111111010110011001011110;
    rom[47501] = 25'b1111111010110011000111001;
    rom[47502] = 25'b1111111010110011000010011;
    rom[47503] = 25'b1111111010110010111101110;
    rom[47504] = 25'b1111111010110010111001001;
    rom[47505] = 25'b1111111010110010110100101;
    rom[47506] = 25'b1111111010110010110000000;
    rom[47507] = 25'b1111111010110010101011100;
    rom[47508] = 25'b1111111010110010100111000;
    rom[47509] = 25'b1111111010110010100010101;
    rom[47510] = 25'b1111111010110010011110001;
    rom[47511] = 25'b1111111010110010011001110;
    rom[47512] = 25'b1111111010110010010101011;
    rom[47513] = 25'b1111111010110010010001001;
    rom[47514] = 25'b1111111010110010001100111;
    rom[47515] = 25'b1111111010110010001000101;
    rom[47516] = 25'b1111111010110010000100011;
    rom[47517] = 25'b1111111010110010000000010;
    rom[47518] = 25'b1111111010110001111100000;
    rom[47519] = 25'b1111111010110001110111111;
    rom[47520] = 25'b1111111010110001110011110;
    rom[47521] = 25'b1111111010110001101111101;
    rom[47522] = 25'b1111111010110001101011101;
    rom[47523] = 25'b1111111010110001100111101;
    rom[47524] = 25'b1111111010110001100011110;
    rom[47525] = 25'b1111111010110001011111110;
    rom[47526] = 25'b1111111010110001011011111;
    rom[47527] = 25'b1111111010110001011000000;
    rom[47528] = 25'b1111111010110001010100001;
    rom[47529] = 25'b1111111010110001010000010;
    rom[47530] = 25'b1111111010110001001100101;
    rom[47531] = 25'b1111111010110001001000111;
    rom[47532] = 25'b1111111010110001000101001;
    rom[47533] = 25'b1111111010110001000001011;
    rom[47534] = 25'b1111111010110000111101110;
    rom[47535] = 25'b1111111010110000111010001;
    rom[47536] = 25'b1111111010110000110110100;
    rom[47537] = 25'b1111111010110000110011000;
    rom[47538] = 25'b1111111010110000101111011;
    rom[47539] = 25'b1111111010110000101100000;
    rom[47540] = 25'b1111111010110000101000011;
    rom[47541] = 25'b1111111010110000100101001;
    rom[47542] = 25'b1111111010110000100001101;
    rom[47543] = 25'b1111111010110000011110010;
    rom[47544] = 25'b1111111010110000011010111;
    rom[47545] = 25'b1111111010110000010111101;
    rom[47546] = 25'b1111111010110000010100011;
    rom[47547] = 25'b1111111010110000010001001;
    rom[47548] = 25'b1111111010110000001101111;
    rom[47549] = 25'b1111111010110000001010110;
    rom[47550] = 25'b1111111010110000000111100;
    rom[47551] = 25'b1111111010110000000100100;
    rom[47552] = 25'b1111111010110000000001011;
    rom[47553] = 25'b1111111010101111111110010;
    rom[47554] = 25'b1111111010101111111011010;
    rom[47555] = 25'b1111111010101111111000010;
    rom[47556] = 25'b1111111010101111110101011;
    rom[47557] = 25'b1111111010101111110010011;
    rom[47558] = 25'b1111111010101111101111100;
    rom[47559] = 25'b1111111010101111101100101;
    rom[47560] = 25'b1111111010101111101001110;
    rom[47561] = 25'b1111111010101111100111000;
    rom[47562] = 25'b1111111010101111100100010;
    rom[47563] = 25'b1111111010101111100001100;
    rom[47564] = 25'b1111111010101111011110110;
    rom[47565] = 25'b1111111010101111011100000;
    rom[47566] = 25'b1111111010101111011001011;
    rom[47567] = 25'b1111111010101111010110110;
    rom[47568] = 25'b1111111010101111010100010;
    rom[47569] = 25'b1111111010101111010001101;
    rom[47570] = 25'b1111111010101111001111001;
    rom[47571] = 25'b1111111010101111001100101;
    rom[47572] = 25'b1111111010101111001010010;
    rom[47573] = 25'b1111111010101111000111110;
    rom[47574] = 25'b1111111010101111000101011;
    rom[47575] = 25'b1111111010101111000011000;
    rom[47576] = 25'b1111111010101111000000101;
    rom[47577] = 25'b1111111010101110111110011;
    rom[47578] = 25'b1111111010101110111100001;
    rom[47579] = 25'b1111111010101110111001111;
    rom[47580] = 25'b1111111010101110110111101;
    rom[47581] = 25'b1111111010101110110101100;
    rom[47582] = 25'b1111111010101110110011011;
    rom[47583] = 25'b1111111010101110110001001;
    rom[47584] = 25'b1111111010101110101111001;
    rom[47585] = 25'b1111111010101110101101000;
    rom[47586] = 25'b1111111010101110101011000;
    rom[47587] = 25'b1111111010101110101001000;
    rom[47588] = 25'b1111111010101110100111001;
    rom[47589] = 25'b1111111010101110100101001;
    rom[47590] = 25'b1111111010101110100011010;
    rom[47591] = 25'b1111111010101110100001011;
    rom[47592] = 25'b1111111010101110011111100;
    rom[47593] = 25'b1111111010101110011101110;
    rom[47594] = 25'b1111111010101110011100000;
    rom[47595] = 25'b1111111010101110011010010;
    rom[47596] = 25'b1111111010101110011000011;
    rom[47597] = 25'b1111111010101110010110110;
    rom[47598] = 25'b1111111010101110010101001;
    rom[47599] = 25'b1111111010101110010011100;
    rom[47600] = 25'b1111111010101110010001111;
    rom[47601] = 25'b1111111010101110010000011;
    rom[47602] = 25'b1111111010101110001110110;
    rom[47603] = 25'b1111111010101110001101010;
    rom[47604] = 25'b1111111010101110001011111;
    rom[47605] = 25'b1111111010101110001010011;
    rom[47606] = 25'b1111111010101110001001000;
    rom[47607] = 25'b1111111010101110000111101;
    rom[47608] = 25'b1111111010101110000110010;
    rom[47609] = 25'b1111111010101110000101000;
    rom[47610] = 25'b1111111010101110000011110;
    rom[47611] = 25'b1111111010101110000010011;
    rom[47612] = 25'b1111111010101110000001001;
    rom[47613] = 25'b1111111010101110000000000;
    rom[47614] = 25'b1111111010101101111110111;
    rom[47615] = 25'b1111111010101101111101110;
    rom[47616] = 25'b1111111010101101111100101;
    rom[47617] = 25'b1111111010101101111011101;
    rom[47618] = 25'b1111111010101101111010100;
    rom[47619] = 25'b1111111010101101111001100;
    rom[47620] = 25'b1111111010101101111000100;
    rom[47621] = 25'b1111111010101101110111100;
    rom[47622] = 25'b1111111010101101110110101;
    rom[47623] = 25'b1111111010101101110101110;
    rom[47624] = 25'b1111111010101101110100111;
    rom[47625] = 25'b1111111010101101110100001;
    rom[47626] = 25'b1111111010101101110011010;
    rom[47627] = 25'b1111111010101101110010100;
    rom[47628] = 25'b1111111010101101110001110;
    rom[47629] = 25'b1111111010101101110001001;
    rom[47630] = 25'b1111111010101101110000011;
    rom[47631] = 25'b1111111010101101101111110;
    rom[47632] = 25'b1111111010101101101111001;
    rom[47633] = 25'b1111111010101101101110101;
    rom[47634] = 25'b1111111010101101101110000;
    rom[47635] = 25'b1111111010101101101101100;
    rom[47636] = 25'b1111111010101101101101000;
    rom[47637] = 25'b1111111010101101101100100;
    rom[47638] = 25'b1111111010101101101100001;
    rom[47639] = 25'b1111111010101101101011110;
    rom[47640] = 25'b1111111010101101101011011;
    rom[47641] = 25'b1111111010101101101011000;
    rom[47642] = 25'b1111111010101101101010101;
    rom[47643] = 25'b1111111010101101101010011;
    rom[47644] = 25'b1111111010101101101010010;
    rom[47645] = 25'b1111111010101101101001111;
    rom[47646] = 25'b1111111010101101101001110;
    rom[47647] = 25'b1111111010101101101001100;
    rom[47648] = 25'b1111111010101101101001100;
    rom[47649] = 25'b1111111010101101101001011;
    rom[47650] = 25'b1111111010101101101001010;
    rom[47651] = 25'b1111111010101101101001010;
    rom[47652] = 25'b1111111010101101101001010;
    rom[47653] = 25'b1111111010101101101001010;
    rom[47654] = 25'b1111111010101101101001010;
    rom[47655] = 25'b1111111010101101101001011;
    rom[47656] = 25'b1111111010101101101001100;
    rom[47657] = 25'b1111111010101101101001101;
    rom[47658] = 25'b1111111010101101101001111;
    rom[47659] = 25'b1111111010101101101010000;
    rom[47660] = 25'b1111111010101101101010010;
    rom[47661] = 25'b1111111010101101101010100;
    rom[47662] = 25'b1111111010101101101010110;
    rom[47663] = 25'b1111111010101101101011001;
    rom[47664] = 25'b1111111010101101101011100;
    rom[47665] = 25'b1111111010101101101011111;
    rom[47666] = 25'b1111111010101101101100010;
    rom[47667] = 25'b1111111010101101101100110;
    rom[47668] = 25'b1111111010101101101101001;
    rom[47669] = 25'b1111111010101101101101101;
    rom[47670] = 25'b1111111010101101101110010;
    rom[47671] = 25'b1111111010101101101110110;
    rom[47672] = 25'b1111111010101101101111011;
    rom[47673] = 25'b1111111010101101110000000;
    rom[47674] = 25'b1111111010101101110000101;
    rom[47675] = 25'b1111111010101101110001010;
    rom[47676] = 25'b1111111010101101110010000;
    rom[47677] = 25'b1111111010101101110010110;
    rom[47678] = 25'b1111111010101101110011100;
    rom[47679] = 25'b1111111010101101110100010;
    rom[47680] = 25'b1111111010101101110101001;
    rom[47681] = 25'b1111111010101101110110000;
    rom[47682] = 25'b1111111010101101110110111;
    rom[47683] = 25'b1111111010101101110111111;
    rom[47684] = 25'b1111111010101101111000110;
    rom[47685] = 25'b1111111010101101111001110;
    rom[47686] = 25'b1111111010101101111010110;
    rom[47687] = 25'b1111111010101101111011110;
    rom[47688] = 25'b1111111010101101111100110;
    rom[47689] = 25'b1111111010101101111101111;
    rom[47690] = 25'b1111111010101101111111000;
    rom[47691] = 25'b1111111010101110000000001;
    rom[47692] = 25'b1111111010101110000001011;
    rom[47693] = 25'b1111111010101110000010101;
    rom[47694] = 25'b1111111010101110000011110;
    rom[47695] = 25'b1111111010101110000101001;
    rom[47696] = 25'b1111111010101110000110011;
    rom[47697] = 25'b1111111010101110000111110;
    rom[47698] = 25'b1111111010101110001001001;
    rom[47699] = 25'b1111111010101110001010011;
    rom[47700] = 25'b1111111010101110001011111;
    rom[47701] = 25'b1111111010101110001101010;
    rom[47702] = 25'b1111111010101110001110110;
    rom[47703] = 25'b1111111010101110010000010;
    rom[47704] = 25'b1111111010101110010001110;
    rom[47705] = 25'b1111111010101110010011011;
    rom[47706] = 25'b1111111010101110010101000;
    rom[47707] = 25'b1111111010101110010110100;
    rom[47708] = 25'b1111111010101110011000010;
    rom[47709] = 25'b1111111010101110011001111;
    rom[47710] = 25'b1111111010101110011011101;
    rom[47711] = 25'b1111111010101110011101011;
    rom[47712] = 25'b1111111010101110011111001;
    rom[47713] = 25'b1111111010101110100000111;
    rom[47714] = 25'b1111111010101110100010110;
    rom[47715] = 25'b1111111010101110100100101;
    rom[47716] = 25'b1111111010101110100110100;
    rom[47717] = 25'b1111111010101110101000011;
    rom[47718] = 25'b1111111010101110101010011;
    rom[47719] = 25'b1111111010101110101100011;
    rom[47720] = 25'b1111111010101110101110010;
    rom[47721] = 25'b1111111010101110110000011;
    rom[47722] = 25'b1111111010101110110010011;
    rom[47723] = 25'b1111111010101110110100100;
    rom[47724] = 25'b1111111010101110110110101;
    rom[47725] = 25'b1111111010101110111000110;
    rom[47726] = 25'b1111111010101110111010111;
    rom[47727] = 25'b1111111010101110111101001;
    rom[47728] = 25'b1111111010101110111111011;
    rom[47729] = 25'b1111111010101111000001101;
    rom[47730] = 25'b1111111010101111000011111;
    rom[47731] = 25'b1111111010101111000110001;
    rom[47732] = 25'b1111111010101111001000100;
    rom[47733] = 25'b1111111010101111001011000;
    rom[47734] = 25'b1111111010101111001101010;
    rom[47735] = 25'b1111111010101111001111110;
    rom[47736] = 25'b1111111010101111010010010;
    rom[47737] = 25'b1111111010101111010100101;
    rom[47738] = 25'b1111111010101111010111001;
    rom[47739] = 25'b1111111010101111011001110;
    rom[47740] = 25'b1111111010101111011100011;
    rom[47741] = 25'b1111111010101111011110111;
    rom[47742] = 25'b1111111010101111100001100;
    rom[47743] = 25'b1111111010101111100100010;
    rom[47744] = 25'b1111111010101111100110111;
    rom[47745] = 25'b1111111010101111101001101;
    rom[47746] = 25'b1111111010101111101100011;
    rom[47747] = 25'b1111111010101111101111001;
    rom[47748] = 25'b1111111010101111110010000;
    rom[47749] = 25'b1111111010101111110100110;
    rom[47750] = 25'b1111111010101111110111101;
    rom[47751] = 25'b1111111010101111111010100;
    rom[47752] = 25'b1111111010101111111101100;
    rom[47753] = 25'b1111111010110000000000011;
    rom[47754] = 25'b1111111010110000000011011;
    rom[47755] = 25'b1111111010110000000110011;
    rom[47756] = 25'b1111111010110000001001011;
    rom[47757] = 25'b1111111010110000001100011;
    rom[47758] = 25'b1111111010110000001111100;
    rom[47759] = 25'b1111111010110000010010101;
    rom[47760] = 25'b1111111010110000010101110;
    rom[47761] = 25'b1111111010110000011000111;
    rom[47762] = 25'b1111111010110000011100001;
    rom[47763] = 25'b1111111010110000011111011;
    rom[47764] = 25'b1111111010110000100010101;
    rom[47765] = 25'b1111111010110000100101111;
    rom[47766] = 25'b1111111010110000101001001;
    rom[47767] = 25'b1111111010110000101100100;
    rom[47768] = 25'b1111111010110000101111111;
    rom[47769] = 25'b1111111010110000110011011;
    rom[47770] = 25'b1111111010110000110110110;
    rom[47771] = 25'b1111111010110000111010001;
    rom[47772] = 25'b1111111010110000111101101;
    rom[47773] = 25'b1111111010110001000001001;
    rom[47774] = 25'b1111111010110001000100110;
    rom[47775] = 25'b1111111010110001001000010;
    rom[47776] = 25'b1111111010110001001011111;
    rom[47777] = 25'b1111111010110001001111100;
    rom[47778] = 25'b1111111010110001010011001;
    rom[47779] = 25'b1111111010110001010110111;
    rom[47780] = 25'b1111111010110001011010100;
    rom[47781] = 25'b1111111010110001011110010;
    rom[47782] = 25'b1111111010110001100010000;
    rom[47783] = 25'b1111111010110001100101110;
    rom[47784] = 25'b1111111010110001101001101;
    rom[47785] = 25'b1111111010110001101101100;
    rom[47786] = 25'b1111111010110001110001010;
    rom[47787] = 25'b1111111010110001110101010;
    rom[47788] = 25'b1111111010110001111001001;
    rom[47789] = 25'b1111111010110001111101000;
    rom[47790] = 25'b1111111010110010000001000;
    rom[47791] = 25'b1111111010110010000101001;
    rom[47792] = 25'b1111111010110010001001001;
    rom[47793] = 25'b1111111010110010001101001;
    rom[47794] = 25'b1111111010110010010001010;
    rom[47795] = 25'b1111111010110010010101011;
    rom[47796] = 25'b1111111010110010011001100;
    rom[47797] = 25'b1111111010110010011101101;
    rom[47798] = 25'b1111111010110010100001111;
    rom[47799] = 25'b1111111010110010100110001;
    rom[47800] = 25'b1111111010110010101010011;
    rom[47801] = 25'b1111111010110010101110101;
    rom[47802] = 25'b1111111010110010110010111;
    rom[47803] = 25'b1111111010110010110111010;
    rom[47804] = 25'b1111111010110010111011101;
    rom[47805] = 25'b1111111010110011000000000;
    rom[47806] = 25'b1111111010110011000100100;
    rom[47807] = 25'b1111111010110011001000111;
    rom[47808] = 25'b1111111010110011001101011;
    rom[47809] = 25'b1111111010110011010001111;
    rom[47810] = 25'b1111111010110011010110011;
    rom[47811] = 25'b1111111010110011011011000;
    rom[47812] = 25'b1111111010110011011111100;
    rom[47813] = 25'b1111111010110011100100001;
    rom[47814] = 25'b1111111010110011101000110;
    rom[47815] = 25'b1111111010110011101101100;
    rom[47816] = 25'b1111111010110011110010001;
    rom[47817] = 25'b1111111010110011110110110;
    rom[47818] = 25'b1111111010110011111011101;
    rom[47819] = 25'b1111111010110100000000011;
    rom[47820] = 25'b1111111010110100000101010;
    rom[47821] = 25'b1111111010110100001010000;
    rom[47822] = 25'b1111111010110100001110110;
    rom[47823] = 25'b1111111010110100010011110;
    rom[47824] = 25'b1111111010110100011000101;
    rom[47825] = 25'b1111111010110100011101101;
    rom[47826] = 25'b1111111010110100100010100;
    rom[47827] = 25'b1111111010110100100111100;
    rom[47828] = 25'b1111111010110100101100100;
    rom[47829] = 25'b1111111010110100110001100;
    rom[47830] = 25'b1111111010110100110110101;
    rom[47831] = 25'b1111111010110100111011110;
    rom[47832] = 25'b1111111010110101000000111;
    rom[47833] = 25'b1111111010110101000110000;
    rom[47834] = 25'b1111111010110101001011001;
    rom[47835] = 25'b1111111010110101010000011;
    rom[47836] = 25'b1111111010110101010101101;
    rom[47837] = 25'b1111111010110101011010111;
    rom[47838] = 25'b1111111010110101100000001;
    rom[47839] = 25'b1111111010110101100101100;
    rom[47840] = 25'b1111111010110101101010110;
    rom[47841] = 25'b1111111010110101110000001;
    rom[47842] = 25'b1111111010110101110101100;
    rom[47843] = 25'b1111111010110101111011000;
    rom[47844] = 25'b1111111010110110000000011;
    rom[47845] = 25'b1111111010110110000101111;
    rom[47846] = 25'b1111111010110110001011011;
    rom[47847] = 25'b1111111010110110010000111;
    rom[47848] = 25'b1111111010110110010110011;
    rom[47849] = 25'b1111111010110110011100000;
    rom[47850] = 25'b1111111010110110100001101;
    rom[47851] = 25'b1111111010110110100111010;
    rom[47852] = 25'b1111111010110110101100111;
    rom[47853] = 25'b1111111010110110110010100;
    rom[47854] = 25'b1111111010110110111000010;
    rom[47855] = 25'b1111111010110110111110000;
    rom[47856] = 25'b1111111010110111000011110;
    rom[47857] = 25'b1111111010110111001001100;
    rom[47858] = 25'b1111111010110111001111011;
    rom[47859] = 25'b1111111010110111010101001;
    rom[47860] = 25'b1111111010110111011011000;
    rom[47861] = 25'b1111111010110111100000111;
    rom[47862] = 25'b1111111010110111100110111;
    rom[47863] = 25'b1111111010110111101100110;
    rom[47864] = 25'b1111111010110111110010110;
    rom[47865] = 25'b1111111010110111111000110;
    rom[47866] = 25'b1111111010110111111110111;
    rom[47867] = 25'b1111111010111000000100110;
    rom[47868] = 25'b1111111010111000001010111;
    rom[47869] = 25'b1111111010111000010001000;
    rom[47870] = 25'b1111111010111000010111001;
    rom[47871] = 25'b1111111010111000011101010;
    rom[47872] = 25'b1111111010111000100011011;
    rom[47873] = 25'b1111111010111000101001101;
    rom[47874] = 25'b1111111010111000101111111;
    rom[47875] = 25'b1111111010111000110110001;
    rom[47876] = 25'b1111111010111000111100011;
    rom[47877] = 25'b1111111010111001000010110;
    rom[47878] = 25'b1111111010111001001001000;
    rom[47879] = 25'b1111111010111001001111011;
    rom[47880] = 25'b1111111010111001010101110;
    rom[47881] = 25'b1111111010111001011100010;
    rom[47882] = 25'b1111111010111001100010101;
    rom[47883] = 25'b1111111010111001101001001;
    rom[47884] = 25'b1111111010111001101111100;
    rom[47885] = 25'b1111111010111001110110001;
    rom[47886] = 25'b1111111010111001111100101;
    rom[47887] = 25'b1111111010111010000011001;
    rom[47888] = 25'b1111111010111010001001110;
    rom[47889] = 25'b1111111010111010010000011;
    rom[47890] = 25'b1111111010111010010111000;
    rom[47891] = 25'b1111111010111010011101101;
    rom[47892] = 25'b1111111010111010100100011;
    rom[47893] = 25'b1111111010111010101011001;
    rom[47894] = 25'b1111111010111010110001111;
    rom[47895] = 25'b1111111010111010111000101;
    rom[47896] = 25'b1111111010111010111111011;
    rom[47897] = 25'b1111111010111011000110010;
    rom[47898] = 25'b1111111010111011001101000;
    rom[47899] = 25'b1111111010111011010011111;
    rom[47900] = 25'b1111111010111011011010110;
    rom[47901] = 25'b1111111010111011100001110;
    rom[47902] = 25'b1111111010111011101000101;
    rom[47903] = 25'b1111111010111011101111101;
    rom[47904] = 25'b1111111010111011110110101;
    rom[47905] = 25'b1111111010111011111101101;
    rom[47906] = 25'b1111111010111100000100101;
    rom[47907] = 25'b1111111010111100001011110;
    rom[47908] = 25'b1111111010111100010010111;
    rom[47909] = 25'b1111111010111100011010000;
    rom[47910] = 25'b1111111010111100100001001;
    rom[47911] = 25'b1111111010111100101000010;
    rom[47912] = 25'b1111111010111100101111100;
    rom[47913] = 25'b1111111010111100110110101;
    rom[47914] = 25'b1111111010111100111101111;
    rom[47915] = 25'b1111111010111101000101010;
    rom[47916] = 25'b1111111010111101001100100;
    rom[47917] = 25'b1111111010111101010011110;
    rom[47918] = 25'b1111111010111101011011001;
    rom[47919] = 25'b1111111010111101100010100;
    rom[47920] = 25'b1111111010111101101001111;
    rom[47921] = 25'b1111111010111101110001010;
    rom[47922] = 25'b1111111010111101111000110;
    rom[47923] = 25'b1111111010111110000000010;
    rom[47924] = 25'b1111111010111110000111110;
    rom[47925] = 25'b1111111010111110001111010;
    rom[47926] = 25'b1111111010111110010110111;
    rom[47927] = 25'b1111111010111110011110011;
    rom[47928] = 25'b1111111010111110100110000;
    rom[47929] = 25'b1111111010111110101101100;
    rom[47930] = 25'b1111111010111110110101001;
    rom[47931] = 25'b1111111010111110111100111;
    rom[47932] = 25'b1111111010111111000100101;
    rom[47933] = 25'b1111111010111111001100010;
    rom[47934] = 25'b1111111010111111010100000;
    rom[47935] = 25'b1111111010111111011011110;
    rom[47936] = 25'b1111111010111111100011101;
    rom[47937] = 25'b1111111010111111101011011;
    rom[47938] = 25'b1111111010111111110011001;
    rom[47939] = 25'b1111111010111111111011000;
    rom[47940] = 25'b1111111011000000000011000;
    rom[47941] = 25'b1111111011000000001010111;
    rom[47942] = 25'b1111111011000000010010110;
    rom[47943] = 25'b1111111011000000011010110;
    rom[47944] = 25'b1111111011000000100010110;
    rom[47945] = 25'b1111111011000000101010110;
    rom[47946] = 25'b1111111011000000110010110;
    rom[47947] = 25'b1111111011000000111010110;
    rom[47948] = 25'b1111111011000001000010111;
    rom[47949] = 25'b1111111011000001001011000;
    rom[47950] = 25'b1111111011000001010011001;
    rom[47951] = 25'b1111111011000001011011010;
    rom[47952] = 25'b1111111011000001100011011;
    rom[47953] = 25'b1111111011000001101011101;
    rom[47954] = 25'b1111111011000001110011111;
    rom[47955] = 25'b1111111011000001111100001;
    rom[47956] = 25'b1111111011000010000100011;
    rom[47957] = 25'b1111111011000010001100110;
    rom[47958] = 25'b1111111011000010010101000;
    rom[47959] = 25'b1111111011000010011101011;
    rom[47960] = 25'b1111111011000010100101110;
    rom[47961] = 25'b1111111011000010101110001;
    rom[47962] = 25'b1111111011000010110110100;
    rom[47963] = 25'b1111111011000010111111000;
    rom[47964] = 25'b1111111011000011000111100;
    rom[47965] = 25'b1111111011000011010000000;
    rom[47966] = 25'b1111111011000011011000100;
    rom[47967] = 25'b1111111011000011100001000;
    rom[47968] = 25'b1111111011000011101001100;
    rom[47969] = 25'b1111111011000011110010001;
    rom[47970] = 25'b1111111011000011111010110;
    rom[47971] = 25'b1111111011000100000011011;
    rom[47972] = 25'b1111111011000100001100000;
    rom[47973] = 25'b1111111011000100010100101;
    rom[47974] = 25'b1111111011000100011101011;
    rom[47975] = 25'b1111111011000100100110000;
    rom[47976] = 25'b1111111011000100101110111;
    rom[47977] = 25'b1111111011000100110111101;
    rom[47978] = 25'b1111111011000101000000011;
    rom[47979] = 25'b1111111011000101001001010;
    rom[47980] = 25'b1111111011000101010010000;
    rom[47981] = 25'b1111111011000101011010111;
    rom[47982] = 25'b1111111011000101100011110;
    rom[47983] = 25'b1111111011000101101100110;
    rom[47984] = 25'b1111111011000101110101101;
    rom[47985] = 25'b1111111011000101111110101;
    rom[47986] = 25'b1111111011000110000111100;
    rom[47987] = 25'b1111111011000110010000101;
    rom[47988] = 25'b1111111011000110011001101;
    rom[47989] = 25'b1111111011000110100010101;
    rom[47990] = 25'b1111111011000110101011110;
    rom[47991] = 25'b1111111011000110110100111;
    rom[47992] = 25'b1111111011000110111110000;
    rom[47993] = 25'b1111111011000111000111001;
    rom[47994] = 25'b1111111011000111010000010;
    rom[47995] = 25'b1111111011000111011001100;
    rom[47996] = 25'b1111111011000111100010110;
    rom[47997] = 25'b1111111011000111101100000;
    rom[47998] = 25'b1111111011000111110101001;
    rom[47999] = 25'b1111111011000111111110011;
    rom[48000] = 25'b1111111011001000000111110;
    rom[48001] = 25'b1111111011001000010001001;
    rom[48002] = 25'b1111111011001000011010100;
    rom[48003] = 25'b1111111011001000100011110;
    rom[48004] = 25'b1111111011001000101101010;
    rom[48005] = 25'b1111111011001000110110100;
    rom[48006] = 25'b1111111011001001000000001;
    rom[48007] = 25'b1111111011001001001001100;
    rom[48008] = 25'b1111111011001001010011000;
    rom[48009] = 25'b1111111011001001011100100;
    rom[48010] = 25'b1111111011001001100110000;
    rom[48011] = 25'b1111111011001001101111101;
    rom[48012] = 25'b1111111011001001111001001;
    rom[48013] = 25'b1111111011001010000010110;
    rom[48014] = 25'b1111111011001010001100011;
    rom[48015] = 25'b1111111011001010010110000;
    rom[48016] = 25'b1111111011001010011111110;
    rom[48017] = 25'b1111111011001010101001011;
    rom[48018] = 25'b1111111011001010110011000;
    rom[48019] = 25'b1111111011001010111100111;
    rom[48020] = 25'b1111111011001011000110100;
    rom[48021] = 25'b1111111011001011010000011;
    rom[48022] = 25'b1111111011001011011010001;
    rom[48023] = 25'b1111111011001011100100000;
    rom[48024] = 25'b1111111011001011101101110;
    rom[48025] = 25'b1111111011001011110111101;
    rom[48026] = 25'b1111111011001100000001101;
    rom[48027] = 25'b1111111011001100001011100;
    rom[48028] = 25'b1111111011001100010101100;
    rom[48029] = 25'b1111111011001100011111011;
    rom[48030] = 25'b1111111011001100101001011;
    rom[48031] = 25'b1111111011001100110011011;
    rom[48032] = 25'b1111111011001100111101011;
    rom[48033] = 25'b1111111011001101000111011;
    rom[48034] = 25'b1111111011001101010001100;
    rom[48035] = 25'b1111111011001101011011101;
    rom[48036] = 25'b1111111011001101100101110;
    rom[48037] = 25'b1111111011001101101111111;
    rom[48038] = 25'b1111111011001101111010000;
    rom[48039] = 25'b1111111011001110000100001;
    rom[48040] = 25'b1111111011001110001110011;
    rom[48041] = 25'b1111111011001110011000101;
    rom[48042] = 25'b1111111011001110100010111;
    rom[48043] = 25'b1111111011001110101101001;
    rom[48044] = 25'b1111111011001110110111011;
    rom[48045] = 25'b1111111011001111000001101;
    rom[48046] = 25'b1111111011001111001100000;
    rom[48047] = 25'b1111111011001111010110011;
    rom[48048] = 25'b1111111011001111100000110;
    rom[48049] = 25'b1111111011001111101011001;
    rom[48050] = 25'b1111111011001111110101100;
    rom[48051] = 25'b1111111011010000000000000;
    rom[48052] = 25'b1111111011010000001010011;
    rom[48053] = 25'b1111111011010000010100111;
    rom[48054] = 25'b1111111011010000011111100;
    rom[48055] = 25'b1111111011010000101010000;
    rom[48056] = 25'b1111111011010000110100100;
    rom[48057] = 25'b1111111011010000111111001;
    rom[48058] = 25'b1111111011010001001001101;
    rom[48059] = 25'b1111111011010001010100010;
    rom[48060] = 25'b1111111011010001011110111;
    rom[48061] = 25'b1111111011010001101001101;
    rom[48062] = 25'b1111111011010001110100010;
    rom[48063] = 25'b1111111011010001111110111;
    rom[48064] = 25'b1111111011010010001001101;
    rom[48065] = 25'b1111111011010010010100011;
    rom[48066] = 25'b1111111011010010011111001;
    rom[48067] = 25'b1111111011010010101001111;
    rom[48068] = 25'b1111111011010010110100101;
    rom[48069] = 25'b1111111011010010111111100;
    rom[48070] = 25'b1111111011010011001010011;
    rom[48071] = 25'b1111111011010011010101010;
    rom[48072] = 25'b1111111011010011100000001;
    rom[48073] = 25'b1111111011010011101011000;
    rom[48074] = 25'b1111111011010011110110000;
    rom[48075] = 25'b1111111011010100000000111;
    rom[48076] = 25'b1111111011010100001011111;
    rom[48077] = 25'b1111111011010100010110111;
    rom[48078] = 25'b1111111011010100100001111;
    rom[48079] = 25'b1111111011010100101101000;
    rom[48080] = 25'b1111111011010100111000000;
    rom[48081] = 25'b1111111011010101000011001;
    rom[48082] = 25'b1111111011010101001110001;
    rom[48083] = 25'b1111111011010101011001010;
    rom[48084] = 25'b1111111011010101100100011;
    rom[48085] = 25'b1111111011010101101111100;
    rom[48086] = 25'b1111111011010101111010110;
    rom[48087] = 25'b1111111011010110000110000;
    rom[48088] = 25'b1111111011010110010001001;
    rom[48089] = 25'b1111111011010110011100011;
    rom[48090] = 25'b1111111011010110100111101;
    rom[48091] = 25'b1111111011010110110011000;
    rom[48092] = 25'b1111111011010110111110010;
    rom[48093] = 25'b1111111011010111001001101;
    rom[48094] = 25'b1111111011010111010100111;
    rom[48095] = 25'b1111111011010111100000010;
    rom[48096] = 25'b1111111011010111101011101;
    rom[48097] = 25'b1111111011010111110111000;
    rom[48098] = 25'b1111111011011000000010011;
    rom[48099] = 25'b1111111011011000001101111;
    rom[48100] = 25'b1111111011011000011001011;
    rom[48101] = 25'b1111111011011000100100111;
    rom[48102] = 25'b1111111011011000110000011;
    rom[48103] = 25'b1111111011011000111011111;
    rom[48104] = 25'b1111111011011001000111100;
    rom[48105] = 25'b1111111011011001010011000;
    rom[48106] = 25'b1111111011011001011110101;
    rom[48107] = 25'b1111111011011001101010010;
    rom[48108] = 25'b1111111011011001110101111;
    rom[48109] = 25'b1111111011011010000001100;
    rom[48110] = 25'b1111111011011010001101001;
    rom[48111] = 25'b1111111011011010011000110;
    rom[48112] = 25'b1111111011011010100100100;
    rom[48113] = 25'b1111111011011010110000010;
    rom[48114] = 25'b1111111011011010111100000;
    rom[48115] = 25'b1111111011011011000111110;
    rom[48116] = 25'b1111111011011011010011100;
    rom[48117] = 25'b1111111011011011011111011;
    rom[48118] = 25'b1111111011011011101011001;
    rom[48119] = 25'b1111111011011011110111000;
    rom[48120] = 25'b1111111011011100000010111;
    rom[48121] = 25'b1111111011011100001110110;
    rom[48122] = 25'b1111111011011100011010110;
    rom[48123] = 25'b1111111011011100100110101;
    rom[48124] = 25'b1111111011011100110010101;
    rom[48125] = 25'b1111111011011100111110100;
    rom[48126] = 25'b1111111011011101001010100;
    rom[48127] = 25'b1111111011011101010110100;
    rom[48128] = 25'b1111111011011101100010100;
    rom[48129] = 25'b1111111011011101101110100;
    rom[48130] = 25'b1111111011011101111010101;
    rom[48131] = 25'b1111111011011110000110110;
    rom[48132] = 25'b1111111011011110010010110;
    rom[48133] = 25'b1111111011011110011110111;
    rom[48134] = 25'b1111111011011110101011001;
    rom[48135] = 25'b1111111011011110110111010;
    rom[48136] = 25'b1111111011011111000011100;
    rom[48137] = 25'b1111111011011111001111101;
    rom[48138] = 25'b1111111011011111011011111;
    rom[48139] = 25'b1111111011011111101000000;
    rom[48140] = 25'b1111111011011111110100010;
    rom[48141] = 25'b1111111011100000000000101;
    rom[48142] = 25'b1111111011100000001100111;
    rom[48143] = 25'b1111111011100000011001001;
    rom[48144] = 25'b1111111011100000100101100;
    rom[48145] = 25'b1111111011100000110001111;
    rom[48146] = 25'b1111111011100000111110010;
    rom[48147] = 25'b1111111011100001001010101;
    rom[48148] = 25'b1111111011100001010111001;
    rom[48149] = 25'b1111111011100001100011100;
    rom[48150] = 25'b1111111011100001101111111;
    rom[48151] = 25'b1111111011100001111100100;
    rom[48152] = 25'b1111111011100010001000111;
    rom[48153] = 25'b1111111011100010010101011;
    rom[48154] = 25'b1111111011100010100001111;
    rom[48155] = 25'b1111111011100010101110011;
    rom[48156] = 25'b1111111011100010111011000;
    rom[48157] = 25'b1111111011100011000111101;
    rom[48158] = 25'b1111111011100011010100010;
    rom[48159] = 25'b1111111011100011100000111;
    rom[48160] = 25'b1111111011100011101101100;
    rom[48161] = 25'b1111111011100011111010000;
    rom[48162] = 25'b1111111011100100000110110;
    rom[48163] = 25'b1111111011100100010011100;
    rom[48164] = 25'b1111111011100100100000001;
    rom[48165] = 25'b1111111011100100101100111;
    rom[48166] = 25'b1111111011100100111001101;
    rom[48167] = 25'b1111111011100101000110011;
    rom[48168] = 25'b1111111011100101010011010;
    rom[48169] = 25'b1111111011100101100000000;
    rom[48170] = 25'b1111111011100101101100111;
    rom[48171] = 25'b1111111011100101111001101;
    rom[48172] = 25'b1111111011100110000110100;
    rom[48173] = 25'b1111111011100110010011011;
    rom[48174] = 25'b1111111011100110100000010;
    rom[48175] = 25'b1111111011100110101101001;
    rom[48176] = 25'b1111111011100110111010001;
    rom[48177] = 25'b1111111011100111000111000;
    rom[48178] = 25'b1111111011100111010100000;
    rom[48179] = 25'b1111111011100111100001000;
    rom[48180] = 25'b1111111011100111101110000;
    rom[48181] = 25'b1111111011100111111011000;
    rom[48182] = 25'b1111111011101000001000001;
    rom[48183] = 25'b1111111011101000010101001;
    rom[48184] = 25'b1111111011101000100010001;
    rom[48185] = 25'b1111111011101000101111011;
    rom[48186] = 25'b1111111011101000111100011;
    rom[48187] = 25'b1111111011101001001001101;
    rom[48188] = 25'b1111111011101001010110101;
    rom[48189] = 25'b1111111011101001100011111;
    rom[48190] = 25'b1111111011101001110001001;
    rom[48191] = 25'b1111111011101001111110010;
    rom[48192] = 25'b1111111011101010001011011;
    rom[48193] = 25'b1111111011101010011000101;
    rom[48194] = 25'b1111111011101010100110000;
    rom[48195] = 25'b1111111011101010110011010;
    rom[48196] = 25'b1111111011101011000000100;
    rom[48197] = 25'b1111111011101011001101111;
    rom[48198] = 25'b1111111011101011011011001;
    rom[48199] = 25'b1111111011101011101000100;
    rom[48200] = 25'b1111111011101011110101111;
    rom[48201] = 25'b1111111011101100000011010;
    rom[48202] = 25'b1111111011101100010000101;
    rom[48203] = 25'b1111111011101100011110000;
    rom[48204] = 25'b1111111011101100101011100;
    rom[48205] = 25'b1111111011101100111000111;
    rom[48206] = 25'b1111111011101101000110011;
    rom[48207] = 25'b1111111011101101010011111;
    rom[48208] = 25'b1111111011101101100001011;
    rom[48209] = 25'b1111111011101101101110111;
    rom[48210] = 25'b1111111011101101111100100;
    rom[48211] = 25'b1111111011101110001010000;
    rom[48212] = 25'b1111111011101110010111100;
    rom[48213] = 25'b1111111011101110100101001;
    rom[48214] = 25'b1111111011101110110010110;
    rom[48215] = 25'b1111111011101111000000011;
    rom[48216] = 25'b1111111011101111001110000;
    rom[48217] = 25'b1111111011101111011011101;
    rom[48218] = 25'b1111111011101111101001011;
    rom[48219] = 25'b1111111011101111110111000;
    rom[48220] = 25'b1111111011110000000100110;
    rom[48221] = 25'b1111111011110000010010011;
    rom[48222] = 25'b1111111011110000100000001;
    rom[48223] = 25'b1111111011110000101101111;
    rom[48224] = 25'b1111111011110000111011110;
    rom[48225] = 25'b1111111011110001001001100;
    rom[48226] = 25'b1111111011110001010111010;
    rom[48227] = 25'b1111111011110001100101001;
    rom[48228] = 25'b1111111011110001110011000;
    rom[48229] = 25'b1111111011110010000000111;
    rom[48230] = 25'b1111111011110010001110110;
    rom[48231] = 25'b1111111011110010011100100;
    rom[48232] = 25'b1111111011110010101010100;
    rom[48233] = 25'b1111111011110010111000011;
    rom[48234] = 25'b1111111011110011000110011;
    rom[48235] = 25'b1111111011110011010100010;
    rom[48236] = 25'b1111111011110011100010011;
    rom[48237] = 25'b1111111011110011110000011;
    rom[48238] = 25'b1111111011110011111110011;
    rom[48239] = 25'b1111111011110100001100011;
    rom[48240] = 25'b1111111011110100011010011;
    rom[48241] = 25'b1111111011110100101000100;
    rom[48242] = 25'b1111111011110100110110100;
    rom[48243] = 25'b1111111011110101000100100;
    rom[48244] = 25'b1111111011110101010010101;
    rom[48245] = 25'b1111111011110101100000111;
    rom[48246] = 25'b1111111011110101101111000;
    rom[48247] = 25'b1111111011110101111101001;
    rom[48248] = 25'b1111111011110110001011010;
    rom[48249] = 25'b1111111011110110011001100;
    rom[48250] = 25'b1111111011110110100111101;
    rom[48251] = 25'b1111111011110110110101111;
    rom[48252] = 25'b1111111011110111000100001;
    rom[48253] = 25'b1111111011110111010010011;
    rom[48254] = 25'b1111111011110111100000101;
    rom[48255] = 25'b1111111011110111101110111;
    rom[48256] = 25'b1111111011110111111101001;
    rom[48257] = 25'b1111111011111000001011101;
    rom[48258] = 25'b1111111011111000011001111;
    rom[48259] = 25'b1111111011111000101000010;
    rom[48260] = 25'b1111111011111000110110101;
    rom[48261] = 25'b1111111011111001000101000;
    rom[48262] = 25'b1111111011111001010011011;
    rom[48263] = 25'b1111111011111001100001110;
    rom[48264] = 25'b1111111011111001110000010;
    rom[48265] = 25'b1111111011111001111110101;
    rom[48266] = 25'b1111111011111010001101001;
    rom[48267] = 25'b1111111011111010011011101;
    rom[48268] = 25'b1111111011111010101010000;
    rom[48269] = 25'b1111111011111010111000101;
    rom[48270] = 25'b1111111011111011000111001;
    rom[48271] = 25'b1111111011111011010101101;
    rom[48272] = 25'b1111111011111011100100010;
    rom[48273] = 25'b1111111011111011110010110;
    rom[48274] = 25'b1111111011111100000001011;
    rom[48275] = 25'b1111111011111100001111111;
    rom[48276] = 25'b1111111011111100011110101;
    rom[48277] = 25'b1111111011111100101101001;
    rom[48278] = 25'b1111111011111100111011111;
    rom[48279] = 25'b1111111011111101001010100;
    rom[48280] = 25'b1111111011111101011001001;
    rom[48281] = 25'b1111111011111101100111111;
    rom[48282] = 25'b1111111011111101110110100;
    rom[48283] = 25'b1111111011111110000101011;
    rom[48284] = 25'b1111111011111110010100000;
    rom[48285] = 25'b1111111011111110100010110;
    rom[48286] = 25'b1111111011111110110001101;
    rom[48287] = 25'b1111111011111111000000011;
    rom[48288] = 25'b1111111011111111001111001;
    rom[48289] = 25'b1111111011111111011110000;
    rom[48290] = 25'b1111111011111111101100110;
    rom[48291] = 25'b1111111011111111111011101;
    rom[48292] = 25'b1111111100000000001010100;
    rom[48293] = 25'b1111111100000000011001011;
    rom[48294] = 25'b1111111100000000101000001;
    rom[48295] = 25'b1111111100000000110111001;
    rom[48296] = 25'b1111111100000001000110001;
    rom[48297] = 25'b1111111100000001010101000;
    rom[48298] = 25'b1111111100000001100100000;
    rom[48299] = 25'b1111111100000001110010111;
    rom[48300] = 25'b1111111100000010000001111;
    rom[48301] = 25'b1111111100000010010000111;
    rom[48302] = 25'b1111111100000010011111110;
    rom[48303] = 25'b1111111100000010101110111;
    rom[48304] = 25'b1111111100000010111101111;
    rom[48305] = 25'b1111111100000011001100111;
    rom[48306] = 25'b1111111100000011011100000;
    rom[48307] = 25'b1111111100000011101011001;
    rom[48308] = 25'b1111111100000011111010010;
    rom[48309] = 25'b1111111100000100001001011;
    rom[48310] = 25'b1111111100000100011000100;
    rom[48311] = 25'b1111111100000100100111101;
    rom[48312] = 25'b1111111100000100110110110;
    rom[48313] = 25'b1111111100000101000101111;
    rom[48314] = 25'b1111111100000101010101001;
    rom[48315] = 25'b1111111100000101100100010;
    rom[48316] = 25'b1111111100000101110011011;
    rom[48317] = 25'b1111111100000110000010101;
    rom[48318] = 25'b1111111100000110010010000;
    rom[48319] = 25'b1111111100000110100001001;
    rom[48320] = 25'b1111111100000110110000011;
    rom[48321] = 25'b1111111100000110111111110;
    rom[48322] = 25'b1111111100000111001111000;
    rom[48323] = 25'b1111111100000111011110011;
    rom[48324] = 25'b1111111100000111101101101;
    rom[48325] = 25'b1111111100000111111101000;
    rom[48326] = 25'b1111111100001000001100010;
    rom[48327] = 25'b1111111100001000011011110;
    rom[48328] = 25'b1111111100001000101011000;
    rom[48329] = 25'b1111111100001000111010011;
    rom[48330] = 25'b1111111100001001001001111;
    rom[48331] = 25'b1111111100001001011001010;
    rom[48332] = 25'b1111111100001001101000110;
    rom[48333] = 25'b1111111100001001111000001;
    rom[48334] = 25'b1111111100001010000111101;
    rom[48335] = 25'b1111111100001010010111001;
    rom[48336] = 25'b1111111100001010100110101;
    rom[48337] = 25'b1111111100001010110110001;
    rom[48338] = 25'b1111111100001011000101101;
    rom[48339] = 25'b1111111100001011010101001;
    rom[48340] = 25'b1111111100001011100100101;
    rom[48341] = 25'b1111111100001011110100010;
    rom[48342] = 25'b1111111100001100000011110;
    rom[48343] = 25'b1111111100001100010011011;
    rom[48344] = 25'b1111111100001100100011000;
    rom[48345] = 25'b1111111100001100110010101;
    rom[48346] = 25'b1111111100001101000010010;
    rom[48347] = 25'b1111111100001101010001111;
    rom[48348] = 25'b1111111100001101100001100;
    rom[48349] = 25'b1111111100001101110001001;
    rom[48350] = 25'b1111111100001110000000111;
    rom[48351] = 25'b1111111100001110010000100;
    rom[48352] = 25'b1111111100001110100000010;
    rom[48353] = 25'b1111111100001110110000000;
    rom[48354] = 25'b1111111100001110111111101;
    rom[48355] = 25'b1111111100001111001111100;
    rom[48356] = 25'b1111111100001111011111001;
    rom[48357] = 25'b1111111100001111101110111;
    rom[48358] = 25'b1111111100001111111110110;
    rom[48359] = 25'b1111111100010000001110100;
    rom[48360] = 25'b1111111100010000011110011;
    rom[48361] = 25'b1111111100010000101110001;
    rom[48362] = 25'b1111111100010000111110000;
    rom[48363] = 25'b1111111100010001001101110;
    rom[48364] = 25'b1111111100010001011101101;
    rom[48365] = 25'b1111111100010001101101100;
    rom[48366] = 25'b1111111100010001111101011;
    rom[48367] = 25'b1111111100010010001101011;
    rom[48368] = 25'b1111111100010010011101010;
    rom[48369] = 25'b1111111100010010101101001;
    rom[48370] = 25'b1111111100010010111101001;
    rom[48371] = 25'b1111111100010011001101001;
    rom[48372] = 25'b1111111100010011011101000;
    rom[48373] = 25'b1111111100010011101101000;
    rom[48374] = 25'b1111111100010011111101000;
    rom[48375] = 25'b1111111100010100001101000;
    rom[48376] = 25'b1111111100010100011101000;
    rom[48377] = 25'b1111111100010100101101001;
    rom[48378] = 25'b1111111100010100111101001;
    rom[48379] = 25'b1111111100010101001101001;
    rom[48380] = 25'b1111111100010101011101010;
    rom[48381] = 25'b1111111100010101101101010;
    rom[48382] = 25'b1111111100010101111101011;
    rom[48383] = 25'b1111111100010110001101100;
    rom[48384] = 25'b1111111100010110011101100;
    rom[48385] = 25'b1111111100010110101101110;
    rom[48386] = 25'b1111111100010110111101111;
    rom[48387] = 25'b1111111100010111001110000;
    rom[48388] = 25'b1111111100010111011110001;
    rom[48389] = 25'b1111111100010111101110010;
    rom[48390] = 25'b1111111100010111111110100;
    rom[48391] = 25'b1111111100011000001110110;
    rom[48392] = 25'b1111111100011000011110111;
    rom[48393] = 25'b1111111100011000101111001;
    rom[48394] = 25'b1111111100011000111111011;
    rom[48395] = 25'b1111111100011001001111101;
    rom[48396] = 25'b1111111100011001011111111;
    rom[48397] = 25'b1111111100011001110000001;
    rom[48398] = 25'b1111111100011010000000100;
    rom[48399] = 25'b1111111100011010010000110;
    rom[48400] = 25'b1111111100011010100001000;
    rom[48401] = 25'b1111111100011010110001010;
    rom[48402] = 25'b1111111100011011000001101;
    rom[48403] = 25'b1111111100011011010010000;
    rom[48404] = 25'b1111111100011011100010011;
    rom[48405] = 25'b1111111100011011110010101;
    rom[48406] = 25'b1111111100011100000011001;
    rom[48407] = 25'b1111111100011100010011100;
    rom[48408] = 25'b1111111100011100100011111;
    rom[48409] = 25'b1111111100011100110100011;
    rom[48410] = 25'b1111111100011101000100101;
    rom[48411] = 25'b1111111100011101010101001;
    rom[48412] = 25'b1111111100011101100101101;
    rom[48413] = 25'b1111111100011101110110001;
    rom[48414] = 25'b1111111100011110000110100;
    rom[48415] = 25'b1111111100011110010111000;
    rom[48416] = 25'b1111111100011110100111100;
    rom[48417] = 25'b1111111100011110111000000;
    rom[48418] = 25'b1111111100011111001000100;
    rom[48419] = 25'b1111111100011111011001000;
    rom[48420] = 25'b1111111100011111101001101;
    rom[48421] = 25'b1111111100011111111010001;
    rom[48422] = 25'b1111111100100000001010101;
    rom[48423] = 25'b1111111100100000011011010;
    rom[48424] = 25'b1111111100100000101011110;
    rom[48425] = 25'b1111111100100000111100011;
    rom[48426] = 25'b1111111100100001001101000;
    rom[48427] = 25'b1111111100100001011101101;
    rom[48428] = 25'b1111111100100001101110010;
    rom[48429] = 25'b1111111100100001111110111;
    rom[48430] = 25'b1111111100100010001111100;
    rom[48431] = 25'b1111111100100010100000001;
    rom[48432] = 25'b1111111100100010110000111;
    rom[48433] = 25'b1111111100100011000001100;
    rom[48434] = 25'b1111111100100011010010010;
    rom[48435] = 25'b1111111100100011100010111;
    rom[48436] = 25'b1111111100100011110011101;
    rom[48437] = 25'b1111111100100100000100011;
    rom[48438] = 25'b1111111100100100010101001;
    rom[48439] = 25'b1111111100100100100101111;
    rom[48440] = 25'b1111111100100100110110101;
    rom[48441] = 25'b1111111100100101000111011;
    rom[48442] = 25'b1111111100100101011000001;
    rom[48443] = 25'b1111111100100101101001000;
    rom[48444] = 25'b1111111100100101111001110;
    rom[48445] = 25'b1111111100100110001010101;
    rom[48446] = 25'b1111111100100110011011011;
    rom[48447] = 25'b1111111100100110101100001;
    rom[48448] = 25'b1111111100100110111101000;
    rom[48449] = 25'b1111111100100111001101111;
    rom[48450] = 25'b1111111100100111011110110;
    rom[48451] = 25'b1111111100100111101111101;
    rom[48452] = 25'b1111111100101000000000100;
    rom[48453] = 25'b1111111100101000010001011;
    rom[48454] = 25'b1111111100101000100010011;
    rom[48455] = 25'b1111111100101000110011010;
    rom[48456] = 25'b1111111100101001000100001;
    rom[48457] = 25'b1111111100101001010101000;
    rom[48458] = 25'b1111111100101001100110000;
    rom[48459] = 25'b1111111100101001110110111;
    rom[48460] = 25'b1111111100101010000111111;
    rom[48461] = 25'b1111111100101010011000111;
    rom[48462] = 25'b1111111100101010101001111;
    rom[48463] = 25'b1111111100101010111010111;
    rom[48464] = 25'b1111111100101011001011111;
    rom[48465] = 25'b1111111100101011011100111;
    rom[48466] = 25'b1111111100101011101101111;
    rom[48467] = 25'b1111111100101011111110111;
    rom[48468] = 25'b1111111100101100010000000;
    rom[48469] = 25'b1111111100101100100001000;
    rom[48470] = 25'b1111111100101100110010001;
    rom[48471] = 25'b1111111100101101000011001;
    rom[48472] = 25'b1111111100101101010100010;
    rom[48473] = 25'b1111111100101101100101011;
    rom[48474] = 25'b1111111100101101110110011;
    rom[48475] = 25'b1111111100101110000111100;
    rom[48476] = 25'b1111111100101110011000101;
    rom[48477] = 25'b1111111100101110101001110;
    rom[48478] = 25'b1111111100101110111010111;
    rom[48479] = 25'b1111111100101111001100001;
    rom[48480] = 25'b1111111100101111011101010;
    rom[48481] = 25'b1111111100101111101110011;
    rom[48482] = 25'b1111111100101111111111101;
    rom[48483] = 25'b1111111100110000010000110;
    rom[48484] = 25'b1111111100110000100010000;
    rom[48485] = 25'b1111111100110000110011001;
    rom[48486] = 25'b1111111100110001000100011;
    rom[48487] = 25'b1111111100110001010101101;
    rom[48488] = 25'b1111111100110001100110110;
    rom[48489] = 25'b1111111100110001111000001;
    rom[48490] = 25'b1111111100110010001001011;
    rom[48491] = 25'b1111111100110010011010101;
    rom[48492] = 25'b1111111100110010101011111;
    rom[48493] = 25'b1111111100110010111101001;
    rom[48494] = 25'b1111111100110011001110100;
    rom[48495] = 25'b1111111100110011011111110;
    rom[48496] = 25'b1111111100110011110001000;
    rom[48497] = 25'b1111111100110100000010011;
    rom[48498] = 25'b1111111100110100010011101;
    rom[48499] = 25'b1111111100110100100101000;
    rom[48500] = 25'b1111111100110100110110011;
    rom[48501] = 25'b1111111100110101000111101;
    rom[48502] = 25'b1111111100110101011001000;
    rom[48503] = 25'b1111111100110101101010011;
    rom[48504] = 25'b1111111100110101111011110;
    rom[48505] = 25'b1111111100110110001101001;
    rom[48506] = 25'b1111111100110110011110101;
    rom[48507] = 25'b1111111100110110110000000;
    rom[48508] = 25'b1111111100110111000001011;
    rom[48509] = 25'b1111111100110111010010111;
    rom[48510] = 25'b1111111100110111100100010;
    rom[48511] = 25'b1111111100110111110101101;
    rom[48512] = 25'b1111111100111000000111001;
    rom[48513] = 25'b1111111100111000011000101;
    rom[48514] = 25'b1111111100111000101010000;
    rom[48515] = 25'b1111111100111000111011100;
    rom[48516] = 25'b1111111100111001001101000;
    rom[48517] = 25'b1111111100111001011110100;
    rom[48518] = 25'b1111111100111001110000000;
    rom[48519] = 25'b1111111100111010000001100;
    rom[48520] = 25'b1111111100111010010011000;
    rom[48521] = 25'b1111111100111010100100101;
    rom[48522] = 25'b1111111100111010110110001;
    rom[48523] = 25'b1111111100111011000111101;
    rom[48524] = 25'b1111111100111011011001001;
    rom[48525] = 25'b1111111100111011101010110;
    rom[48526] = 25'b1111111100111011111100010;
    rom[48527] = 25'b1111111100111100001101111;
    rom[48528] = 25'b1111111100111100011111100;
    rom[48529] = 25'b1111111100111100110001000;
    rom[48530] = 25'b1111111100111101000010101;
    rom[48531] = 25'b1111111100111101010100010;
    rom[48532] = 25'b1111111100111101100101111;
    rom[48533] = 25'b1111111100111101110111100;
    rom[48534] = 25'b1111111100111110001001001;
    rom[48535] = 25'b1111111100111110011010110;
    rom[48536] = 25'b1111111100111110101100011;
    rom[48537] = 25'b1111111100111110111110000;
    rom[48538] = 25'b1111111100111111001111110;
    rom[48539] = 25'b1111111100111111100001011;
    rom[48540] = 25'b1111111100111111110011001;
    rom[48541] = 25'b1111111101000000000100110;
    rom[48542] = 25'b1111111101000000010110011;
    rom[48543] = 25'b1111111101000000101000001;
    rom[48544] = 25'b1111111101000000111001110;
    rom[48545] = 25'b1111111101000001001011100;
    rom[48546] = 25'b1111111101000001011101010;
    rom[48547] = 25'b1111111101000001101111000;
    rom[48548] = 25'b1111111101000010000000110;
    rom[48549] = 25'b1111111101000010010010100;
    rom[48550] = 25'b1111111101000010100100010;
    rom[48551] = 25'b1111111101000010110110000;
    rom[48552] = 25'b1111111101000011000111110;
    rom[48553] = 25'b1111111101000011011001101;
    rom[48554] = 25'b1111111101000011101011011;
    rom[48555] = 25'b1111111101000011111101000;
    rom[48556] = 25'b1111111101000100001110111;
    rom[48557] = 25'b1111111101000100100000110;
    rom[48558] = 25'b1111111101000100110010100;
    rom[48559] = 25'b1111111101000101000100011;
    rom[48560] = 25'b1111111101000101010110001;
    rom[48561] = 25'b1111111101000101101000000;
    rom[48562] = 25'b1111111101000101111001111;
    rom[48563] = 25'b1111111101000110001011101;
    rom[48564] = 25'b1111111101000110011101100;
    rom[48565] = 25'b1111111101000110101111011;
    rom[48566] = 25'b1111111101000111000001010;
    rom[48567] = 25'b1111111101000111010011001;
    rom[48568] = 25'b1111111101000111100101000;
    rom[48569] = 25'b1111111101000111110110111;
    rom[48570] = 25'b1111111101001000001000110;
    rom[48571] = 25'b1111111101001000011010110;
    rom[48572] = 25'b1111111101001000101100101;
    rom[48573] = 25'b1111111101001000111110100;
    rom[48574] = 25'b1111111101001001010000011;
    rom[48575] = 25'b1111111101001001100010011;
    rom[48576] = 25'b1111111101001001110100010;
    rom[48577] = 25'b1111111101001010000110010;
    rom[48578] = 25'b1111111101001010011000010;
    rom[48579] = 25'b1111111101001010101010001;
    rom[48580] = 25'b1111111101001010111100001;
    rom[48581] = 25'b1111111101001011001110001;
    rom[48582] = 25'b1111111101001011100000000;
    rom[48583] = 25'b1111111101001011110010001;
    rom[48584] = 25'b1111111101001100000100000;
    rom[48585] = 25'b1111111101001100010110000;
    rom[48586] = 25'b1111111101001100101000000;
    rom[48587] = 25'b1111111101001100111010001;
    rom[48588] = 25'b1111111101001101001100001;
    rom[48589] = 25'b1111111101001101011110001;
    rom[48590] = 25'b1111111101001101110000001;
    rom[48591] = 25'b1111111101001110000010001;
    rom[48592] = 25'b1111111101001110010100010;
    rom[48593] = 25'b1111111101001110100110010;
    rom[48594] = 25'b1111111101001110111000010;
    rom[48595] = 25'b1111111101001111001010011;
    rom[48596] = 25'b1111111101001111011100011;
    rom[48597] = 25'b1111111101001111101110100;
    rom[48598] = 25'b1111111101010000000000100;
    rom[48599] = 25'b1111111101010000010010101;
    rom[48600] = 25'b1111111101010000100100110;
    rom[48601] = 25'b1111111101010000110110110;
    rom[48602] = 25'b1111111101010001001000111;
    rom[48603] = 25'b1111111101010001011011000;
    rom[48604] = 25'b1111111101010001101101001;
    rom[48605] = 25'b1111111101010001111111010;
    rom[48606] = 25'b1111111101010010010001011;
    rom[48607] = 25'b1111111101010010100011100;
    rom[48608] = 25'b1111111101010010110101110;
    rom[48609] = 25'b1111111101010011000111111;
    rom[48610] = 25'b1111111101010011011001111;
    rom[48611] = 25'b1111111101010011101100001;
    rom[48612] = 25'b1111111101010011111110010;
    rom[48613] = 25'b1111111101010100010000011;
    rom[48614] = 25'b1111111101010100100010101;
    rom[48615] = 25'b1111111101010100110100110;
    rom[48616] = 25'b1111111101010101000110111;
    rom[48617] = 25'b1111111101010101011001001;
    rom[48618] = 25'b1111111101010101101011011;
    rom[48619] = 25'b1111111101010101111101100;
    rom[48620] = 25'b1111111101010110001111110;
    rom[48621] = 25'b1111111101010110100010000;
    rom[48622] = 25'b1111111101010110110100001;
    rom[48623] = 25'b1111111101010111000110011;
    rom[48624] = 25'b1111111101010111011000101;
    rom[48625] = 25'b1111111101010111101010110;
    rom[48626] = 25'b1111111101010111111101001;
    rom[48627] = 25'b1111111101011000001111011;
    rom[48628] = 25'b1111111101011000100001100;
    rom[48629] = 25'b1111111101011000110011111;
    rom[48630] = 25'b1111111101011001000110000;
    rom[48631] = 25'b1111111101011001011000011;
    rom[48632] = 25'b1111111101011001101010101;
    rom[48633] = 25'b1111111101011001111100111;
    rom[48634] = 25'b1111111101011010001111001;
    rom[48635] = 25'b1111111101011010100001100;
    rom[48636] = 25'b1111111101011010110011101;
    rom[48637] = 25'b1111111101011011000110000;
    rom[48638] = 25'b1111111101011011011000010;
    rom[48639] = 25'b1111111101011011101010101;
    rom[48640] = 25'b1111111101011011111100111;
    rom[48641] = 25'b1111111101011100001111010;
    rom[48642] = 25'b1111111101011100100001100;
    rom[48643] = 25'b1111111101011100110011111;
    rom[48644] = 25'b1111111101011101000110010;
    rom[48645] = 25'b1111111101011101011000100;
    rom[48646] = 25'b1111111101011101101010111;
    rom[48647] = 25'b1111111101011101111101010;
    rom[48648] = 25'b1111111101011110001111100;
    rom[48649] = 25'b1111111101011110100001111;
    rom[48650] = 25'b1111111101011110110100010;
    rom[48651] = 25'b1111111101011111000110101;
    rom[48652] = 25'b1111111101011111011001000;
    rom[48653] = 25'b1111111101011111101011011;
    rom[48654] = 25'b1111111101011111111101110;
    rom[48655] = 25'b1111111101100000010000001;
    rom[48656] = 25'b1111111101100000100010100;
    rom[48657] = 25'b1111111101100000110100111;
    rom[48658] = 25'b1111111101100001000111010;
    rom[48659] = 25'b1111111101100001011001101;
    rom[48660] = 25'b1111111101100001101100000;
    rom[48661] = 25'b1111111101100001111110100;
    rom[48662] = 25'b1111111101100010010000111;
    rom[48663] = 25'b1111111101100010100011010;
    rom[48664] = 25'b1111111101100010110101110;
    rom[48665] = 25'b1111111101100011001000001;
    rom[48666] = 25'b1111111101100011011010101;
    rom[48667] = 25'b1111111101100011101101000;
    rom[48668] = 25'b1111111101100011111111011;
    rom[48669] = 25'b1111111101100100010001111;
    rom[48670] = 25'b1111111101100100100100010;
    rom[48671] = 25'b1111111101100100110110110;
    rom[48672] = 25'b1111111101100101001001001;
    rom[48673] = 25'b1111111101100101011011101;
    rom[48674] = 25'b1111111101100101101110000;
    rom[48675] = 25'b1111111101100110000000100;
    rom[48676] = 25'b1111111101100110010011000;
    rom[48677] = 25'b1111111101100110100101100;
    rom[48678] = 25'b1111111101100110110111111;
    rom[48679] = 25'b1111111101100111001010011;
    rom[48680] = 25'b1111111101100111011100111;
    rom[48681] = 25'b1111111101100111101111011;
    rom[48682] = 25'b1111111101101000000001111;
    rom[48683] = 25'b1111111101101000010100011;
    rom[48684] = 25'b1111111101101000100110111;
    rom[48685] = 25'b1111111101101000111001011;
    rom[48686] = 25'b1111111101101001001011111;
    rom[48687] = 25'b1111111101101001011110011;
    rom[48688] = 25'b1111111101101001110000111;
    rom[48689] = 25'b1111111101101010000011011;
    rom[48690] = 25'b1111111101101010010101111;
    rom[48691] = 25'b1111111101101010101000011;
    rom[48692] = 25'b1111111101101010111011000;
    rom[48693] = 25'b1111111101101011001101100;
    rom[48694] = 25'b1111111101101011100000000;
    rom[48695] = 25'b1111111101101011110010100;
    rom[48696] = 25'b1111111101101100000101001;
    rom[48697] = 25'b1111111101101100010111101;
    rom[48698] = 25'b1111111101101100101010001;
    rom[48699] = 25'b1111111101101100111100101;
    rom[48700] = 25'b1111111101101101001111010;
    rom[48701] = 25'b1111111101101101100001111;
    rom[48702] = 25'b1111111101101101110100011;
    rom[48703] = 25'b1111111101101110000110111;
    rom[48704] = 25'b1111111101101110011001100;
    rom[48705] = 25'b1111111101101110101100001;
    rom[48706] = 25'b1111111101101110111110101;
    rom[48707] = 25'b1111111101101111010001001;
    rom[48708] = 25'b1111111101101111100011110;
    rom[48709] = 25'b1111111101101111110110011;
    rom[48710] = 25'b1111111101110000001000111;
    rom[48711] = 25'b1111111101110000011011100;
    rom[48712] = 25'b1111111101110000101110001;
    rom[48713] = 25'b1111111101110001000000101;
    rom[48714] = 25'b1111111101110001010011010;
    rom[48715] = 25'b1111111101110001100101111;
    rom[48716] = 25'b1111111101110001111000011;
    rom[48717] = 25'b1111111101110010001011001;
    rom[48718] = 25'b1111111101110010011101101;
    rom[48719] = 25'b1111111101110010110000010;
    rom[48720] = 25'b1111111101110011000010111;
    rom[48721] = 25'b1111111101110011010101100;
    rom[48722] = 25'b1111111101110011101000001;
    rom[48723] = 25'b1111111101110011111010110;
    rom[48724] = 25'b1111111101110100001101011;
    rom[48725] = 25'b1111111101110100100000000;
    rom[48726] = 25'b1111111101110100110010100;
    rom[48727] = 25'b1111111101110101000101010;
    rom[48728] = 25'b1111111101110101010111110;
    rom[48729] = 25'b1111111101110101101010100;
    rom[48730] = 25'b1111111101110101111101000;
    rom[48731] = 25'b1111111101110110001111110;
    rom[48732] = 25'b1111111101110110100010011;
    rom[48733] = 25'b1111111101110110110101000;
    rom[48734] = 25'b1111111101110111000111101;
    rom[48735] = 25'b1111111101110111011010010;
    rom[48736] = 25'b1111111101110111101100111;
    rom[48737] = 25'b1111111101110111111111101;
    rom[48738] = 25'b1111111101111000010010010;
    rom[48739] = 25'b1111111101111000100100111;
    rom[48740] = 25'b1111111101111000110111100;
    rom[48741] = 25'b1111111101111001001010010;
    rom[48742] = 25'b1111111101111001011100111;
    rom[48743] = 25'b1111111101111001101111100;
    rom[48744] = 25'b1111111101111010000010001;
    rom[48745] = 25'b1111111101111010010100111;
    rom[48746] = 25'b1111111101111010100111100;
    rom[48747] = 25'b1111111101111010111010010;
    rom[48748] = 25'b1111111101111011001100111;
    rom[48749] = 25'b1111111101111011011111100;
    rom[48750] = 25'b1111111101111011110010010;
    rom[48751] = 25'b1111111101111100000100111;
    rom[48752] = 25'b1111111101111100010111101;
    rom[48753] = 25'b1111111101111100101010010;
    rom[48754] = 25'b1111111101111100111101000;
    rom[48755] = 25'b1111111101111101001111101;
    rom[48756] = 25'b1111111101111101100010010;
    rom[48757] = 25'b1111111101111101110101000;
    rom[48758] = 25'b1111111101111110000111101;
    rom[48759] = 25'b1111111101111110011010011;
    rom[48760] = 25'b1111111101111110101101000;
    rom[48761] = 25'b1111111101111110111111110;
    rom[48762] = 25'b1111111101111111010010100;
    rom[48763] = 25'b1111111101111111100101001;
    rom[48764] = 25'b1111111101111111110111110;
    rom[48765] = 25'b1111111110000000001010100;
    rom[48766] = 25'b1111111110000000011101010;
    rom[48767] = 25'b1111111110000000101111111;
    rom[48768] = 25'b1111111110000001000010101;
    rom[48769] = 25'b1111111110000001010101010;
    rom[48770] = 25'b1111111110000001101000000;
    rom[48771] = 25'b1111111110000001111010110;
    rom[48772] = 25'b1111111110000010001101011;
    rom[48773] = 25'b1111111110000010100000001;
    rom[48774] = 25'b1111111110000010110010111;
    rom[48775] = 25'b1111111110000011000101100;
    rom[48776] = 25'b1111111110000011011000011;
    rom[48777] = 25'b1111111110000011101011000;
    rom[48778] = 25'b1111111110000011111101110;
    rom[48779] = 25'b1111111110000100010000100;
    rom[48780] = 25'b1111111110000100100011001;
    rom[48781] = 25'b1111111110000100110101111;
    rom[48782] = 25'b1111111110000101001000101;
    rom[48783] = 25'b1111111110000101011011011;
    rom[48784] = 25'b1111111110000101101110000;
    rom[48785] = 25'b1111111110000110000000110;
    rom[48786] = 25'b1111111110000110010011100;
    rom[48787] = 25'b1111111110000110100110010;
    rom[48788] = 25'b1111111110000110111000111;
    rom[48789] = 25'b1111111110000111001011101;
    rom[48790] = 25'b1111111110000111011110011;
    rom[48791] = 25'b1111111110000111110001001;
    rom[48792] = 25'b1111111110001000000011110;
    rom[48793] = 25'b1111111110001000010110101;
    rom[48794] = 25'b1111111110001000101001010;
    rom[48795] = 25'b1111111110001000111100000;
    rom[48796] = 25'b1111111110001001001110110;
    rom[48797] = 25'b1111111110001001100001100;
    rom[48798] = 25'b1111111110001001110100010;
    rom[48799] = 25'b1111111110001010000110111;
    rom[48800] = 25'b1111111110001010011001110;
    rom[48801] = 25'b1111111110001010101100011;
    rom[48802] = 25'b1111111110001010111111001;
    rom[48803] = 25'b1111111110001011010001111;
    rom[48804] = 25'b1111111110001011100100101;
    rom[48805] = 25'b1111111110001011110111011;
    rom[48806] = 25'b1111111110001100001010000;
    rom[48807] = 25'b1111111110001100011100110;
    rom[48808] = 25'b1111111110001100101111101;
    rom[48809] = 25'b1111111110001101000010010;
    rom[48810] = 25'b1111111110001101010101000;
    rom[48811] = 25'b1111111110001101100111110;
    rom[48812] = 25'b1111111110001101111010100;
    rom[48813] = 25'b1111111110001110001101010;
    rom[48814] = 25'b1111111110001110011111111;
    rom[48815] = 25'b1111111110001110110010110;
    rom[48816] = 25'b1111111110001111000101011;
    rom[48817] = 25'b1111111110001111011000001;
    rom[48818] = 25'b1111111110001111101010111;
    rom[48819] = 25'b1111111110001111111101101;
    rom[48820] = 25'b1111111110010000010000011;
    rom[48821] = 25'b1111111110010000100011001;
    rom[48822] = 25'b1111111110010000110101110;
    rom[48823] = 25'b1111111110010001001000101;
    rom[48824] = 25'b1111111110010001011011010;
    rom[48825] = 25'b1111111110010001101110000;
    rom[48826] = 25'b1111111110010010000000110;
    rom[48827] = 25'b1111111110010010010011100;
    rom[48828] = 25'b1111111110010010100110010;
    rom[48829] = 25'b1111111110010010111001000;
    rom[48830] = 25'b1111111110010011001011110;
    rom[48831] = 25'b1111111110010011011110100;
    rom[48832] = 25'b1111111110010011110001001;
    rom[48833] = 25'b1111111110010100000011111;
    rom[48834] = 25'b1111111110010100010110101;
    rom[48835] = 25'b1111111110010100101001011;
    rom[48836] = 25'b1111111110010100111100001;
    rom[48837] = 25'b1111111110010101001110110;
    rom[48838] = 25'b1111111110010101100001101;
    rom[48839] = 25'b1111111110010101110100010;
    rom[48840] = 25'b1111111110010110000111000;
    rom[48841] = 25'b1111111110010110011001110;
    rom[48842] = 25'b1111111110010110101100100;
    rom[48843] = 25'b1111111110010110111111010;
    rom[48844] = 25'b1111111110010111010001111;
    rom[48845] = 25'b1111111110010111100100110;
    rom[48846] = 25'b1111111110010111110111011;
    rom[48847] = 25'b1111111110011000001010001;
    rom[48848] = 25'b1111111110011000011100111;
    rom[48849] = 25'b1111111110011000101111101;
    rom[48850] = 25'b1111111110011001000010010;
    rom[48851] = 25'b1111111110011001010101000;
    rom[48852] = 25'b1111111110011001100111110;
    rom[48853] = 25'b1111111110011001111010011;
    rom[48854] = 25'b1111111110011010001101001;
    rom[48855] = 25'b1111111110011010011111111;
    rom[48856] = 25'b1111111110011010110010101;
    rom[48857] = 25'b1111111110011011000101010;
    rom[48858] = 25'b1111111110011011011000000;
    rom[48859] = 25'b1111111110011011101010110;
    rom[48860] = 25'b1111111110011011111101011;
    rom[48861] = 25'b1111111110011100010000010;
    rom[48862] = 25'b1111111110011100100010111;
    rom[48863] = 25'b1111111110011100110101100;
    rom[48864] = 25'b1111111110011101001000011;
    rom[48865] = 25'b1111111110011101011011000;
    rom[48866] = 25'b1111111110011101101101101;
    rom[48867] = 25'b1111111110011110000000100;
    rom[48868] = 25'b1111111110011110010011001;
    rom[48869] = 25'b1111111110011110100101110;
    rom[48870] = 25'b1111111110011110111000100;
    rom[48871] = 25'b1111111110011111001011010;
    rom[48872] = 25'b1111111110011111011101111;
    rom[48873] = 25'b1111111110011111110000101;
    rom[48874] = 25'b1111111110100000000011010;
    rom[48875] = 25'b1111111110100000010110000;
    rom[48876] = 25'b1111111110100000101000101;
    rom[48877] = 25'b1111111110100000111011011;
    rom[48878] = 25'b1111111110100001001110001;
    rom[48879] = 25'b1111111110100001100000110;
    rom[48880] = 25'b1111111110100001110011011;
    rom[48881] = 25'b1111111110100010000110001;
    rom[48882] = 25'b1111111110100010011000110;
    rom[48883] = 25'b1111111110100010101011100;
    rom[48884] = 25'b1111111110100010111110001;
    rom[48885] = 25'b1111111110100011010000111;
    rom[48886] = 25'b1111111110100011100011100;
    rom[48887] = 25'b1111111110100011110110001;
    rom[48888] = 25'b1111111110100100001000111;
    rom[48889] = 25'b1111111110100100011011100;
    rom[48890] = 25'b1111111110100100101110010;
    rom[48891] = 25'b1111111110100101000000111;
    rom[48892] = 25'b1111111110100101010011100;
    rom[48893] = 25'b1111111110100101100110001;
    rom[48894] = 25'b1111111110100101111000111;
    rom[48895] = 25'b1111111110100110001011100;
    rom[48896] = 25'b1111111110100110011110001;
    rom[48897] = 25'b1111111110100110110000110;
    rom[48898] = 25'b1111111110100111000011100;
    rom[48899] = 25'b1111111110100111010110001;
    rom[48900] = 25'b1111111110100111101000110;
    rom[48901] = 25'b1111111110100111111011011;
    rom[48902] = 25'b1111111110101000001110000;
    rom[48903] = 25'b1111111110101000100000101;
    rom[48904] = 25'b1111111110101000110011011;
    rom[48905] = 25'b1111111110101001000101111;
    rom[48906] = 25'b1111111110101001011000101;
    rom[48907] = 25'b1111111110101001101011010;
    rom[48908] = 25'b1111111110101001111101111;
    rom[48909] = 25'b1111111110101010010000011;
    rom[48910] = 25'b1111111110101010100011001;
    rom[48911] = 25'b1111111110101010110101101;
    rom[48912] = 25'b1111111110101011001000011;
    rom[48913] = 25'b1111111110101011011011000;
    rom[48914] = 25'b1111111110101011101101100;
    rom[48915] = 25'b1111111110101100000000010;
    rom[48916] = 25'b1111111110101100010010110;
    rom[48917] = 25'b1111111110101100100101011;
    rom[48918] = 25'b1111111110101100111000000;
    rom[48919] = 25'b1111111110101101001010101;
    rom[48920] = 25'b1111111110101101011101010;
    rom[48921] = 25'b1111111110101101101111110;
    rom[48922] = 25'b1111111110101110000010011;
    rom[48923] = 25'b1111111110101110010101000;
    rom[48924] = 25'b1111111110101110100111100;
    rom[48925] = 25'b1111111110101110111010001;
    rom[48926] = 25'b1111111110101111001100110;
    rom[48927] = 25'b1111111110101111011111010;
    rom[48928] = 25'b1111111110101111110001111;
    rom[48929] = 25'b1111111110110000000100100;
    rom[48930] = 25'b1111111110110000010111000;
    rom[48931] = 25'b1111111110110000101001101;
    rom[48932] = 25'b1111111110110000111100010;
    rom[48933] = 25'b1111111110110001001110110;
    rom[48934] = 25'b1111111110110001100001010;
    rom[48935] = 25'b1111111110110001110011111;
    rom[48936] = 25'b1111111110110010000110100;
    rom[48937] = 25'b1111111110110010011001000;
    rom[48938] = 25'b1111111110110010101011100;
    rom[48939] = 25'b1111111110110010111110000;
    rom[48940] = 25'b1111111110110011010000101;
    rom[48941] = 25'b1111111110110011100011010;
    rom[48942] = 25'b1111111110110011110101110;
    rom[48943] = 25'b1111111110110100001000001;
    rom[48944] = 25'b1111111110110100011010110;
    rom[48945] = 25'b1111111110110100101101010;
    rom[48946] = 25'b1111111110110100111111111;
    rom[48947] = 25'b1111111110110101010010011;
    rom[48948] = 25'b1111111110110101100100111;
    rom[48949] = 25'b1111111110110101110111011;
    rom[48950] = 25'b1111111110110110001001111;
    rom[48951] = 25'b1111111110110110011100011;
    rom[48952] = 25'b1111111110110110101110111;
    rom[48953] = 25'b1111111110110111000001011;
    rom[48954] = 25'b1111111110110111010011111;
    rom[48955] = 25'b1111111110110111100110011;
    rom[48956] = 25'b1111111110110111111000111;
    rom[48957] = 25'b1111111110111000001011011;
    rom[48958] = 25'b1111111110111000011101111;
    rom[48959] = 25'b1111111110111000110000011;
    rom[48960] = 25'b1111111110111001000010110;
    rom[48961] = 25'b1111111110111001010101010;
    rom[48962] = 25'b1111111110111001100111110;
    rom[48963] = 25'b1111111110111001111010001;
    rom[48964] = 25'b1111111110111010001100101;
    rom[48965] = 25'b1111111110111010011111001;
    rom[48966] = 25'b1111111110111010110001101;
    rom[48967] = 25'b1111111110111011000100000;
    rom[48968] = 25'b1111111110111011010110100;
    rom[48969] = 25'b1111111110111011101000111;
    rom[48970] = 25'b1111111110111011111011011;
    rom[48971] = 25'b1111111110111100001101110;
    rom[48972] = 25'b1111111110111100100000010;
    rom[48973] = 25'b1111111110111100110010101;
    rom[48974] = 25'b1111111110111101000101000;
    rom[48975] = 25'b1111111110111101010111011;
    rom[48976] = 25'b1111111110111101101001111;
    rom[48977] = 25'b1111111110111101111100010;
    rom[48978] = 25'b1111111110111110001110110;
    rom[48979] = 25'b1111111110111110100001001;
    rom[48980] = 25'b1111111110111110110011100;
    rom[48981] = 25'b1111111110111111000101111;
    rom[48982] = 25'b1111111110111111011000010;
    rom[48983] = 25'b1111111110111111101010110;
    rom[48984] = 25'b1111111110111111111101001;
    rom[48985] = 25'b1111111111000000001111011;
    rom[48986] = 25'b1111111111000000100001110;
    rom[48987] = 25'b1111111111000000110100001;
    rom[48988] = 25'b1111111111000001000110100;
    rom[48989] = 25'b1111111111000001011000111;
    rom[48990] = 25'b1111111111000001101011010;
    rom[48991] = 25'b1111111111000001111101101;
    rom[48992] = 25'b1111111111000010010000000;
    rom[48993] = 25'b1111111111000010100010010;
    rom[48994] = 25'b1111111111000010110100101;
    rom[48995] = 25'b1111111111000011000111000;
    rom[48996] = 25'b1111111111000011011001010;
    rom[48997] = 25'b1111111111000011101011101;
    rom[48998] = 25'b1111111111000011111101111;
    rom[48999] = 25'b1111111111000100010000010;
    rom[49000] = 25'b1111111111000100100010101;
    rom[49001] = 25'b1111111111000100110100111;
    rom[49002] = 25'b1111111111000101000111010;
    rom[49003] = 25'b1111111111000101011001100;
    rom[49004] = 25'b1111111111000101101011110;
    rom[49005] = 25'b1111111111000101111110000;
    rom[49006] = 25'b1111111111000110010000011;
    rom[49007] = 25'b1111111111000110100010101;
    rom[49008] = 25'b1111111111000110110100111;
    rom[49009] = 25'b1111111111000111000111001;
    rom[49010] = 25'b1111111111000111011001100;
    rom[49011] = 25'b1111111111000111101011101;
    rom[49012] = 25'b1111111111000111111110000;
    rom[49013] = 25'b1111111111001000010000001;
    rom[49014] = 25'b1111111111001000100010100;
    rom[49015] = 25'b1111111111001000110100110;
    rom[49016] = 25'b1111111111001001000110111;
    rom[49017] = 25'b1111111111001001011001001;
    rom[49018] = 25'b1111111111001001101011011;
    rom[49019] = 25'b1111111111001001111101101;
    rom[49020] = 25'b1111111111001010001111111;
    rom[49021] = 25'b1111111111001010100010000;
    rom[49022] = 25'b1111111111001010110100010;
    rom[49023] = 25'b1111111111001011000110100;
    rom[49024] = 25'b1111111111001011011000101;
    rom[49025] = 25'b1111111111001011101010110;
    rom[49026] = 25'b1111111111001011111101000;
    rom[49027] = 25'b1111111111001100001111010;
    rom[49028] = 25'b1111111111001100100001011;
    rom[49029] = 25'b1111111111001100110011100;
    rom[49030] = 25'b1111111111001101000101101;
    rom[49031] = 25'b1111111111001101010111111;
    rom[49032] = 25'b1111111111001101101010000;
    rom[49033] = 25'b1111111111001101111100001;
    rom[49034] = 25'b1111111111001110001110011;
    rom[49035] = 25'b1111111111001110100000011;
    rom[49036] = 25'b1111111111001110110010100;
    rom[49037] = 25'b1111111111001111000100101;
    rom[49038] = 25'b1111111111001111010110110;
    rom[49039] = 25'b1111111111001111101000111;
    rom[49040] = 25'b1111111111001111111011000;
    rom[49041] = 25'b1111111111010000001101001;
    rom[49042] = 25'b1111111111010000011111010;
    rom[49043] = 25'b1111111111010000110001011;
    rom[49044] = 25'b1111111111010001000011011;
    rom[49045] = 25'b1111111111010001010101100;
    rom[49046] = 25'b1111111111010001100111101;
    rom[49047] = 25'b1111111111010001111001101;
    rom[49048] = 25'b1111111111010010001011110;
    rom[49049] = 25'b1111111111010010011101110;
    rom[49050] = 25'b1111111111010010101111111;
    rom[49051] = 25'b1111111111010011000001111;
    rom[49052] = 25'b1111111111010011010100000;
    rom[49053] = 25'b1111111111010011100110000;
    rom[49054] = 25'b1111111111010011111000000;
    rom[49055] = 25'b1111111111010100001010000;
    rom[49056] = 25'b1111111111010100011100000;
    rom[49057] = 25'b1111111111010100101110001;
    rom[49058] = 25'b1111111111010101000000001;
    rom[49059] = 25'b1111111111010101010010001;
    rom[49060] = 25'b1111111111010101100100000;
    rom[49061] = 25'b1111111111010101110110001;
    rom[49062] = 25'b1111111111010110001000001;
    rom[49063] = 25'b1111111111010110011010000;
    rom[49064] = 25'b1111111111010110101100000;
    rom[49065] = 25'b1111111111010110111110000;
    rom[49066] = 25'b1111111111010111001111111;
    rom[49067] = 25'b1111111111010111100001111;
    rom[49068] = 25'b1111111111010111110011111;
    rom[49069] = 25'b1111111111011000000101110;
    rom[49070] = 25'b1111111111011000010111110;
    rom[49071] = 25'b1111111111011000101001101;
    rom[49072] = 25'b1111111111011000111011101;
    rom[49073] = 25'b1111111111011001001101100;
    rom[49074] = 25'b1111111111011001011111100;
    rom[49075] = 25'b1111111111011001110001010;
    rom[49076] = 25'b1111111111011010000011010;
    rom[49077] = 25'b1111111111011010010101001;
    rom[49078] = 25'b1111111111011010100111000;
    rom[49079] = 25'b1111111111011010111000111;
    rom[49080] = 25'b1111111111011011001010110;
    rom[49081] = 25'b1111111111011011011100101;
    rom[49082] = 25'b1111111111011011101110100;
    rom[49083] = 25'b1111111111011100000000011;
    rom[49084] = 25'b1111111111011100010010010;
    rom[49085] = 25'b1111111111011100100100000;
    rom[49086] = 25'b1111111111011100110101111;
    rom[49087] = 25'b1111111111011101000111110;
    rom[49088] = 25'b1111111111011101011001100;
    rom[49089] = 25'b1111111111011101101011010;
    rom[49090] = 25'b1111111111011101111101001;
    rom[49091] = 25'b1111111111011110001111000;
    rom[49092] = 25'b1111111111011110100000110;
    rom[49093] = 25'b1111111111011110110010100;
    rom[49094] = 25'b1111111111011111000100010;
    rom[49095] = 25'b1111111111011111010110001;
    rom[49096] = 25'b1111111111011111100111111;
    rom[49097] = 25'b1111111111011111111001101;
    rom[49098] = 25'b1111111111100000001011011;
    rom[49099] = 25'b1111111111100000011101001;
    rom[49100] = 25'b1111111111100000101110111;
    rom[49101] = 25'b1111111111100001000000101;
    rom[49102] = 25'b1111111111100001010010011;
    rom[49103] = 25'b1111111111100001100100001;
    rom[49104] = 25'b1111111111100001110101110;
    rom[49105] = 25'b1111111111100010000111100;
    rom[49106] = 25'b1111111111100010011001010;
    rom[49107] = 25'b1111111111100010101010111;
    rom[49108] = 25'b1111111111100010111100100;
    rom[49109] = 25'b1111111111100011001110010;
    rom[49110] = 25'b1111111111100011011111111;
    rom[49111] = 25'b1111111111100011110001100;
    rom[49112] = 25'b1111111111100100000011010;
    rom[49113] = 25'b1111111111100100010100111;
    rom[49114] = 25'b1111111111100100100110100;
    rom[49115] = 25'b1111111111100100111000001;
    rom[49116] = 25'b1111111111100101001001110;
    rom[49117] = 25'b1111111111100101011011100;
    rom[49118] = 25'b1111111111100101101101000;
    rom[49119] = 25'b1111111111100101111110101;
    rom[49120] = 25'b1111111111100110010000010;
    rom[49121] = 25'b1111111111100110100001111;
    rom[49122] = 25'b1111111111100110110011011;
    rom[49123] = 25'b1111111111100111000101000;
    rom[49124] = 25'b1111111111100111010110101;
    rom[49125] = 25'b1111111111100111101000010;
    rom[49126] = 25'b1111111111100111111001110;
    rom[49127] = 25'b1111111111101000001011010;
    rom[49128] = 25'b1111111111101000011100110;
    rom[49129] = 25'b1111111111101000101110011;
    rom[49130] = 25'b1111111111101000111111111;
    rom[49131] = 25'b1111111111101001010001011;
    rom[49132] = 25'b1111111111101001100010111;
    rom[49133] = 25'b1111111111101001110100100;
    rom[49134] = 25'b1111111111101010000101111;
    rom[49135] = 25'b1111111111101010010111011;
    rom[49136] = 25'b1111111111101010101000111;
    rom[49137] = 25'b1111111111101010111010011;
    rom[49138] = 25'b1111111111101011001011111;
    rom[49139] = 25'b1111111111101011011101011;
    rom[49140] = 25'b1111111111101011101110110;
    rom[49141] = 25'b1111111111101100000000001;
    rom[49142] = 25'b1111111111101100010001101;
    rom[49143] = 25'b1111111111101100100011001;
    rom[49144] = 25'b1111111111101100110100100;
    rom[49145] = 25'b1111111111101101000101111;
    rom[49146] = 25'b1111111111101101010111010;
    rom[49147] = 25'b1111111111101101101000110;
    rom[49148] = 25'b1111111111101101111010001;
    rom[49149] = 25'b1111111111101110001011100;
    rom[49150] = 25'b1111111111101110011100111;
    rom[49151] = 25'b1111111111101110101110010;
    rom[49152] = 25'b1111111111101110111111101;
    rom[49153] = 25'b1111111111101111010001000;
    rom[49154] = 25'b1111111111101111100010010;
    rom[49155] = 25'b1111111111101111110011101;
    rom[49156] = 25'b1111111111110000000101000;
    rom[49157] = 25'b1111111111110000010110010;
    rom[49158] = 25'b1111111111110000100111100;
    rom[49159] = 25'b1111111111110000111000111;
    rom[49160] = 25'b1111111111110001001010010;
    rom[49161] = 25'b1111111111110001011011100;
    rom[49162] = 25'b1111111111110001101100110;
    rom[49163] = 25'b1111111111110001111110000;
    rom[49164] = 25'b1111111111110010001111010;
    rom[49165] = 25'b1111111111110010100000101;
    rom[49166] = 25'b1111111111110010110001110;
    rom[49167] = 25'b1111111111110011000011000;
    rom[49168] = 25'b1111111111110011010100010;
    rom[49169] = 25'b1111111111110011100101100;
    rom[49170] = 25'b1111111111110011110110101;
    rom[49171] = 25'b1111111111110100001000000;
    rom[49172] = 25'b1111111111110100011001001;
    rom[49173] = 25'b1111111111110100101010011;
    rom[49174] = 25'b1111111111110100111011100;
    rom[49175] = 25'b1111111111110101001100101;
    rom[49176] = 25'b1111111111110101011101111;
    rom[49177] = 25'b1111111111110101101111000;
    rom[49178] = 25'b1111111111110110000000001;
    rom[49179] = 25'b1111111111110110010001010;
    rom[49180] = 25'b1111111111110110100010011;
    rom[49181] = 25'b1111111111110110110011100;
    rom[49182] = 25'b1111111111110111000100110;
    rom[49183] = 25'b1111111111110111010101110;
    rom[49184] = 25'b1111111111110111100110111;
    rom[49185] = 25'b1111111111110111111000000;
    rom[49186] = 25'b1111111111111000001001000;
    rom[49187] = 25'b1111111111111000011010001;
    rom[49188] = 25'b1111111111111000101011001;
    rom[49189] = 25'b1111111111111000111100010;
    rom[49190] = 25'b1111111111111001001101010;
    rom[49191] = 25'b1111111111111001011110010;
    rom[49192] = 25'b1111111111111001101111010;
    rom[49193] = 25'b1111111111111010000000010;
    rom[49194] = 25'b1111111111111010010001011;
    rom[49195] = 25'b1111111111111010100010011;
    rom[49196] = 25'b1111111111111010110011011;
    rom[49197] = 25'b1111111111111011000100011;
    rom[49198] = 25'b1111111111111011010101010;
    rom[49199] = 25'b1111111111111011100110010;
    rom[49200] = 25'b1111111111111011110111010;
    rom[49201] = 25'b1111111111111100001000001;
    rom[49202] = 25'b1111111111111100011001001;
    rom[49203] = 25'b1111111111111100101010001;
    rom[49204] = 25'b1111111111111100111011000;
    rom[49205] = 25'b1111111111111101001011111;
    rom[49206] = 25'b1111111111111101011100110;
    rom[49207] = 25'b1111111111111101101101110;
    rom[49208] = 25'b1111111111111101111110101;
    rom[49209] = 25'b1111111111111110001111100;
    rom[49210] = 25'b1111111111111110100000010;
    rom[49211] = 25'b1111111111111110110001010;
    rom[49212] = 25'b1111111111111111000010000;
    rom[49213] = 25'b1111111111111111010010111;
    rom[49214] = 25'b1111111111111111100011110;
    rom[49215] = 25'b1111111111111111110100100;
    rom[49216] = 25'b0000000000000000000101010;
    rom[49217] = 25'b0000000000000000010110001;
    rom[49218] = 25'b0000000000000000100110111;
    rom[49219] = 25'b0000000000000000110111110;
    rom[49220] = 25'b0000000000000001001000100;
    rom[49221] = 25'b0000000000000001011001010;
    rom[49222] = 25'b0000000000000001101010000;
    rom[49223] = 25'b0000000000000001111010110;
    rom[49224] = 25'b0000000000000010001011100;
    rom[49225] = 25'b0000000000000010011100001;
    rom[49226] = 25'b0000000000000010101100111;
    rom[49227] = 25'b0000000000000010111101101;
    rom[49228] = 25'b0000000000000011001110011;
    rom[49229] = 25'b0000000000000011011111000;
    rom[49230] = 25'b0000000000000011101111110;
    rom[49231] = 25'b0000000000000100000000011;
    rom[49232] = 25'b0000000000000100010001001;
    rom[49233] = 25'b0000000000000100100001110;
    rom[49234] = 25'b0000000000000100110010011;
    rom[49235] = 25'b0000000000000101000011000;
    rom[49236] = 25'b0000000000000101010011101;
    rom[49237] = 25'b0000000000000101100100010;
    rom[49238] = 25'b0000000000000101110100111;
    rom[49239] = 25'b0000000000000110000101100;
    rom[49240] = 25'b0000000000000110010110001;
    rom[49241] = 25'b0000000000000110100110101;
    rom[49242] = 25'b0000000000000110110111010;
    rom[49243] = 25'b0000000000000111000111110;
    rom[49244] = 25'b0000000000000111011000011;
    rom[49245] = 25'b0000000000000111101000111;
    rom[49246] = 25'b0000000000000111111001100;
    rom[49247] = 25'b0000000000001000001010000;
    rom[49248] = 25'b0000000000001000011010011;
    rom[49249] = 25'b0000000000001000101010111;
    rom[49250] = 25'b0000000000001000111011100;
    rom[49251] = 25'b0000000000001001001011111;
    rom[49252] = 25'b0000000000001001011100011;
    rom[49253] = 25'b0000000000001001101100111;
    rom[49254] = 25'b0000000000001001111101010;
    rom[49255] = 25'b0000000000001010001101110;
    rom[49256] = 25'b0000000000001010011110001;
    rom[49257] = 25'b0000000000001010101110101;
    rom[49258] = 25'b0000000000001010111111000;
    rom[49259] = 25'b0000000000001011001111100;
    rom[49260] = 25'b0000000000001011011111111;
    rom[49261] = 25'b0000000000001011110000010;
    rom[49262] = 25'b0000000000001100000000101;
    rom[49263] = 25'b0000000000001100010001000;
    rom[49264] = 25'b0000000000001100100001010;
    rom[49265] = 25'b0000000000001100110001110;
    rom[49266] = 25'b0000000000001101000010000;
    rom[49267] = 25'b0000000000001101010010011;
    rom[49268] = 25'b0000000000001101100010101;
    rom[49269] = 25'b0000000000001101110011000;
    rom[49270] = 25'b0000000000001110000011010;
    rom[49271] = 25'b0000000000001110010011100;
    rom[49272] = 25'b0000000000001110100011111;
    rom[49273] = 25'b0000000000001110110100001;
    rom[49274] = 25'b0000000000001111000100011;
    rom[49275] = 25'b0000000000001111010100101;
    rom[49276] = 25'b0000000000001111100100111;
    rom[49277] = 25'b0000000000001111110101000;
    rom[49278] = 25'b0000000000010000000101010;
    rom[49279] = 25'b0000000000010000010101100;
    rom[49280] = 25'b0000000000010000100101101;
    rom[49281] = 25'b0000000000010000110101110;
    rom[49282] = 25'b0000000000010001000110000;
    rom[49283] = 25'b0000000000010001010110010;
    rom[49284] = 25'b0000000000010001100110011;
    rom[49285] = 25'b0000000000010001110110011;
    rom[49286] = 25'b0000000000010010000110101;
    rom[49287] = 25'b0000000000010010010110110;
    rom[49288] = 25'b0000000000010010100110110;
    rom[49289] = 25'b0000000000010010110111000;
    rom[49290] = 25'b0000000000010011000111000;
    rom[49291] = 25'b0000000000010011010111001;
    rom[49292] = 25'b0000000000010011100111001;
    rom[49293] = 25'b0000000000010011110111010;
    rom[49294] = 25'b0000000000010100000111010;
    rom[49295] = 25'b0000000000010100010111011;
    rom[49296] = 25'b0000000000010100100111010;
    rom[49297] = 25'b0000000000010100110111011;
    rom[49298] = 25'b0000000000010101000111011;
    rom[49299] = 25'b0000000000010101010111010;
    rom[49300] = 25'b0000000000010101100111011;
    rom[49301] = 25'b0000000000010101110111011;
    rom[49302] = 25'b0000000000010110000111010;
    rom[49303] = 25'b0000000000010110010111001;
    rom[49304] = 25'b0000000000010110100111001;
    rom[49305] = 25'b0000000000010110110111001;
    rom[49306] = 25'b0000000000010111000111000;
    rom[49307] = 25'b0000000000010111010111000;
    rom[49308] = 25'b0000000000010111100110111;
    rom[49309] = 25'b0000000000010111110110110;
    rom[49310] = 25'b0000000000011000000110101;
    rom[49311] = 25'b0000000000011000010110100;
    rom[49312] = 25'b0000000000011000100110011;
    rom[49313] = 25'b0000000000011000110110001;
    rom[49314] = 25'b0000000000011001000110000;
    rom[49315] = 25'b0000000000011001010101110;
    rom[49316] = 25'b0000000000011001100101101;
    rom[49317] = 25'b0000000000011001110101100;
    rom[49318] = 25'b0000000000011010000101010;
    rom[49319] = 25'b0000000000011010010101000;
    rom[49320] = 25'b0000000000011010100100110;
    rom[49321] = 25'b0000000000011010110100100;
    rom[49322] = 25'b0000000000011011000100010;
    rom[49323] = 25'b0000000000011011010100000;
    rom[49324] = 25'b0000000000011011100011110;
    rom[49325] = 25'b0000000000011011110011011;
    rom[49326] = 25'b0000000000011100000011001;
    rom[49327] = 25'b0000000000011100010010110;
    rom[49328] = 25'b0000000000011100100010100;
    rom[49329] = 25'b0000000000011100110010001;
    rom[49330] = 25'b0000000000011101000001111;
    rom[49331] = 25'b0000000000011101010001100;
    rom[49332] = 25'b0000000000011101100001001;
    rom[49333] = 25'b0000000000011101110000110;
    rom[49334] = 25'b0000000000011110000000011;
    rom[49335] = 25'b0000000000011110010000000;
    rom[49336] = 25'b0000000000011110011111100;
    rom[49337] = 25'b0000000000011110101111001;
    rom[49338] = 25'b0000000000011110111110110;
    rom[49339] = 25'b0000000000011111001110010;
    rom[49340] = 25'b0000000000011111011101111;
    rom[49341] = 25'b0000000000011111101101011;
    rom[49342] = 25'b0000000000011111111100111;
    rom[49343] = 25'b0000000000100000001100011;
    rom[49344] = 25'b0000000000100000011011111;
    rom[49345] = 25'b0000000000100000101011011;
    rom[49346] = 25'b0000000000100000111010111;
    rom[49347] = 25'b0000000000100001001010011;
    rom[49348] = 25'b0000000000100001011001110;
    rom[49349] = 25'b0000000000100001101001010;
    rom[49350] = 25'b0000000000100001111000101;
    rom[49351] = 25'b0000000000100010001000001;
    rom[49352] = 25'b0000000000100010010111100;
    rom[49353] = 25'b0000000000100010100110111;
    rom[49354] = 25'b0000000000100010110110010;
    rom[49355] = 25'b0000000000100011000101101;
    rom[49356] = 25'b0000000000100011010101000;
    rom[49357] = 25'b0000000000100011100100011;
    rom[49358] = 25'b0000000000100011110011101;
    rom[49359] = 25'b0000000000100100000011000;
    rom[49360] = 25'b0000000000100100010010010;
    rom[49361] = 25'b0000000000100100100001101;
    rom[49362] = 25'b0000000000100100110000111;
    rom[49363] = 25'b0000000000100101000000010;
    rom[49364] = 25'b0000000000100101001111100;
    rom[49365] = 25'b0000000000100101011110110;
    rom[49366] = 25'b0000000000100101101110000;
    rom[49367] = 25'b0000000000100101111101010;
    rom[49368] = 25'b0000000000100110001100011;
    rom[49369] = 25'b0000000000100110011011101;
    rom[49370] = 25'b0000000000100110101010111;
    rom[49371] = 25'b0000000000100110111010000;
    rom[49372] = 25'b0000000000100111001001010;
    rom[49373] = 25'b0000000000100111011000011;
    rom[49374] = 25'b0000000000100111100111101;
    rom[49375] = 25'b0000000000100111110110110;
    rom[49376] = 25'b0000000000101000000101111;
    rom[49377] = 25'b0000000000101000010101000;
    rom[49378] = 25'b0000000000101000100100000;
    rom[49379] = 25'b0000000000101000110011001;
    rom[49380] = 25'b0000000000101001000010001;
    rom[49381] = 25'b0000000000101001010001010;
    rom[49382] = 25'b0000000000101001100000011;
    rom[49383] = 25'b0000000000101001101111011;
    rom[49384] = 25'b0000000000101001111110011;
    rom[49385] = 25'b0000000000101010001101011;
    rom[49386] = 25'b0000000000101010011100100;
    rom[49387] = 25'b0000000000101010101011011;
    rom[49388] = 25'b0000000000101010111010100;
    rom[49389] = 25'b0000000000101011001001011;
    rom[49390] = 25'b0000000000101011011000011;
    rom[49391] = 25'b0000000000101011100111011;
    rom[49392] = 25'b0000000000101011110110010;
    rom[49393] = 25'b0000000000101100000101001;
    rom[49394] = 25'b0000000000101100010100001;
    rom[49395] = 25'b0000000000101100100011000;
    rom[49396] = 25'b0000000000101100110001111;
    rom[49397] = 25'b0000000000101101000000110;
    rom[49398] = 25'b0000000000101101001111101;
    rom[49399] = 25'b0000000000101101011110100;
    rom[49400] = 25'b0000000000101101101101010;
    rom[49401] = 25'b0000000000101101111100001;
    rom[49402] = 25'b0000000000101110001011000;
    rom[49403] = 25'b0000000000101110011001110;
    rom[49404] = 25'b0000000000101110101000101;
    rom[49405] = 25'b0000000000101110110111011;
    rom[49406] = 25'b0000000000101111000110001;
    rom[49407] = 25'b0000000000101111010100111;
    rom[49408] = 25'b0000000000101111100011101;
    rom[49409] = 25'b0000000000101111110010011;
    rom[49410] = 25'b0000000000110000000001000;
    rom[49411] = 25'b0000000000110000001111110;
    rom[49412] = 25'b0000000000110000011110100;
    rom[49413] = 25'b0000000000110000101101001;
    rom[49414] = 25'b0000000000110000111011111;
    rom[49415] = 25'b0000000000110001001010100;
    rom[49416] = 25'b0000000000110001011001001;
    rom[49417] = 25'b0000000000110001100111110;
    rom[49418] = 25'b0000000000110001110110011;
    rom[49419] = 25'b0000000000110010000101000;
    rom[49420] = 25'b0000000000110010010011100;
    rom[49421] = 25'b0000000000110010100010001;
    rom[49422] = 25'b0000000000110010110000101;
    rom[49423] = 25'b0000000000110010111111010;
    rom[49424] = 25'b0000000000110011001101111;
    rom[49425] = 25'b0000000000110011011100011;
    rom[49426] = 25'b0000000000110011101010111;
    rom[49427] = 25'b0000000000110011111001011;
    rom[49428] = 25'b0000000000110100000111111;
    rom[49429] = 25'b0000000000110100010110011;
    rom[49430] = 25'b0000000000110100100100111;
    rom[49431] = 25'b0000000000110100110011010;
    rom[49432] = 25'b0000000000110101000001110;
    rom[49433] = 25'b0000000000110101010000010;
    rom[49434] = 25'b0000000000110101011110101;
    rom[49435] = 25'b0000000000110101101101000;
    rom[49436] = 25'b0000000000110101111011011;
    rom[49437] = 25'b0000000000110110001001110;
    rom[49438] = 25'b0000000000110110011000001;
    rom[49439] = 25'b0000000000110110100110100;
    rom[49440] = 25'b0000000000110110110100111;
    rom[49441] = 25'b0000000000110111000011001;
    rom[49442] = 25'b0000000000110111010001100;
    rom[49443] = 25'b0000000000110111011111110;
    rom[49444] = 25'b0000000000110111101110000;
    rom[49445] = 25'b0000000000110111111100010;
    rom[49446] = 25'b0000000000111000001010101;
    rom[49447] = 25'b0000000000111000011000111;
    rom[49448] = 25'b0000000000111000100111001;
    rom[49449] = 25'b0000000000111000110101011;
    rom[49450] = 25'b0000000000111001000011100;
    rom[49451] = 25'b0000000000111001010001110;
    rom[49452] = 25'b0000000000111001100000000;
    rom[49453] = 25'b0000000000111001101110001;
    rom[49454] = 25'b0000000000111001111100010;
    rom[49455] = 25'b0000000000111010001010011;
    rom[49456] = 25'b0000000000111010011000100;
    rom[49457] = 25'b0000000000111010100110101;
    rom[49458] = 25'b0000000000111010110100110;
    rom[49459] = 25'b0000000000111011000010111;
    rom[49460] = 25'b0000000000111011010001000;
    rom[49461] = 25'b0000000000111011011111000;
    rom[49462] = 25'b0000000000111011101101000;
    rom[49463] = 25'b0000000000111011111011001;
    rom[49464] = 25'b0000000000111100001001001;
    rom[49465] = 25'b0000000000111100010111001;
    rom[49466] = 25'b0000000000111100100101001;
    rom[49467] = 25'b0000000000111100110011010;
    rom[49468] = 25'b0000000000111101000001010;
    rom[49469] = 25'b0000000000111101001111001;
    rom[49470] = 25'b0000000000111101011101001;
    rom[49471] = 25'b0000000000111101101011000;
    rom[49472] = 25'b0000000000111101111001000;
    rom[49473] = 25'b0000000000111110000110111;
    rom[49474] = 25'b0000000000111110010100110;
    rom[49475] = 25'b0000000000111110100010110;
    rom[49476] = 25'b0000000000111110110000100;
    rom[49477] = 25'b0000000000111110111110011;
    rom[49478] = 25'b0000000000111111001100010;
    rom[49479] = 25'b0000000000111111011010001;
    rom[49480] = 25'b0000000000111111100111111;
    rom[49481] = 25'b0000000000111111110101110;
    rom[49482] = 25'b0000000001000000000011100;
    rom[49483] = 25'b0000000001000000010001010;
    rom[49484] = 25'b0000000001000000011111001;
    rom[49485] = 25'b0000000001000000101100110;
    rom[49486] = 25'b0000000001000000111010100;
    rom[49487] = 25'b0000000001000001001000010;
    rom[49488] = 25'b0000000001000001010110000;
    rom[49489] = 25'b0000000001000001100011110;
    rom[49490] = 25'b0000000001000001110001011;
    rom[49491] = 25'b0000000001000001111111001;
    rom[49492] = 25'b0000000001000010001100110;
    rom[49493] = 25'b0000000001000010011010011;
    rom[49494] = 25'b0000000001000010101000000;
    rom[49495] = 25'b0000000001000010110101101;
    rom[49496] = 25'b0000000001000011000011010;
    rom[49497] = 25'b0000000001000011010000110;
    rom[49498] = 25'b0000000001000011011110011;
    rom[49499] = 25'b0000000001000011101100000;
    rom[49500] = 25'b0000000001000011111001100;
    rom[49501] = 25'b0000000001000100000111000;
    rom[49502] = 25'b0000000001000100010100101;
    rom[49503] = 25'b0000000001000100100010001;
    rom[49504] = 25'b0000000001000100101111101;
    rom[49505] = 25'b0000000001000100111101001;
    rom[49506] = 25'b0000000001000101001010101;
    rom[49507] = 25'b0000000001000101011000000;
    rom[49508] = 25'b0000000001000101100101100;
    rom[49509] = 25'b0000000001000101110010111;
    rom[49510] = 25'b0000000001000110000000011;
    rom[49511] = 25'b0000000001000110001101110;
    rom[49512] = 25'b0000000001000110011011001;
    rom[49513] = 25'b0000000001000110101000100;
    rom[49514] = 25'b0000000001000110110101111;
    rom[49515] = 25'b0000000001000111000011010;
    rom[49516] = 25'b0000000001000111010000101;
    rom[49517] = 25'b0000000001000111011101111;
    rom[49518] = 25'b0000000001000111101011010;
    rom[49519] = 25'b0000000001000111111000100;
    rom[49520] = 25'b0000000001001000000101111;
    rom[49521] = 25'b0000000001001000010011001;
    rom[49522] = 25'b0000000001001000100000011;
    rom[49523] = 25'b0000000001001000101101100;
    rom[49524] = 25'b0000000001001000111010110;
    rom[49525] = 25'b0000000001001001000111111;
    rom[49526] = 25'b0000000001001001010101010;
    rom[49527] = 25'b0000000001001001100010011;
    rom[49528] = 25'b0000000001001001101111100;
    rom[49529] = 25'b0000000001001001111100110;
    rom[49530] = 25'b0000000001001010001001111;
    rom[49531] = 25'b0000000001001010010111000;
    rom[49532] = 25'b0000000001001010100100001;
    rom[49533] = 25'b0000000001001010110001001;
    rom[49534] = 25'b0000000001001010111110010;
    rom[49535] = 25'b0000000001001011001011011;
    rom[49536] = 25'b0000000001001011011000011;
    rom[49537] = 25'b0000000001001011100101100;
    rom[49538] = 25'b0000000001001011110010100;
    rom[49539] = 25'b0000000001001011111111100;
    rom[49540] = 25'b0000000001001100001100100;
    rom[49541] = 25'b0000000001001100011001100;
    rom[49542] = 25'b0000000001001100100110100;
    rom[49543] = 25'b0000000001001100110011100;
    rom[49544] = 25'b0000000001001101000000011;
    rom[49545] = 25'b0000000001001101001101011;
    rom[49546] = 25'b0000000001001101011010010;
    rom[49547] = 25'b0000000001001101100111010;
    rom[49548] = 25'b0000000001001101110100001;
    rom[49549] = 25'b0000000001001110000001000;
    rom[49550] = 25'b0000000001001110001101110;
    rom[49551] = 25'b0000000001001110011010101;
    rom[49552] = 25'b0000000001001110100111100;
    rom[49553] = 25'b0000000001001110110100011;
    rom[49554] = 25'b0000000001001111000001001;
    rom[49555] = 25'b0000000001001111001101111;
    rom[49556] = 25'b0000000001001111011010110;
    rom[49557] = 25'b0000000001001111100111011;
    rom[49558] = 25'b0000000001001111110100010;
    rom[49559] = 25'b0000000001010000000000111;
    rom[49560] = 25'b0000000001010000001101110;
    rom[49561] = 25'b0000000001010000011010011;
    rom[49562] = 25'b0000000001010000100111001;
    rom[49563] = 25'b0000000001010000110011110;
    rom[49564] = 25'b0000000001010001000000011;
    rom[49565] = 25'b0000000001010001001101001;
    rom[49566] = 25'b0000000001010001011001110;
    rom[49567] = 25'b0000000001010001100110011;
    rom[49568] = 25'b0000000001010001110010111;
    rom[49569] = 25'b0000000001010001111111100;
    rom[49570] = 25'b0000000001010010001100001;
    rom[49571] = 25'b0000000001010010011000101;
    rom[49572] = 25'b0000000001010010100101010;
    rom[49573] = 25'b0000000001010010110001110;
    rom[49574] = 25'b0000000001010010111110010;
    rom[49575] = 25'b0000000001010011001010110;
    rom[49576] = 25'b0000000001010011010111011;
    rom[49577] = 25'b0000000001010011100011111;
    rom[49578] = 25'b0000000001010011110000010;
    rom[49579] = 25'b0000000001010011111100101;
    rom[49580] = 25'b0000000001010100001001010;
    rom[49581] = 25'b0000000001010100010101101;
    rom[49582] = 25'b0000000001010100100010000;
    rom[49583] = 25'b0000000001010100101110011;
    rom[49584] = 25'b0000000001010100111010110;
    rom[49585] = 25'b0000000001010101000111001;
    rom[49586] = 25'b0000000001010101010011011;
    rom[49587] = 25'b0000000001010101011111111;
    rom[49588] = 25'b0000000001010101101100001;
    rom[49589] = 25'b0000000001010101111000011;
    rom[49590] = 25'b0000000001010110000100110;
    rom[49591] = 25'b0000000001010110010001001;
    rom[49592] = 25'b0000000001010110011101010;
    rom[49593] = 25'b0000000001010110101001100;
    rom[49594] = 25'b0000000001010110110101110;
    rom[49595] = 25'b0000000001010111000010000;
    rom[49596] = 25'b0000000001010111001110010;
    rom[49597] = 25'b0000000001010111011010011;
    rom[49598] = 25'b0000000001010111100110101;
    rom[49599] = 25'b0000000001010111110010110;
    rom[49600] = 25'b0000000001010111111110111;
    rom[49601] = 25'b0000000001011000001011000;
    rom[49602] = 25'b0000000001011000010111001;
    rom[49603] = 25'b0000000001011000100011010;
    rom[49604] = 25'b0000000001011000101111011;
    rom[49605] = 25'b0000000001011000111011011;
    rom[49606] = 25'b0000000001011001000111100;
    rom[49607] = 25'b0000000001011001010011100;
    rom[49608] = 25'b0000000001011001011111100;
    rom[49609] = 25'b0000000001011001101011101;
    rom[49610] = 25'b0000000001011001110111100;
    rom[49611] = 25'b0000000001011010000011101;
    rom[49612] = 25'b0000000001011010001111100;
    rom[49613] = 25'b0000000001011010011011100;
    rom[49614] = 25'b0000000001011010100111100;
    rom[49615] = 25'b0000000001011010110011011;
    rom[49616] = 25'b0000000001011010111111010;
    rom[49617] = 25'b0000000001011011001011010;
    rom[49618] = 25'b0000000001011011010111001;
    rom[49619] = 25'b0000000001011011100011000;
    rom[49620] = 25'b0000000001011011101110110;
    rom[49621] = 25'b0000000001011011111010101;
    rom[49622] = 25'b0000000001011100000110011;
    rom[49623] = 25'b0000000001011100010010010;
    rom[49624] = 25'b0000000001011100011110000;
    rom[49625] = 25'b0000000001011100101001111;
    rom[49626] = 25'b0000000001011100110101101;
    rom[49627] = 25'b0000000001011101000001011;
    rom[49628] = 25'b0000000001011101001101001;
    rom[49629] = 25'b0000000001011101011000111;
    rom[49630] = 25'b0000000001011101100100101;
    rom[49631] = 25'b0000000001011101110000010;
    rom[49632] = 25'b0000000001011101111011111;
    rom[49633] = 25'b0000000001011110000111101;
    rom[49634] = 25'b0000000001011110010011010;
    rom[49635] = 25'b0000000001011110011110111;
    rom[49636] = 25'b0000000001011110101010100;
    rom[49637] = 25'b0000000001011110110110001;
    rom[49638] = 25'b0000000001011111000001101;
    rom[49639] = 25'b0000000001011111001101010;
    rom[49640] = 25'b0000000001011111011000111;
    rom[49641] = 25'b0000000001011111100100011;
    rom[49642] = 25'b0000000001011111101111111;
    rom[49643] = 25'b0000000001011111111011011;
    rom[49644] = 25'b0000000001100000000111000;
    rom[49645] = 25'b0000000001100000010010100;
    rom[49646] = 25'b0000000001100000011101111;
    rom[49647] = 25'b0000000001100000101001011;
    rom[49648] = 25'b0000000001100000110100111;
    rom[49649] = 25'b0000000001100001000000010;
    rom[49650] = 25'b0000000001100001001011101;
    rom[49651] = 25'b0000000001100001010111000;
    rom[49652] = 25'b0000000001100001100010011;
    rom[49653] = 25'b0000000001100001101101110;
    rom[49654] = 25'b0000000001100001111001001;
    rom[49655] = 25'b0000000001100010000100100;
    rom[49656] = 25'b0000000001100010001111110;
    rom[49657] = 25'b0000000001100010011011001;
    rom[49658] = 25'b0000000001100010100110011;
    rom[49659] = 25'b0000000001100010110001101;
    rom[49660] = 25'b0000000001100010111100111;
    rom[49661] = 25'b0000000001100011001000001;
    rom[49662] = 25'b0000000001100011010011011;
    rom[49663] = 25'b0000000001100011011110101;
    rom[49664] = 25'b0000000001100011101001110;
    rom[49665] = 25'b0000000001100011110101000;
    rom[49666] = 25'b0000000001100100000000001;
    rom[49667] = 25'b0000000001100100001011011;
    rom[49668] = 25'b0000000001100100010110100;
    rom[49669] = 25'b0000000001100100100001100;
    rom[49670] = 25'b0000000001100100101100101;
    rom[49671] = 25'b0000000001100100110111110;
    rom[49672] = 25'b0000000001100101000010110;
    rom[49673] = 25'b0000000001100101001101111;
    rom[49674] = 25'b0000000001100101011000111;
    rom[49675] = 25'b0000000001100101100100000;
    rom[49676] = 25'b0000000001100101101111000;
    rom[49677] = 25'b0000000001100101111010000;
    rom[49678] = 25'b0000000001100110000101000;
    rom[49679] = 25'b0000000001100110010000000;
    rom[49680] = 25'b0000000001100110011011000;
    rom[49681] = 25'b0000000001100110100101111;
    rom[49682] = 25'b0000000001100110110000110;
    rom[49683] = 25'b0000000001100110111011110;
    rom[49684] = 25'b0000000001100111000110101;
    rom[49685] = 25'b0000000001100111010001100;
    rom[49686] = 25'b0000000001100111011100011;
    rom[49687] = 25'b0000000001100111100111001;
    rom[49688] = 25'b0000000001100111110010000;
    rom[49689] = 25'b0000000001100111111100111;
    rom[49690] = 25'b0000000001101000000111101;
    rom[49691] = 25'b0000000001101000010010100;
    rom[49692] = 25'b0000000001101000011101010;
    rom[49693] = 25'b0000000001101000101000000;
    rom[49694] = 25'b0000000001101000110010110;
    rom[49695] = 25'b0000000001101000111101100;
    rom[49696] = 25'b0000000001101001001000010;
    rom[49697] = 25'b0000000001101001010010111;
    rom[49698] = 25'b0000000001101001011101101;
    rom[49699] = 25'b0000000001101001101000010;
    rom[49700] = 25'b0000000001101001110010111;
    rom[49701] = 25'b0000000001101001111101100;
    rom[49702] = 25'b0000000001101010001000001;
    rom[49703] = 25'b0000000001101010010010110;
    rom[49704] = 25'b0000000001101010011101011;
    rom[49705] = 25'b0000000001101010100111111;
    rom[49706] = 25'b0000000001101010110010100;
    rom[49707] = 25'b0000000001101010111101000;
    rom[49708] = 25'b0000000001101011000111101;
    rom[49709] = 25'b0000000001101011010010000;
    rom[49710] = 25'b0000000001101011011100101;
    rom[49711] = 25'b0000000001101011100111000;
    rom[49712] = 25'b0000000001101011110001100;
    rom[49713] = 25'b0000000001101011111100000;
    rom[49714] = 25'b0000000001101100000110011;
    rom[49715] = 25'b0000000001101100010000110;
    rom[49716] = 25'b0000000001101100011011010;
    rom[49717] = 25'b0000000001101100100101101;
    rom[49718] = 25'b0000000001101100110000000;
    rom[49719] = 25'b0000000001101100111010011;
    rom[49720] = 25'b0000000001101101000100110;
    rom[49721] = 25'b0000000001101101001111000;
    rom[49722] = 25'b0000000001101101011001011;
    rom[49723] = 25'b0000000001101101100011101;
    rom[49724] = 25'b0000000001101101101101111;
    rom[49725] = 25'b0000000001101101111000001;
    rom[49726] = 25'b0000000001101110000010100;
    rom[49727] = 25'b0000000001101110001100101;
    rom[49728] = 25'b0000000001101110010110111;
    rom[49729] = 25'b0000000001101110100001001;
    rom[49730] = 25'b0000000001101110101011010;
    rom[49731] = 25'b0000000001101110110101011;
    rom[49732] = 25'b0000000001101110111111101;
    rom[49733] = 25'b0000000001101111001001110;
    rom[49734] = 25'b0000000001101111010011111;
    rom[49735] = 25'b0000000001101111011110000;
    rom[49736] = 25'b0000000001101111101000000;
    rom[49737] = 25'b0000000001101111110010001;
    rom[49738] = 25'b0000000001101111111100010;
    rom[49739] = 25'b0000000001110000000110010;
    rom[49740] = 25'b0000000001110000010000010;
    rom[49741] = 25'b0000000001110000011010010;
    rom[49742] = 25'b0000000001110000100100010;
    rom[49743] = 25'b0000000001110000101110010;
    rom[49744] = 25'b0000000001110000111000010;
    rom[49745] = 25'b0000000001110001000010010;
    rom[49746] = 25'b0000000001110001001100001;
    rom[49747] = 25'b0000000001110001010110000;
    rom[49748] = 25'b0000000001110001100000000;
    rom[49749] = 25'b0000000001110001101001111;
    rom[49750] = 25'b0000000001110001110011110;
    rom[49751] = 25'b0000000001110001111101101;
    rom[49752] = 25'b0000000001110010000111100;
    rom[49753] = 25'b0000000001110010010001011;
    rom[49754] = 25'b0000000001110010011011001;
    rom[49755] = 25'b0000000001110010100101000;
    rom[49756] = 25'b0000000001110010101110101;
    rom[49757] = 25'b0000000001110010111000100;
    rom[49758] = 25'b0000000001110011000010010;
    rom[49759] = 25'b0000000001110011001100000;
    rom[49760] = 25'b0000000001110011010101110;
    rom[49761] = 25'b0000000001110011011111011;
    rom[49762] = 25'b0000000001110011101001000;
    rom[49763] = 25'b0000000001110011110010110;
    rom[49764] = 25'b0000000001110011111100011;
    rom[49765] = 25'b0000000001110100000110001;
    rom[49766] = 25'b0000000001110100001111110;
    rom[49767] = 25'b0000000001110100011001011;
    rom[49768] = 25'b0000000001110100100010111;
    rom[49769] = 25'b0000000001110100101100100;
    rom[49770] = 25'b0000000001110100110110000;
    rom[49771] = 25'b0000000001110100111111100;
    rom[49772] = 25'b0000000001110101001001001;
    rom[49773] = 25'b0000000001110101010010101;
    rom[49774] = 25'b0000000001110101011100001;
    rom[49775] = 25'b0000000001110101100101101;
    rom[49776] = 25'b0000000001110101101111000;
    rom[49777] = 25'b0000000001110101111000100;
    rom[49778] = 25'b0000000001110110000001111;
    rom[49779] = 25'b0000000001110110001011011;
    rom[49780] = 25'b0000000001110110010100110;
    rom[49781] = 25'b0000000001110110011110001;
    rom[49782] = 25'b0000000001110110100111100;
    rom[49783] = 25'b0000000001110110110000111;
    rom[49784] = 25'b0000000001110110111010010;
    rom[49785] = 25'b0000000001110111000011101;
    rom[49786] = 25'b0000000001110111001100111;
    rom[49787] = 25'b0000000001110111010110001;
    rom[49788] = 25'b0000000001110111011111100;
    rom[49789] = 25'b0000000001110111101000110;
    rom[49790] = 25'b0000000001110111110010000;
    rom[49791] = 25'b0000000001110111111011010;
    rom[49792] = 25'b0000000001111000000100011;
    rom[49793] = 25'b0000000001111000001101101;
    rom[49794] = 25'b0000000001111000010110110;
    rom[49795] = 25'b0000000001111000011111111;
    rom[49796] = 25'b0000000001111000101001001;
    rom[49797] = 25'b0000000001111000110010010;
    rom[49798] = 25'b0000000001111000111011011;
    rom[49799] = 25'b0000000001111001000100100;
    rom[49800] = 25'b0000000001111001001101101;
    rom[49801] = 25'b0000000001111001010110101;
    rom[49802] = 25'b0000000001111001011111110;
    rom[49803] = 25'b0000000001111001101000101;
    rom[49804] = 25'b0000000001111001110001110;
    rom[49805] = 25'b0000000001111001111010110;
    rom[49806] = 25'b0000000001111010000011110;
    rom[49807] = 25'b0000000001111010001100110;
    rom[49808] = 25'b0000000001111010010101110;
    rom[49809] = 25'b0000000001111010011110101;
    rom[49810] = 25'b0000000001111010100111100;
    rom[49811] = 25'b0000000001111010110000100;
    rom[49812] = 25'b0000000001111010111001011;
    rom[49813] = 25'b0000000001111011000010010;
    rom[49814] = 25'b0000000001111011001011001;
    rom[49815] = 25'b0000000001111011010100000;
    rom[49816] = 25'b0000000001111011011100110;
    rom[49817] = 25'b0000000001111011100101101;
    rom[49818] = 25'b0000000001111011101110011;
    rom[49819] = 25'b0000000001111011110111010;
    rom[49820] = 25'b0000000001111100000000000;
    rom[49821] = 25'b0000000001111100001000110;
    rom[49822] = 25'b0000000001111100010001011;
    rom[49823] = 25'b0000000001111100011010010;
    rom[49824] = 25'b0000000001111100100010111;
    rom[49825] = 25'b0000000001111100101011101;
    rom[49826] = 25'b0000000001111100110100010;
    rom[49827] = 25'b0000000001111100111101000;
    rom[49828] = 25'b0000000001111101000101100;
    rom[49829] = 25'b0000000001111101001110010;
    rom[49830] = 25'b0000000001111101010110111;
    rom[49831] = 25'b0000000001111101011111011;
    rom[49832] = 25'b0000000001111101101000000;
    rom[49833] = 25'b0000000001111101110000100;
    rom[49834] = 25'b0000000001111101111001001;
    rom[49835] = 25'b0000000001111110000001101;
    rom[49836] = 25'b0000000001111110001010001;
    rom[49837] = 25'b0000000001111110010010101;
    rom[49838] = 25'b0000000001111110011011001;
    rom[49839] = 25'b0000000001111110100011101;
    rom[49840] = 25'b0000000001111110101100000;
    rom[49841] = 25'b0000000001111110110100100;
    rom[49842] = 25'b0000000001111110111100111;
    rom[49843] = 25'b0000000001111111000101010;
    rom[49844] = 25'b0000000001111111001101101;
    rom[49845] = 25'b0000000001111111010110000;
    rom[49846] = 25'b0000000001111111011110011;
    rom[49847] = 25'b0000000001111111100110110;
    rom[49848] = 25'b0000000001111111101111000;
    rom[49849] = 25'b0000000001111111110111011;
    rom[49850] = 25'b0000000001111111111111101;
    rom[49851] = 25'b0000000010000000000111111;
    rom[49852] = 25'b0000000010000000010000010;
    rom[49853] = 25'b0000000010000000011000011;
    rom[49854] = 25'b0000000010000000100000101;
    rom[49855] = 25'b0000000010000000101000111;
    rom[49856] = 25'b0000000010000000110001000;
    rom[49857] = 25'b0000000010000000111001001;
    rom[49858] = 25'b0000000010000001000001010;
    rom[49859] = 25'b0000000010000001001001100;
    rom[49860] = 25'b0000000010000001010001101;
    rom[49861] = 25'b0000000010000001011001110;
    rom[49862] = 25'b0000000010000001100001110;
    rom[49863] = 25'b0000000010000001101001111;
    rom[49864] = 25'b0000000010000001110010000;
    rom[49865] = 25'b0000000010000001111010000;
    rom[49866] = 25'b0000000010000010000010000;
    rom[49867] = 25'b0000000010000010001010000;
    rom[49868] = 25'b0000000010000010010010001;
    rom[49869] = 25'b0000000010000010011010000;
    rom[49870] = 25'b0000000010000010100010000;
    rom[49871] = 25'b0000000010000010101010000;
    rom[49872] = 25'b0000000010000010110001111;
    rom[49873] = 25'b0000000010000010111001111;
    rom[49874] = 25'b0000000010000011000001110;
    rom[49875] = 25'b0000000010000011001001101;
    rom[49876] = 25'b0000000010000011010001100;
    rom[49877] = 25'b0000000010000011011001011;
    rom[49878] = 25'b0000000010000011100001010;
    rom[49879] = 25'b0000000010000011101001000;
    rom[49880] = 25'b0000000010000011110000110;
    rom[49881] = 25'b0000000010000011111000101;
    rom[49882] = 25'b0000000010000100000000011;
    rom[49883] = 25'b0000000010000100001000001;
    rom[49884] = 25'b0000000010000100001111111;
    rom[49885] = 25'b0000000010000100010111101;
    rom[49886] = 25'b0000000010000100011111010;
    rom[49887] = 25'b0000000010000100100111000;
    rom[49888] = 25'b0000000010000100101110110;
    rom[49889] = 25'b0000000010000100110110011;
    rom[49890] = 25'b0000000010000100111110000;
    rom[49891] = 25'b0000000010000101000101101;
    rom[49892] = 25'b0000000010000101001101010;
    rom[49893] = 25'b0000000010000101010100110;
    rom[49894] = 25'b0000000010000101011100011;
    rom[49895] = 25'b0000000010000101100011111;
    rom[49896] = 25'b0000000010000101101011100;
    rom[49897] = 25'b0000000010000101110011000;
    rom[49898] = 25'b0000000010000101111010100;
    rom[49899] = 25'b0000000010000110000010001;
    rom[49900] = 25'b0000000010000110001001101;
    rom[49901] = 25'b0000000010000110010001000;
    rom[49902] = 25'b0000000010000110011000011;
    rom[49903] = 25'b0000000010000110011111111;
    rom[49904] = 25'b0000000010000110100111011;
    rom[49905] = 25'b0000000010000110101110110;
    rom[49906] = 25'b0000000010000110110110001;
    rom[49907] = 25'b0000000010000110111101100;
    rom[49908] = 25'b0000000010000111000100111;
    rom[49909] = 25'b0000000010000111001100001;
    rom[49910] = 25'b0000000010000111010011100;
    rom[49911] = 25'b0000000010000111011010111;
    rom[49912] = 25'b0000000010000111100010001;
    rom[49913] = 25'b0000000010000111101001011;
    rom[49914] = 25'b0000000010000111110000101;
    rom[49915] = 25'b0000000010000111110111111;
    rom[49916] = 25'b0000000010000111111111000;
    rom[49917] = 25'b0000000010001000000110010;
    rom[49918] = 25'b0000000010001000001101011;
    rom[49919] = 25'b0000000010001000010100101;
    rom[49920] = 25'b0000000010001000011011110;
    rom[49921] = 25'b0000000010001000100010111;
    rom[49922] = 25'b0000000010001000101010001;
    rom[49923] = 25'b0000000010001000110001010;
    rom[49924] = 25'b0000000010001000111000010;
    rom[49925] = 25'b0000000010001000111111011;
    rom[49926] = 25'b0000000010001001000110011;
    rom[49927] = 25'b0000000010001001001101100;
    rom[49928] = 25'b0000000010001001010100100;
    rom[49929] = 25'b0000000010001001011011100;
    rom[49930] = 25'b0000000010001001100010100;
    rom[49931] = 25'b0000000010001001101001100;
    rom[49932] = 25'b0000000010001001110000011;
    rom[49933] = 25'b0000000010001001110111011;
    rom[49934] = 25'b0000000010001001111110011;
    rom[49935] = 25'b0000000010001010000101010;
    rom[49936] = 25'b0000000010001010001100001;
    rom[49937] = 25'b0000000010001010010011001;
    rom[49938] = 25'b0000000010001010011001111;
    rom[49939] = 25'b0000000010001010100000110;
    rom[49940] = 25'b0000000010001010100111101;
    rom[49941] = 25'b0000000010001010101110011;
    rom[49942] = 25'b0000000010001010110101010;
    rom[49943] = 25'b0000000010001010111100000;
    rom[49944] = 25'b0000000010001011000010110;
    rom[49945] = 25'b0000000010001011001001100;
    rom[49946] = 25'b0000000010001011010000010;
    rom[49947] = 25'b0000000010001011010111000;
    rom[49948] = 25'b0000000010001011011101101;
    rom[49949] = 25'b0000000010001011100100011;
    rom[49950] = 25'b0000000010001011101011000;
    rom[49951] = 25'b0000000010001011110001101;
    rom[49952] = 25'b0000000010001011111000010;
    rom[49953] = 25'b0000000010001011111110111;
    rom[49954] = 25'b0000000010001100000101100;
    rom[49955] = 25'b0000000010001100001100010;
    rom[49956] = 25'b0000000010001100010010110;
    rom[49957] = 25'b0000000010001100011001010;
    rom[49958] = 25'b0000000010001100011111110;
    rom[49959] = 25'b0000000010001100100110011;
    rom[49960] = 25'b0000000010001100101100111;
    rom[49961] = 25'b0000000010001100110011011;
    rom[49962] = 25'b0000000010001100111001111;
    rom[49963] = 25'b0000000010001101000000010;
    rom[49964] = 25'b0000000010001101000110110;
    rom[49965] = 25'b0000000010001101001101001;
    rom[49966] = 25'b0000000010001101010011101;
    rom[49967] = 25'b0000000010001101011010000;
    rom[49968] = 25'b0000000010001101100000011;
    rom[49969] = 25'b0000000010001101100110101;
    rom[49970] = 25'b0000000010001101101101000;
    rom[49971] = 25'b0000000010001101110011011;
    rom[49972] = 25'b0000000010001101111001110;
    rom[49973] = 25'b0000000010001110000000000;
    rom[49974] = 25'b0000000010001110000110011;
    rom[49975] = 25'b0000000010001110001100101;
    rom[49976] = 25'b0000000010001110010010111;
    rom[49977] = 25'b0000000010001110011001000;
    rom[49978] = 25'b0000000010001110011111010;
    rom[49979] = 25'b0000000010001110100101011;
    rom[49980] = 25'b0000000010001110101011110;
    rom[49981] = 25'b0000000010001110110001111;
    rom[49982] = 25'b0000000010001110111000000;
    rom[49983] = 25'b0000000010001110111110001;
    rom[49984] = 25'b0000000010001111000100010;
    rom[49985] = 25'b0000000010001111001010011;
    rom[49986] = 25'b0000000010001111010000011;
    rom[49987] = 25'b0000000010001111010110100;
    rom[49988] = 25'b0000000010001111011100100;
    rom[49989] = 25'b0000000010001111100010101;
    rom[49990] = 25'b0000000010001111101000101;
    rom[49991] = 25'b0000000010001111101110101;
    rom[49992] = 25'b0000000010001111110100101;
    rom[49993] = 25'b0000000010001111111010101;
    rom[49994] = 25'b0000000010010000000000101;
    rom[49995] = 25'b0000000010010000000110100;
    rom[49996] = 25'b0000000010010000001100100;
    rom[49997] = 25'b0000000010010000010010011;
    rom[49998] = 25'b0000000010010000011000010;
    rom[49999] = 25'b0000000010010000011110001;
    rom[50000] = 25'b0000000010010000100100000;
    rom[50001] = 25'b0000000010010000101001110;
    rom[50002] = 25'b0000000010010000101111101;
    rom[50003] = 25'b0000000010010000110101100;
    rom[50004] = 25'b0000000010010000111011010;
    rom[50005] = 25'b0000000010010001000001000;
    rom[50006] = 25'b0000000010010001000110110;
    rom[50007] = 25'b0000000010010001001100100;
    rom[50008] = 25'b0000000010010001010010010;
    rom[50009] = 25'b0000000010010001011000000;
    rom[50010] = 25'b0000000010010001011101110;
    rom[50011] = 25'b0000000010010001100011011;
    rom[50012] = 25'b0000000010010001101001000;
    rom[50013] = 25'b0000000010010001101110101;
    rom[50014] = 25'b0000000010010001110100010;
    rom[50015] = 25'b0000000010010001111001111;
    rom[50016] = 25'b0000000010010001111111100;
    rom[50017] = 25'b0000000010010010000101001;
    rom[50018] = 25'b0000000010010010001010110;
    rom[50019] = 25'b0000000010010010010000010;
    rom[50020] = 25'b0000000010010010010101111;
    rom[50021] = 25'b0000000010010010011011011;
    rom[50022] = 25'b0000000010010010100000111;
    rom[50023] = 25'b0000000010010010100110010;
    rom[50024] = 25'b0000000010010010101011110;
    rom[50025] = 25'b0000000010010010110001001;
    rom[50026] = 25'b0000000010010010110110101;
    rom[50027] = 25'b0000000010010010111100001;
    rom[50028] = 25'b0000000010010011000001100;
    rom[50029] = 25'b0000000010010011000110111;
    rom[50030] = 25'b0000000010010011001100010;
    rom[50031] = 25'b0000000010010011010001101;
    rom[50032] = 25'b0000000010010011010110111;
    rom[50033] = 25'b0000000010010011011100010;
    rom[50034] = 25'b0000000010010011100001100;
    rom[50035] = 25'b0000000010010011100110111;
    rom[50036] = 25'b0000000010010011101100010;
    rom[50037] = 25'b0000000010010011110001011;
    rom[50038] = 25'b0000000010010011110110101;
    rom[50039] = 25'b0000000010010011111011111;
    rom[50040] = 25'b0000000010010100000001001;
    rom[50041] = 25'b0000000010010100000110010;
    rom[50042] = 25'b0000000010010100001011100;
    rom[50043] = 25'b0000000010010100010000101;
    rom[50044] = 25'b0000000010010100010101110;
    rom[50045] = 25'b0000000010010100011010111;
    rom[50046] = 25'b0000000010010100100000000;
    rom[50047] = 25'b0000000010010100100101001;
    rom[50048] = 25'b0000000010010100101010010;
    rom[50049] = 25'b0000000010010100101111010;
    rom[50050] = 25'b0000000010010100110100010;
    rom[50051] = 25'b0000000010010100111001011;
    rom[50052] = 25'b0000000010010100111110011;
    rom[50053] = 25'b0000000010010101000011011;
    rom[50054] = 25'b0000000010010101001000011;
    rom[50055] = 25'b0000000010010101001101011;
    rom[50056] = 25'b0000000010010101010010010;
    rom[50057] = 25'b0000000010010101010111010;
    rom[50058] = 25'b0000000010010101011100001;
    rom[50059] = 25'b0000000010010101100001000;
    rom[50060] = 25'b0000000010010101100110000;
    rom[50061] = 25'b0000000010010101101010111;
    rom[50062] = 25'b0000000010010101101111101;
    rom[50063] = 25'b0000000010010101110100100;
    rom[50064] = 25'b0000000010010101111001010;
    rom[50065] = 25'b0000000010010101111110001;
    rom[50066] = 25'b0000000010010110000010111;
    rom[50067] = 25'b0000000010010110000111101;
    rom[50068] = 25'b0000000010010110001100100;
    rom[50069] = 25'b0000000010010110010001010;
    rom[50070] = 25'b0000000010010110010110000;
    rom[50071] = 25'b0000000010010110011010101;
    rom[50072] = 25'b0000000010010110011111011;
    rom[50073] = 25'b0000000010010110100100001;
    rom[50074] = 25'b0000000010010110101000110;
    rom[50075] = 25'b0000000010010110101101011;
    rom[50076] = 25'b0000000010010110110010000;
    rom[50077] = 25'b0000000010010110110110101;
    rom[50078] = 25'b0000000010010110111011010;
    rom[50079] = 25'b0000000010010110111111111;
    rom[50080] = 25'b0000000010010111000100011;
    rom[50081] = 25'b0000000010010111001000111;
    rom[50082] = 25'b0000000010010111001101100;
    rom[50083] = 25'b0000000010010111010001111;
    rom[50084] = 25'b0000000010010111010110100;
    rom[50085] = 25'b0000000010010111011011000;
    rom[50086] = 25'b0000000010010111011111011;
    rom[50087] = 25'b0000000010010111100011111;
    rom[50088] = 25'b0000000010010111101000011;
    rom[50089] = 25'b0000000010010111101100110;
    rom[50090] = 25'b0000000010010111110001001;
    rom[50091] = 25'b0000000010010111110101100;
    rom[50092] = 25'b0000000010010111111001111;
    rom[50093] = 25'b0000000010010111111110010;
    rom[50094] = 25'b0000000010011000000010101;
    rom[50095] = 25'b0000000010011000000111000;
    rom[50096] = 25'b0000000010011000001011010;
    rom[50097] = 25'b0000000010011000001111101;
    rom[50098] = 25'b0000000010011000010011110;
    rom[50099] = 25'b0000000010011000011000001;
    rom[50100] = 25'b0000000010011000011100011;
    rom[50101] = 25'b0000000010011000100000100;
    rom[50102] = 25'b0000000010011000100100110;
    rom[50103] = 25'b0000000010011000101001000;
    rom[50104] = 25'b0000000010011000101101001;
    rom[50105] = 25'b0000000010011000110001010;
    rom[50106] = 25'b0000000010011000110101100;
    rom[50107] = 25'b0000000010011000111001101;
    rom[50108] = 25'b0000000010011000111101110;
    rom[50109] = 25'b0000000010011001000001110;
    rom[50110] = 25'b0000000010011001000101111;
    rom[50111] = 25'b0000000010011001001001111;
    rom[50112] = 25'b0000000010011001001110000;
    rom[50113] = 25'b0000000010011001010010000;
    rom[50114] = 25'b0000000010011001010110001;
    rom[50115] = 25'b0000000010011001011010001;
    rom[50116] = 25'b0000000010011001011110001;
    rom[50117] = 25'b0000000010011001100010000;
    rom[50118] = 25'b0000000010011001100110000;
    rom[50119] = 25'b0000000010011001101010000;
    rom[50120] = 25'b0000000010011001101101111;
    rom[50121] = 25'b0000000010011001110001110;
    rom[50122] = 25'b0000000010011001110101101;
    rom[50123] = 25'b0000000010011001111001100;
    rom[50124] = 25'b0000000010011001111101011;
    rom[50125] = 25'b0000000010011010000001010;
    rom[50126] = 25'b0000000010011010000101000;
    rom[50127] = 25'b0000000010011010001000111;
    rom[50128] = 25'b0000000010011010001100110;
    rom[50129] = 25'b0000000010011010010000100;
    rom[50130] = 25'b0000000010011010010100010;
    rom[50131] = 25'b0000000010011010011000000;
    rom[50132] = 25'b0000000010011010011011110;
    rom[50133] = 25'b0000000010011010011111100;
    rom[50134] = 25'b0000000010011010100011001;
    rom[50135] = 25'b0000000010011010100110111;
    rom[50136] = 25'b0000000010011010101010100;
    rom[50137] = 25'b0000000010011010101110001;
    rom[50138] = 25'b0000000010011010110001110;
    rom[50139] = 25'b0000000010011010110101011;
    rom[50140] = 25'b0000000010011010111001000;
    rom[50141] = 25'b0000000010011010111100101;
    rom[50142] = 25'b0000000010011011000000001;
    rom[50143] = 25'b0000000010011011000011110;
    rom[50144] = 25'b0000000010011011000111010;
    rom[50145] = 25'b0000000010011011001010110;
    rom[50146] = 25'b0000000010011011001110011;
    rom[50147] = 25'b0000000010011011010001110;
    rom[50148] = 25'b0000000010011011010101010;
    rom[50149] = 25'b0000000010011011011000110;
    rom[50150] = 25'b0000000010011011011100001;
    rom[50151] = 25'b0000000010011011011111101;
    rom[50152] = 25'b0000000010011011100011001;
    rom[50153] = 25'b0000000010011011100110100;
    rom[50154] = 25'b0000000010011011101001110;
    rom[50155] = 25'b0000000010011011101101001;
    rom[50156] = 25'b0000000010011011110000100;
    rom[50157] = 25'b0000000010011011110011111;
    rom[50158] = 25'b0000000010011011110111001;
    rom[50159] = 25'b0000000010011011111010100;
    rom[50160] = 25'b0000000010011011111101110;
    rom[50161] = 25'b0000000010011100000001001;
    rom[50162] = 25'b0000000010011100000100011;
    rom[50163] = 25'b0000000010011100000111101;
    rom[50164] = 25'b0000000010011100001010110;
    rom[50165] = 25'b0000000010011100001110000;
    rom[50166] = 25'b0000000010011100010001010;
    rom[50167] = 25'b0000000010011100010100011;
    rom[50168] = 25'b0000000010011100010111101;
    rom[50169] = 25'b0000000010011100011010101;
    rom[50170] = 25'b0000000010011100011101111;
    rom[50171] = 25'b0000000010011100100000111;
    rom[50172] = 25'b0000000010011100100100000;
    rom[50173] = 25'b0000000010011100100111001;
    rom[50174] = 25'b0000000010011100101010001;
    rom[50175] = 25'b0000000010011100101101010;
    rom[50176] = 25'b0000000010011100110000011;
    rom[50177] = 25'b0000000010011100110011010;
    rom[50178] = 25'b0000000010011100110110010;
    rom[50179] = 25'b0000000010011100111001010;
    rom[50180] = 25'b0000000010011100111100010;
    rom[50181] = 25'b0000000010011100111111010;
    rom[50182] = 25'b0000000010011101000010001;
    rom[50183] = 25'b0000000010011101000101000;
    rom[50184] = 25'b0000000010011101001000000;
    rom[50185] = 25'b0000000010011101001010111;
    rom[50186] = 25'b0000000010011101001101110;
    rom[50187] = 25'b0000000010011101010000101;
    rom[50188] = 25'b0000000010011101010011011;
    rom[50189] = 25'b0000000010011101010110011;
    rom[50190] = 25'b0000000010011101011001001;
    rom[50191] = 25'b0000000010011101011011111;
    rom[50192] = 25'b0000000010011101011110110;
    rom[50193] = 25'b0000000010011101100001100;
    rom[50194] = 25'b0000000010011101100100010;
    rom[50195] = 25'b0000000010011101100111000;
    rom[50196] = 25'b0000000010011101101001101;
    rom[50197] = 25'b0000000010011101101100011;
    rom[50198] = 25'b0000000010011101101111001;
    rom[50199] = 25'b0000000010011101110001110;
    rom[50200] = 25'b0000000010011101110100011;
    rom[50201] = 25'b0000000010011101110111001;
    rom[50202] = 25'b0000000010011101111001110;
    rom[50203] = 25'b0000000010011101111100011;
    rom[50204] = 25'b0000000010011101111110111;
    rom[50205] = 25'b0000000010011110000001100;
    rom[50206] = 25'b0000000010011110000100001;
    rom[50207] = 25'b0000000010011110000110101;
    rom[50208] = 25'b0000000010011110001001001;
    rom[50209] = 25'b0000000010011110001011101;
    rom[50210] = 25'b0000000010011110001110001;
    rom[50211] = 25'b0000000010011110010000101;
    rom[50212] = 25'b0000000010011110010011001;
    rom[50213] = 25'b0000000010011110010101100;
    rom[50214] = 25'b0000000010011110011000000;
    rom[50215] = 25'b0000000010011110011010011;
    rom[50216] = 25'b0000000010011110011100111;
    rom[50217] = 25'b0000000010011110011111010;
    rom[50218] = 25'b0000000010011110100001101;
    rom[50219] = 25'b0000000010011110100011111;
    rom[50220] = 25'b0000000010011110100110011;
    rom[50221] = 25'b0000000010011110101000110;
    rom[50222] = 25'b0000000010011110101010111;
    rom[50223] = 25'b0000000010011110101101010;
    rom[50224] = 25'b0000000010011110101111100;
    rom[50225] = 25'b0000000010011110110001111;
    rom[50226] = 25'b0000000010011110110100001;
    rom[50227] = 25'b0000000010011110110110011;
    rom[50228] = 25'b0000000010011110111000101;
    rom[50229] = 25'b0000000010011110111010110;
    rom[50230] = 25'b0000000010011110111101000;
    rom[50231] = 25'b0000000010011110111111001;
    rom[50232] = 25'b0000000010011111000001010;
    rom[50233] = 25'b0000000010011111000011011;
    rom[50234] = 25'b0000000010011111000101100;
    rom[50235] = 25'b0000000010011111000111110;
    rom[50236] = 25'b0000000010011111001001110;
    rom[50237] = 25'b0000000010011111001011110;
    rom[50238] = 25'b0000000010011111001110000;
    rom[50239] = 25'b0000000010011111010000000;
    rom[50240] = 25'b0000000010011111010010000;
    rom[50241] = 25'b0000000010011111010100000;
    rom[50242] = 25'b0000000010011111010110000;
    rom[50243] = 25'b0000000010011111011000000;
    rom[50244] = 25'b0000000010011111011010000;
    rom[50245] = 25'b0000000010011111011100000;
    rom[50246] = 25'b0000000010011111011101111;
    rom[50247] = 25'b0000000010011111011111110;
    rom[50248] = 25'b0000000010011111100001110;
    rom[50249] = 25'b0000000010011111100011101;
    rom[50250] = 25'b0000000010011111100101100;
    rom[50251] = 25'b0000000010011111100111011;
    rom[50252] = 25'b0000000010011111101001010;
    rom[50253] = 25'b0000000010011111101011001;
    rom[50254] = 25'b0000000010011111101100111;
    rom[50255] = 25'b0000000010011111101110110;
    rom[50256] = 25'b0000000010011111110000100;
    rom[50257] = 25'b0000000010011111110010010;
    rom[50258] = 25'b0000000010011111110100000;
    rom[50259] = 25'b0000000010011111110101110;
    rom[50260] = 25'b0000000010011111110111100;
    rom[50261] = 25'b0000000010011111111001010;
    rom[50262] = 25'b0000000010011111111011000;
    rom[50263] = 25'b0000000010011111111100101;
    rom[50264] = 25'b0000000010011111111110010;
    rom[50265] = 25'b0000000010011111111111111;
    rom[50266] = 25'b0000000010100000000001101;
    rom[50267] = 25'b0000000010100000000011001;
    rom[50268] = 25'b0000000010100000000100110;
    rom[50269] = 25'b0000000010100000000110011;
    rom[50270] = 25'b0000000010100000001000000;
    rom[50271] = 25'b0000000010100000001001100;
    rom[50272] = 25'b0000000010100000001011000;
    rom[50273] = 25'b0000000010100000001100101;
    rom[50274] = 25'b0000000010100000001110001;
    rom[50275] = 25'b0000000010100000001111101;
    rom[50276] = 25'b0000000010100000010001001;
    rom[50277] = 25'b0000000010100000010010101;
    rom[50278] = 25'b0000000010100000010100000;
    rom[50279] = 25'b0000000010100000010101100;
    rom[50280] = 25'b0000000010100000010110111;
    rom[50281] = 25'b0000000010100000011000010;
    rom[50282] = 25'b0000000010100000011001110;
    rom[50283] = 25'b0000000010100000011011001;
    rom[50284] = 25'b0000000010100000011100011;
    rom[50285] = 25'b0000000010100000011101110;
    rom[50286] = 25'b0000000010100000011111001;
    rom[50287] = 25'b0000000010100000100000011;
    rom[50288] = 25'b0000000010100000100001110;
    rom[50289] = 25'b0000000010100000100011000;
    rom[50290] = 25'b0000000010100000100100011;
    rom[50291] = 25'b0000000010100000100101100;
    rom[50292] = 25'b0000000010100000100110110;
    rom[50293] = 25'b0000000010100000101000001;
    rom[50294] = 25'b0000000010100000101001010;
    rom[50295] = 25'b0000000010100000101010011;
    rom[50296] = 25'b0000000010100000101011101;
    rom[50297] = 25'b0000000010100000101100110;
    rom[50298] = 25'b0000000010100000101110000;
    rom[50299] = 25'b0000000010100000101111001;
    rom[50300] = 25'b0000000010100000110000010;
    rom[50301] = 25'b0000000010100000110001011;
    rom[50302] = 25'b0000000010100000110010100;
    rom[50303] = 25'b0000000010100000110011100;
    rom[50304] = 25'b0000000010100000110100100;
    rom[50305] = 25'b0000000010100000110101101;
    rom[50306] = 25'b0000000010100000110110101;
    rom[50307] = 25'b0000000010100000110111101;
    rom[50308] = 25'b0000000010100000111000101;
    rom[50309] = 25'b0000000010100000111001101;
    rom[50310] = 25'b0000000010100000111010101;
    rom[50311] = 25'b0000000010100000111011101;
    rom[50312] = 25'b0000000010100000111100100;
    rom[50313] = 25'b0000000010100000111101100;
    rom[50314] = 25'b0000000010100000111110010;
    rom[50315] = 25'b0000000010100000111111010;
    rom[50316] = 25'b0000000010100001000000001;
    rom[50317] = 25'b0000000010100001000001000;
    rom[50318] = 25'b0000000010100001000001111;
    rom[50319] = 25'b0000000010100001000010110;
    rom[50320] = 25'b0000000010100001000011100;
    rom[50321] = 25'b0000000010100001000100010;
    rom[50322] = 25'b0000000010100001000101001;
    rom[50323] = 25'b0000000010100001000101111;
    rom[50324] = 25'b0000000010100001000110101;
    rom[50325] = 25'b0000000010100001000111011;
    rom[50326] = 25'b0000000010100001001000001;
    rom[50327] = 25'b0000000010100001001000111;
    rom[50328] = 25'b0000000010100001001001100;
    rom[50329] = 25'b0000000010100001001010010;
    rom[50330] = 25'b0000000010100001001010111;
    rom[50331] = 25'b0000000010100001001011100;
    rom[50332] = 25'b0000000010100001001100010;
    rom[50333] = 25'b0000000010100001001100110;
    rom[50334] = 25'b0000000010100001001101011;
    rom[50335] = 25'b0000000010100001001110000;
    rom[50336] = 25'b0000000010100001001110101;
    rom[50337] = 25'b0000000010100001001111010;
    rom[50338] = 25'b0000000010100001001111110;
    rom[50339] = 25'b0000000010100001010000011;
    rom[50340] = 25'b0000000010100001010000110;
    rom[50341] = 25'b0000000010100001010001011;
    rom[50342] = 25'b0000000010100001010001111;
    rom[50343] = 25'b0000000010100001010010010;
    rom[50344] = 25'b0000000010100001010010110;
    rom[50345] = 25'b0000000010100001010011010;
    rom[50346] = 25'b0000000010100001010011101;
    rom[50347] = 25'b0000000010100001010100000;
    rom[50348] = 25'b0000000010100001010100011;
    rom[50349] = 25'b0000000010100001010100111;
    rom[50350] = 25'b0000000010100001010101010;
    rom[50351] = 25'b0000000010100001010101101;
    rom[50352] = 25'b0000000010100001010101111;
    rom[50353] = 25'b0000000010100001010110010;
    rom[50354] = 25'b0000000010100001010110101;
    rom[50355] = 25'b0000000010100001010111000;
    rom[50356] = 25'b0000000010100001010111010;
    rom[50357] = 25'b0000000010100001010111100;
    rom[50358] = 25'b0000000010100001010111110;
    rom[50359] = 25'b0000000010100001011000000;
    rom[50360] = 25'b0000000010100001011000010;
    rom[50361] = 25'b0000000010100001011000100;
    rom[50362] = 25'b0000000010100001011000101;
    rom[50363] = 25'b0000000010100001011000111;
    rom[50364] = 25'b0000000010100001011001000;
    rom[50365] = 25'b0000000010100001011001010;
    rom[50366] = 25'b0000000010100001011001010;
    rom[50367] = 25'b0000000010100001011001011;
    rom[50368] = 25'b0000000010100001011001101;
    rom[50369] = 25'b0000000010100001011001101;
    rom[50370] = 25'b0000000010100001011001110;
    rom[50371] = 25'b0000000010100001011001110;
    rom[50372] = 25'b0000000010100001011001111;
    rom[50373] = 25'b0000000010100001011001111;
    rom[50374] = 25'b0000000010100001011010000;
    rom[50375] = 25'b0000000010100001011010000;
    rom[50376] = 25'b0000000010100001011010000;
    rom[50377] = 25'b0000000010100001011010000;
    rom[50378] = 25'b0000000010100001011001111;
    rom[50379] = 25'b0000000010100001011001111;
    rom[50380] = 25'b0000000010100001011001110;
    rom[50381] = 25'b0000000010100001011001101;
    rom[50382] = 25'b0000000010100001011001101;
    rom[50383] = 25'b0000000010100001011001100;
    rom[50384] = 25'b0000000010100001011001011;
    rom[50385] = 25'b0000000010100001011001010;
    rom[50386] = 25'b0000000010100001011001001;
    rom[50387] = 25'b0000000010100001011000111;
    rom[50388] = 25'b0000000010100001011000111;
    rom[50389] = 25'b0000000010100001011000101;
    rom[50390] = 25'b0000000010100001011000011;
    rom[50391] = 25'b0000000010100001011000001;
    rom[50392] = 25'b0000000010100001011000000;
    rom[50393] = 25'b0000000010100001010111110;
    rom[50394] = 25'b0000000010100001010111011;
    rom[50395] = 25'b0000000010100001010111001;
    rom[50396] = 25'b0000000010100001010110111;
    rom[50397] = 25'b0000000010100001010110101;
    rom[50398] = 25'b0000000010100001010110010;
    rom[50399] = 25'b0000000010100001010101111;
    rom[50400] = 25'b0000000010100001010101100;
    rom[50401] = 25'b0000000010100001010101001;
    rom[50402] = 25'b0000000010100001010100110;
    rom[50403] = 25'b0000000010100001010100011;
    rom[50404] = 25'b0000000010100001010100000;
    rom[50405] = 25'b0000000010100001010011101;
    rom[50406] = 25'b0000000010100001010011010;
    rom[50407] = 25'b0000000010100001010010110;
    rom[50408] = 25'b0000000010100001010010010;
    rom[50409] = 25'b0000000010100001010001111;
    rom[50410] = 25'b0000000010100001010001011;
    rom[50411] = 25'b0000000010100001010000110;
    rom[50412] = 25'b0000000010100001010000011;
    rom[50413] = 25'b0000000010100001001111110;
    rom[50414] = 25'b0000000010100001001111010;
    rom[50415] = 25'b0000000010100001001110101;
    rom[50416] = 25'b0000000010100001001110001;
    rom[50417] = 25'b0000000010100001001101100;
    rom[50418] = 25'b0000000010100001001100111;
    rom[50419] = 25'b0000000010100001001100010;
    rom[50420] = 25'b0000000010100001001011101;
    rom[50421] = 25'b0000000010100001001011000;
    rom[50422] = 25'b0000000010100001001010011;
    rom[50423] = 25'b0000000010100001001001110;
    rom[50424] = 25'b0000000010100001001001000;
    rom[50425] = 25'b0000000010100001001000010;
    rom[50426] = 25'b0000000010100001000111100;
    rom[50427] = 25'b0000000010100001000110110;
    rom[50428] = 25'b0000000010100001000110000;
    rom[50429] = 25'b0000000010100001000101010;
    rom[50430] = 25'b0000000010100001000100100;
    rom[50431] = 25'b0000000010100001000011110;
    rom[50432] = 25'b0000000010100001000011000;
    rom[50433] = 25'b0000000010100001000010001;
    rom[50434] = 25'b0000000010100001000001010;
    rom[50435] = 25'b0000000010100001000000100;
    rom[50436] = 25'b0000000010100000111111101;
    rom[50437] = 25'b0000000010100000111110110;
    rom[50438] = 25'b0000000010100000111101111;
    rom[50439] = 25'b0000000010100000111101000;
    rom[50440] = 25'b0000000010100000111100000;
    rom[50441] = 25'b0000000010100000111011001;
    rom[50442] = 25'b0000000010100000111010010;
    rom[50443] = 25'b0000000010100000111001010;
    rom[50444] = 25'b0000000010100000111000011;
    rom[50445] = 25'b0000000010100000110111010;
    rom[50446] = 25'b0000000010100000110110010;
    rom[50447] = 25'b0000000010100000110101011;
    rom[50448] = 25'b0000000010100000110100010;
    rom[50449] = 25'b0000000010100000110011001;
    rom[50450] = 25'b0000000010100000110010001;
    rom[50451] = 25'b0000000010100000110001001;
    rom[50452] = 25'b0000000010100000110000000;
    rom[50453] = 25'b0000000010100000101111000;
    rom[50454] = 25'b0000000010100000101101111;
    rom[50455] = 25'b0000000010100000101100110;
    rom[50456] = 25'b0000000010100000101011101;
    rom[50457] = 25'b0000000010100000101010011;
    rom[50458] = 25'b0000000010100000101001010;
    rom[50459] = 25'b0000000010100000101000001;
    rom[50460] = 25'b0000000010100000100111000;
    rom[50461] = 25'b0000000010100000100101110;
    rom[50462] = 25'b0000000010100000100100100;
    rom[50463] = 25'b0000000010100000100011010;
    rom[50464] = 25'b0000000010100000100010000;
    rom[50465] = 25'b0000000010100000100000110;
    rom[50466] = 25'b0000000010100000011111100;
    rom[50467] = 25'b0000000010100000011110001;
    rom[50468] = 25'b0000000010100000011100111;
    rom[50469] = 25'b0000000010100000011011100;
    rom[50470] = 25'b0000000010100000011010010;
    rom[50471] = 25'b0000000010100000011001000;
    rom[50472] = 25'b0000000010100000010111100;
    rom[50473] = 25'b0000000010100000010110010;
    rom[50474] = 25'b0000000010100000010100111;
    rom[50475] = 25'b0000000010100000010011011;
    rom[50476] = 25'b0000000010100000010010000;
    rom[50477] = 25'b0000000010100000010000101;
    rom[50478] = 25'b0000000010100000001111001;
    rom[50479] = 25'b0000000010100000001101110;
    rom[50480] = 25'b0000000010100000001100010;
    rom[50481] = 25'b0000000010100000001010110;
    rom[50482] = 25'b0000000010100000001001011;
    rom[50483] = 25'b0000000010100000000111110;
    rom[50484] = 25'b0000000010100000000110010;
    rom[50485] = 25'b0000000010100000000100110;
    rom[50486] = 25'b0000000010100000000011001;
    rom[50487] = 25'b0000000010100000000001110;
    rom[50488] = 25'b0000000010100000000000001;
    rom[50489] = 25'b0000000010011111111110100;
    rom[50490] = 25'b0000000010011111111100111;
    rom[50491] = 25'b0000000010011111111011011;
    rom[50492] = 25'b0000000010011111111001101;
    rom[50493] = 25'b0000000010011111111000001;
    rom[50494] = 25'b0000000010011111110110011;
    rom[50495] = 25'b0000000010011111110100110;
    rom[50496] = 25'b0000000010011111110011000;
    rom[50497] = 25'b0000000010011111110001011;
    rom[50498] = 25'b0000000010011111101111101;
    rom[50499] = 25'b0000000010011111101101111;
    rom[50500] = 25'b0000000010011111101100010;
    rom[50501] = 25'b0000000010011111101010100;
    rom[50502] = 25'b0000000010011111101000101;
    rom[50503] = 25'b0000000010011111100110111;
    rom[50504] = 25'b0000000010011111100101001;
    rom[50505] = 25'b0000000010011111100011011;
    rom[50506] = 25'b0000000010011111100001101;
    rom[50507] = 25'b0000000010011111011111110;
    rom[50508] = 25'b0000000010011111011101111;
    rom[50509] = 25'b0000000010011111011100000;
    rom[50510] = 25'b0000000010011111011010010;
    rom[50511] = 25'b0000000010011111011000011;
    rom[50512] = 25'b0000000010011111010110011;
    rom[50513] = 25'b0000000010011111010100100;
    rom[50514] = 25'b0000000010011111010010100;
    rom[50515] = 25'b0000000010011111010000101;
    rom[50516] = 25'b0000000010011111001110110;
    rom[50517] = 25'b0000000010011111001100110;
    rom[50518] = 25'b0000000010011111001010110;
    rom[50519] = 25'b0000000010011111001000111;
    rom[50520] = 25'b0000000010011111000110110;
    rom[50521] = 25'b0000000010011111000100110;
    rom[50522] = 25'b0000000010011111000010110;
    rom[50523] = 25'b0000000010011111000000110;
    rom[50524] = 25'b0000000010011110111110101;
    rom[50525] = 25'b0000000010011110111100101;
    rom[50526] = 25'b0000000010011110111010100;
    rom[50527] = 25'b0000000010011110111000100;
    rom[50528] = 25'b0000000010011110110110011;
    rom[50529] = 25'b0000000010011110110100010;
    rom[50530] = 25'b0000000010011110110010001;
    rom[50531] = 25'b0000000010011110110000000;
    rom[50532] = 25'b0000000010011110101101111;
    rom[50533] = 25'b0000000010011110101011101;
    rom[50534] = 25'b0000000010011110101001100;
    rom[50535] = 25'b0000000010011110100111010;
    rom[50536] = 25'b0000000010011110100101000;
    rom[50537] = 25'b0000000010011110100010110;
    rom[50538] = 25'b0000000010011110100000101;
    rom[50539] = 25'b0000000010011110011110011;
    rom[50540] = 25'b0000000010011110011100001;
    rom[50541] = 25'b0000000010011110011001111;
    rom[50542] = 25'b0000000010011110010111101;
    rom[50543] = 25'b0000000010011110010101010;
    rom[50544] = 25'b0000000010011110010010111;
    rom[50545] = 25'b0000000010011110010000101;
    rom[50546] = 25'b0000000010011110001110010;
    rom[50547] = 25'b0000000010011110001011111;
    rom[50548] = 25'b0000000010011110001001101;
    rom[50549] = 25'b0000000010011110000111010;
    rom[50550] = 25'b0000000010011110000100111;
    rom[50551] = 25'b0000000010011110000010011;
    rom[50552] = 25'b0000000010011110000000000;
    rom[50553] = 25'b0000000010011101111101100;
    rom[50554] = 25'b0000000010011101111011001;
    rom[50555] = 25'b0000000010011101111000110;
    rom[50556] = 25'b0000000010011101110110010;
    rom[50557] = 25'b0000000010011101110011110;
    rom[50558] = 25'b0000000010011101110001011;
    rom[50559] = 25'b0000000010011101101110110;
    rom[50560] = 25'b0000000010011101101100010;
    rom[50561] = 25'b0000000010011101101001110;
    rom[50562] = 25'b0000000010011101100111010;
    rom[50563] = 25'b0000000010011101100100101;
    rom[50564] = 25'b0000000010011101100010001;
    rom[50565] = 25'b0000000010011101011111100;
    rom[50566] = 25'b0000000010011101011100111;
    rom[50567] = 25'b0000000010011101011010011;
    rom[50568] = 25'b0000000010011101010111110;
    rom[50569] = 25'b0000000010011101010101000;
    rom[50570] = 25'b0000000010011101010010011;
    rom[50571] = 25'b0000000010011101001111110;
    rom[50572] = 25'b0000000010011101001101001;
    rom[50573] = 25'b0000000010011101001010100;
    rom[50574] = 25'b0000000010011101000111110;
    rom[50575] = 25'b0000000010011101000101000;
    rom[50576] = 25'b0000000010011101000010011;
    rom[50577] = 25'b0000000010011100111111100;
    rom[50578] = 25'b0000000010011100111100111;
    rom[50579] = 25'b0000000010011100111010001;
    rom[50580] = 25'b0000000010011100110111011;
    rom[50581] = 25'b0000000010011100110100100;
    rom[50582] = 25'b0000000010011100110001110;
    rom[50583] = 25'b0000000010011100101110111;
    rom[50584] = 25'b0000000010011100101100001;
    rom[50585] = 25'b0000000010011100101001011;
    rom[50586] = 25'b0000000010011100100110011;
    rom[50587] = 25'b0000000010011100100011101;
    rom[50588] = 25'b0000000010011100100000110;
    rom[50589] = 25'b0000000010011100011101111;
    rom[50590] = 25'b0000000010011100011010111;
    rom[50591] = 25'b0000000010011100011000000;
    rom[50592] = 25'b0000000010011100010101001;
    rom[50593] = 25'b0000000010011100010010010;
    rom[50594] = 25'b0000000010011100001111010;
    rom[50595] = 25'b0000000010011100001100010;
    rom[50596] = 25'b0000000010011100001001011;
    rom[50597] = 25'b0000000010011100000110011;
    rom[50598] = 25'b0000000010011100000011011;
    rom[50599] = 25'b0000000010011100000000011;
    rom[50600] = 25'b0000000010011011111101011;
    rom[50601] = 25'b0000000010011011111010011;
    rom[50602] = 25'b0000000010011011110111010;
    rom[50603] = 25'b0000000010011011110100010;
    rom[50604] = 25'b0000000010011011110001010;
    rom[50605] = 25'b0000000010011011101110001;
    rom[50606] = 25'b0000000010011011101011000;
    rom[50607] = 25'b0000000010011011101000000;
    rom[50608] = 25'b0000000010011011100100110;
    rom[50609] = 25'b0000000010011011100001101;
    rom[50610] = 25'b0000000010011011011110100;
    rom[50611] = 25'b0000000010011011011011011;
    rom[50612] = 25'b0000000010011011011000010;
    rom[50613] = 25'b0000000010011011010101001;
    rom[50614] = 25'b0000000010011011010001111;
    rom[50615] = 25'b0000000010011011001110101;
    rom[50616] = 25'b0000000010011011001011100;
    rom[50617] = 25'b0000000010011011001000010;
    rom[50618] = 25'b0000000010011011000101000;
    rom[50619] = 25'b0000000010011011000001110;
    rom[50620] = 25'b0000000010011010111110100;
    rom[50621] = 25'b0000000010011010111011010;
    rom[50622] = 25'b0000000010011010111000000;
    rom[50623] = 25'b0000000010011010110100101;
    rom[50624] = 25'b0000000010011010110001010;
    rom[50625] = 25'b0000000010011010101110000;
    rom[50626] = 25'b0000000010011010101010101;
    rom[50627] = 25'b0000000010011010100111011;
    rom[50628] = 25'b0000000010011010100100000;
    rom[50629] = 25'b0000000010011010100000101;
    rom[50630] = 25'b0000000010011010011101010;
    rom[50631] = 25'b0000000010011010011001111;
    rom[50632] = 25'b0000000010011010010110011;
    rom[50633] = 25'b0000000010011010010011000;
    rom[50634] = 25'b0000000010011010001111101;
    rom[50635] = 25'b0000000010011010001100001;
    rom[50636] = 25'b0000000010011010001000110;
    rom[50637] = 25'b0000000010011010000101010;
    rom[50638] = 25'b0000000010011010000001110;
    rom[50639] = 25'b0000000010011001111110011;
    rom[50640] = 25'b0000000010011001111010110;
    rom[50641] = 25'b0000000010011001110111011;
    rom[50642] = 25'b0000000010011001110011110;
    rom[50643] = 25'b0000000010011001110000010;
    rom[50644] = 25'b0000000010011001101100101;
    rom[50645] = 25'b0000000010011001101001001;
    rom[50646] = 25'b0000000010011001100101101;
    rom[50647] = 25'b0000000010011001100001111;
    rom[50648] = 25'b0000000010011001011110011;
    rom[50649] = 25'b0000000010011001011010110;
    rom[50650] = 25'b0000000010011001010111010;
    rom[50651] = 25'b0000000010011001010011100;
    rom[50652] = 25'b0000000010011001001111111;
    rom[50653] = 25'b0000000010011001001100010;
    rom[50654] = 25'b0000000010011001001000101;
    rom[50655] = 25'b0000000010011001000100111;
    rom[50656] = 25'b0000000010011001000001010;
    rom[50657] = 25'b0000000010011000111101100;
    rom[50658] = 25'b0000000010011000111001110;
    rom[50659] = 25'b0000000010011000110110001;
    rom[50660] = 25'b0000000010011000110010011;
    rom[50661] = 25'b0000000010011000101110101;
    rom[50662] = 25'b0000000010011000101010111;
    rom[50663] = 25'b0000000010011000100111001;
    rom[50664] = 25'b0000000010011000100011010;
    rom[50665] = 25'b0000000010011000011111100;
    rom[50666] = 25'b0000000010011000011011110;
    rom[50667] = 25'b0000000010011000010111111;
    rom[50668] = 25'b0000000010011000010100000;
    rom[50669] = 25'b0000000010011000010000010;
    rom[50670] = 25'b0000000010011000001100011;
    rom[50671] = 25'b0000000010011000001000100;
    rom[50672] = 25'b0000000010011000000100101;
    rom[50673] = 25'b0000000010011000000000110;
    rom[50674] = 25'b0000000010010111111100111;
    rom[50675] = 25'b0000000010010111111001000;
    rom[50676] = 25'b0000000010010111110101000;
    rom[50677] = 25'b0000000010010111110001001;
    rom[50678] = 25'b0000000010010111101101010;
    rom[50679] = 25'b0000000010010111101001010;
    rom[50680] = 25'b0000000010010111100101010;
    rom[50681] = 25'b0000000010010111100001011;
    rom[50682] = 25'b0000000010010111011101011;
    rom[50683] = 25'b0000000010010111011001010;
    rom[50684] = 25'b0000000010010111010101010;
    rom[50685] = 25'b0000000010010111010001010;
    rom[50686] = 25'b0000000010010111001101010;
    rom[50687] = 25'b0000000010010111001001010;
    rom[50688] = 25'b0000000010010111000101001;
    rom[50689] = 25'b0000000010010111000001001;
    rom[50690] = 25'b0000000010010110111101000;
    rom[50691] = 25'b0000000010010110111001000;
    rom[50692] = 25'b0000000010010110110100111;
    rom[50693] = 25'b0000000010010110110000110;
    rom[50694] = 25'b0000000010010110101100101;
    rom[50695] = 25'b0000000010010110101000100;
    rom[50696] = 25'b0000000010010110100100011;
    rom[50697] = 25'b0000000010010110100000001;
    rom[50698] = 25'b0000000010010110011100000;
    rom[50699] = 25'b0000000010010110010111111;
    rom[50700] = 25'b0000000010010110010011101;
    rom[50701] = 25'b0000000010010110001111100;
    rom[50702] = 25'b0000000010010110001011010;
    rom[50703] = 25'b0000000010010110000111000;
    rom[50704] = 25'b0000000010010110000010111;
    rom[50705] = 25'b0000000010010101111110100;
    rom[50706] = 25'b0000000010010101111010011;
    rom[50707] = 25'b0000000010010101110110000;
    rom[50708] = 25'b0000000010010101110001110;
    rom[50709] = 25'b0000000010010101101101100;
    rom[50710] = 25'b0000000010010101101001001;
    rom[50711] = 25'b0000000010010101100100111;
    rom[50712] = 25'b0000000010010101100000100;
    rom[50713] = 25'b0000000010010101011100010;
    rom[50714] = 25'b0000000010010101010111111;
    rom[50715] = 25'b0000000010010101010011101;
    rom[50716] = 25'b0000000010010101001111010;
    rom[50717] = 25'b0000000010010101001010110;
    rom[50718] = 25'b0000000010010101000110011;
    rom[50719] = 25'b0000000010010101000010000;
    rom[50720] = 25'b0000000010010100111101101;
    rom[50721] = 25'b0000000010010100111001001;
    rom[50722] = 25'b0000000010010100110100110;
    rom[50723] = 25'b0000000010010100110000010;
    rom[50724] = 25'b0000000010010100101011111;
    rom[50725] = 25'b0000000010010100100111011;
    rom[50726] = 25'b0000000010010100100010111;
    rom[50727] = 25'b0000000010010100011110100;
    rom[50728] = 25'b0000000010010100011010000;
    rom[50729] = 25'b0000000010010100010101100;
    rom[50730] = 25'b0000000010010100010000111;
    rom[50731] = 25'b0000000010010100001100011;
    rom[50732] = 25'b0000000010010100000111111;
    rom[50733] = 25'b0000000010010100000011011;
    rom[50734] = 25'b0000000010010011111110110;
    rom[50735] = 25'b0000000010010011111010010;
    rom[50736] = 25'b0000000010010011110101101;
    rom[50737] = 25'b0000000010010011110001000;
    rom[50738] = 25'b0000000010010011101100011;
    rom[50739] = 25'b0000000010010011100111110;
    rom[50740] = 25'b0000000010010011100011010;
    rom[50741] = 25'b0000000010010011011110101;
    rom[50742] = 25'b0000000010010011011001111;
    rom[50743] = 25'b0000000010010011010101010;
    rom[50744] = 25'b0000000010010011010000100;
    rom[50745] = 25'b0000000010010011001011111;
    rom[50746] = 25'b0000000010010011000111010;
    rom[50747] = 25'b0000000010010011000010100;
    rom[50748] = 25'b0000000010010010111101111;
    rom[50749] = 25'b0000000010010010111001001;
    rom[50750] = 25'b0000000010010010110100011;
    rom[50751] = 25'b0000000010010010101111101;
    rom[50752] = 25'b0000000010010010101010111;
    rom[50753] = 25'b0000000010010010100110001;
    rom[50754] = 25'b0000000010010010100001011;
    rom[50755] = 25'b0000000010010010011100101;
    rom[50756] = 25'b0000000010010010010111110;
    rom[50757] = 25'b0000000010010010010011000;
    rom[50758] = 25'b0000000010010010001110001;
    rom[50759] = 25'b0000000010010010001001011;
    rom[50760] = 25'b0000000010010010000100100;
    rom[50761] = 25'b0000000010010001111111101;
    rom[50762] = 25'b0000000010010001111010111;
    rom[50763] = 25'b0000000010010001110110000;
    rom[50764] = 25'b0000000010010001110001001;
    rom[50765] = 25'b0000000010010001101100010;
    rom[50766] = 25'b0000000010010001100111010;
    rom[50767] = 25'b0000000010010001100010100;
    rom[50768] = 25'b0000000010010001011101100;
    rom[50769] = 25'b0000000010010001011000100;
    rom[50770] = 25'b0000000010010001010011101;
    rom[50771] = 25'b0000000010010001001110110;
    rom[50772] = 25'b0000000010010001001001110;
    rom[50773] = 25'b0000000010010001000100110;
    rom[50774] = 25'b0000000010010000111111110;
    rom[50775] = 25'b0000000010010000111010111;
    rom[50776] = 25'b0000000010010000110101111;
    rom[50777] = 25'b0000000010010000110000110;
    rom[50778] = 25'b0000000010010000101011111;
    rom[50779] = 25'b0000000010010000100110110;
    rom[50780] = 25'b0000000010010000100001110;
    rom[50781] = 25'b0000000010010000011100110;
    rom[50782] = 25'b0000000010010000010111101;
    rom[50783] = 25'b0000000010010000010010101;
    rom[50784] = 25'b0000000010010000001101100;
    rom[50785] = 25'b0000000010010000001000011;
    rom[50786] = 25'b0000000010010000000011010;
    rom[50787] = 25'b0000000010001111111110001;
    rom[50788] = 25'b0000000010001111111001001;
    rom[50789] = 25'b0000000010001111110100000;
    rom[50790] = 25'b0000000010001111101110111;
    rom[50791] = 25'b0000000010001111101001110;
    rom[50792] = 25'b0000000010001111100100100;
    rom[50793] = 25'b0000000010001111011111011;
    rom[50794] = 25'b0000000010001111011010010;
    rom[50795] = 25'b0000000010001111010101000;
    rom[50796] = 25'b0000000010001111001111110;
    rom[50797] = 25'b0000000010001111001010101;
    rom[50798] = 25'b0000000010001111000101011;
    rom[50799] = 25'b0000000010001111000000001;
    rom[50800] = 25'b0000000010001110111010111;
    rom[50801] = 25'b0000000010001110110101101;
    rom[50802] = 25'b0000000010001110110000011;
    rom[50803] = 25'b0000000010001110101011001;
    rom[50804] = 25'b0000000010001110100101110;
    rom[50805] = 25'b0000000010001110100000101;
    rom[50806] = 25'b0000000010001110011011010;
    rom[50807] = 25'b0000000010001110010101111;
    rom[50808] = 25'b0000000010001110010000101;
    rom[50809] = 25'b0000000010001110001011010;
    rom[50810] = 25'b0000000010001110000110000;
    rom[50811] = 25'b0000000010001110000000101;
    rom[50812] = 25'b0000000010001101111011011;
    rom[50813] = 25'b0000000010001101110101111;
    rom[50814] = 25'b0000000010001101110000101;
    rom[50815] = 25'b0000000010001101101011001;
    rom[50816] = 25'b0000000010001101100101110;
    rom[50817] = 25'b0000000010001101100000011;
    rom[50818] = 25'b0000000010001101011010111;
    rom[50819] = 25'b0000000010001101010101100;
    rom[50820] = 25'b0000000010001101010000001;
    rom[50821] = 25'b0000000010001101001010101;
    rom[50822] = 25'b0000000010001101000101010;
    rom[50823] = 25'b0000000010001100111111110;
    rom[50824] = 25'b0000000010001100111010010;
    rom[50825] = 25'b0000000010001100110100110;
    rom[50826] = 25'b0000000010001100101111010;
    rom[50827] = 25'b0000000010001100101001110;
    rom[50828] = 25'b0000000010001100100100010;
    rom[50829] = 25'b0000000010001100011110110;
    rom[50830] = 25'b0000000010001100011001010;
    rom[50831] = 25'b0000000010001100010011110;
    rom[50832] = 25'b0000000010001100001110001;
    rom[50833] = 25'b0000000010001100001000101;
    rom[50834] = 25'b0000000010001100000011000;
    rom[50835] = 25'b0000000010001011111101100;
    rom[50836] = 25'b0000000010001011110111111;
    rom[50837] = 25'b0000000010001011110010011;
    rom[50838] = 25'b0000000010001011101100110;
    rom[50839] = 25'b0000000010001011100111001;
    rom[50840] = 25'b0000000010001011100001100;
    rom[50841] = 25'b0000000010001011011011111;
    rom[50842] = 25'b0000000010001011010110010;
    rom[50843] = 25'b0000000010001011010000100;
    rom[50844] = 25'b0000000010001011001010111;
    rom[50845] = 25'b0000000010001011000101010;
    rom[50846] = 25'b0000000010001010111111100;
    rom[50847] = 25'b0000000010001010111001111;
    rom[50848] = 25'b0000000010001010110100010;
    rom[50849] = 25'b0000000010001010101110011;
    rom[50850] = 25'b0000000010001010101000110;
    rom[50851] = 25'b0000000010001010100011000;
    rom[50852] = 25'b0000000010001010011101011;
    rom[50853] = 25'b0000000010001010010111100;
    rom[50854] = 25'b0000000010001010010001111;
    rom[50855] = 25'b0000000010001010001100000;
    rom[50856] = 25'b0000000010001010000110010;
    rom[50857] = 25'b0000000010001010000000100;
    rom[50858] = 25'b0000000010001001111010110;
    rom[50859] = 25'b0000000010001001110100111;
    rom[50860] = 25'b0000000010001001101111001;
    rom[50861] = 25'b0000000010001001101001011;
    rom[50862] = 25'b0000000010001001100011100;
    rom[50863] = 25'b0000000010001001011101101;
    rom[50864] = 25'b0000000010001001010111111;
    rom[50865] = 25'b0000000010001001010010000;
    rom[50866] = 25'b0000000010001001001100001;
    rom[50867] = 25'b0000000010001001000110010;
    rom[50868] = 25'b0000000010001001000000011;
    rom[50869] = 25'b0000000010001000111010100;
    rom[50870] = 25'b0000000010001000110100100;
    rom[50871] = 25'b0000000010001000101110101;
    rom[50872] = 25'b0000000010001000101000110;
    rom[50873] = 25'b0000000010001000100010111;
    rom[50874] = 25'b0000000010001000011100111;
    rom[50875] = 25'b0000000010001000010111000;
    rom[50876] = 25'b0000000010001000010001001;
    rom[50877] = 25'b0000000010001000001011001;
    rom[50878] = 25'b0000000010001000000101001;
    rom[50879] = 25'b0000000010000111111111001;
    rom[50880] = 25'b0000000010000111111001001;
    rom[50881] = 25'b0000000010000111110011001;
    rom[50882] = 25'b0000000010000111101101001;
    rom[50883] = 25'b0000000010000111100111001;
    rom[50884] = 25'b0000000010000111100001001;
    rom[50885] = 25'b0000000010000111011011001;
    rom[50886] = 25'b0000000010000111010101000;
    rom[50887] = 25'b0000000010000111001111000;
    rom[50888] = 25'b0000000010000111001001000;
    rom[50889] = 25'b0000000010000111000010111;
    rom[50890] = 25'b0000000010000110111100111;
    rom[50891] = 25'b0000000010000110110110110;
    rom[50892] = 25'b0000000010000110110000110;
    rom[50893] = 25'b0000000010000110101010100;
    rom[50894] = 25'b0000000010000110100100100;
    rom[50895] = 25'b0000000010000110011110011;
    rom[50896] = 25'b0000000010000110011000010;
    rom[50897] = 25'b0000000010000110010010001;
    rom[50898] = 25'b0000000010000110001100000;
    rom[50899] = 25'b0000000010000110000101111;
    rom[50900] = 25'b0000000010000101111111101;
    rom[50901] = 25'b0000000010000101111001100;
    rom[50902] = 25'b0000000010000101110011011;
    rom[50903] = 25'b0000000010000101101101001;
    rom[50904] = 25'b0000000010000101100110111;
    rom[50905] = 25'b0000000010000101100000110;
    rom[50906] = 25'b0000000010000101011010100;
    rom[50907] = 25'b0000000010000101010100011;
    rom[50908] = 25'b0000000010000101001110001;
    rom[50909] = 25'b0000000010000101000111111;
    rom[50910] = 25'b0000000010000101000001101;
    rom[50911] = 25'b0000000010000100111011011;
    rom[50912] = 25'b0000000010000100110101001;
    rom[50913] = 25'b0000000010000100101110111;
    rom[50914] = 25'b0000000010000100101000101;
    rom[50915] = 25'b0000000010000100100010010;
    rom[50916] = 25'b0000000010000100011100000;
    rom[50917] = 25'b0000000010000100010101101;
    rom[50918] = 25'b0000000010000100001111011;
    rom[50919] = 25'b0000000010000100001001001;
    rom[50920] = 25'b0000000010000100000010110;
    rom[50921] = 25'b0000000010000011111100100;
    rom[50922] = 25'b0000000010000011110110001;
    rom[50923] = 25'b0000000010000011101111110;
    rom[50924] = 25'b0000000010000011101001011;
    rom[50925] = 25'b0000000010000011100011000;
    rom[50926] = 25'b0000000010000011011100101;
    rom[50927] = 25'b0000000010000011010110010;
    rom[50928] = 25'b0000000010000011001111111;
    rom[50929] = 25'b0000000010000011001001100;
    rom[50930] = 25'b0000000010000011000011001;
    rom[50931] = 25'b0000000010000010111100101;
    rom[50932] = 25'b0000000010000010110110010;
    rom[50933] = 25'b0000000010000010101111110;
    rom[50934] = 25'b0000000010000010101001011;
    rom[50935] = 25'b0000000010000010100010111;
    rom[50936] = 25'b0000000010000010011100100;
    rom[50937] = 25'b0000000010000010010110000;
    rom[50938] = 25'b0000000010000010001111101;
    rom[50939] = 25'b0000000010000010001001000;
    rom[50940] = 25'b0000000010000010000010101;
    rom[50941] = 25'b0000000010000001111100000;
    rom[50942] = 25'b0000000010000001110101101;
    rom[50943] = 25'b0000000010000001101111001;
    rom[50944] = 25'b0000000010000001101000100;
    rom[50945] = 25'b0000000010000001100010000;
    rom[50946] = 25'b0000000010000001011011100;
    rom[50947] = 25'b0000000010000001010100111;
    rom[50948] = 25'b0000000010000001001110011;
    rom[50949] = 25'b0000000010000001000111111;
    rom[50950] = 25'b0000000010000001000001010;
    rom[50951] = 25'b0000000010000000111010101;
    rom[50952] = 25'b0000000010000000110100001;
    rom[50953] = 25'b0000000010000000101101100;
    rom[50954] = 25'b0000000010000000100111000;
    rom[50955] = 25'b0000000010000000100000011;
    rom[50956] = 25'b0000000010000000011001110;
    rom[50957] = 25'b0000000010000000010011001;
    rom[50958] = 25'b0000000010000000001100100;
    rom[50959] = 25'b0000000010000000000101111;
    rom[50960] = 25'b0000000001111111111111010;
    rom[50961] = 25'b0000000001111111111000101;
    rom[50962] = 25'b0000000001111111110001111;
    rom[50963] = 25'b0000000001111111101011010;
    rom[50964] = 25'b0000000001111111100100101;
    rom[50965] = 25'b0000000001111111011101111;
    rom[50966] = 25'b0000000001111111010111010;
    rom[50967] = 25'b0000000001111111010000100;
    rom[50968] = 25'b0000000001111111001001110;
    rom[50969] = 25'b0000000001111111000011000;
    rom[50970] = 25'b0000000001111110111100011;
    rom[50971] = 25'b0000000001111110110101101;
    rom[50972] = 25'b0000000001111110101110111;
    rom[50973] = 25'b0000000001111110101000001;
    rom[50974] = 25'b0000000001111110100001011;
    rom[50975] = 25'b0000000001111110011010101;
    rom[50976] = 25'b0000000001111110010011111;
    rom[50977] = 25'b0000000001111110001101001;
    rom[50978] = 25'b0000000001111110000110011;
    rom[50979] = 25'b0000000001111101111111100;
    rom[50980] = 25'b0000000001111101111000110;
    rom[50981] = 25'b0000000001111101110010000;
    rom[50982] = 25'b0000000001111101101011001;
    rom[50983] = 25'b0000000001111101100100011;
    rom[50984] = 25'b0000000001111101011101100;
    rom[50985] = 25'b0000000001111101010110110;
    rom[50986] = 25'b0000000001111101001111110;
    rom[50987] = 25'b0000000001111101001001000;
    rom[50988] = 25'b0000000001111101000010001;
    rom[50989] = 25'b0000000001111100111011010;
    rom[50990] = 25'b0000000001111100110100100;
    rom[50991] = 25'b0000000001111100101101100;
    rom[50992] = 25'b0000000001111100100110101;
    rom[50993] = 25'b0000000001111100011111110;
    rom[50994] = 25'b0000000001111100011000111;
    rom[50995] = 25'b0000000001111100010010000;
    rom[50996] = 25'b0000000001111100001011001;
    rom[50997] = 25'b0000000001111100000100001;
    rom[50998] = 25'b0000000001111011111101010;
    rom[50999] = 25'b0000000001111011110110010;
    rom[51000] = 25'b0000000001111011101111011;
    rom[51001] = 25'b0000000001111011101000011;
    rom[51002] = 25'b0000000001111011100001011;
    rom[51003] = 25'b0000000001111011011010100;
    rom[51004] = 25'b0000000001111011010011100;
    rom[51005] = 25'b0000000001111011001100100;
    rom[51006] = 25'b0000000001111011000101101;
    rom[51007] = 25'b0000000001111010111110101;
    rom[51008] = 25'b0000000001111010110111101;
    rom[51009] = 25'b0000000001111010110000101;
    rom[51010] = 25'b0000000001111010101001101;
    rom[51011] = 25'b0000000001111010100010101;
    rom[51012] = 25'b0000000001111010011011100;
    rom[51013] = 25'b0000000001111010010100100;
    rom[51014] = 25'b0000000001111010001101100;
    rom[51015] = 25'b0000000001111010000110011;
    rom[51016] = 25'b0000000001111001111111011;
    rom[51017] = 25'b0000000001111001111000010;
    rom[51018] = 25'b0000000001111001110001010;
    rom[51019] = 25'b0000000001111001101010001;
    rom[51020] = 25'b0000000001111001100011001;
    rom[51021] = 25'b0000000001111001011100000;
    rom[51022] = 25'b0000000001111001010100111;
    rom[51023] = 25'b0000000001111001001101110;
    rom[51024] = 25'b0000000001111001000110101;
    rom[51025] = 25'b0000000001111000111111101;
    rom[51026] = 25'b0000000001111000111000100;
    rom[51027] = 25'b0000000001111000110001010;
    rom[51028] = 25'b0000000001111000101010010;
    rom[51029] = 25'b0000000001111000100011001;
    rom[51030] = 25'b0000000001111000011011111;
    rom[51031] = 25'b0000000001111000010100110;
    rom[51032] = 25'b0000000001111000001101101;
    rom[51033] = 25'b0000000001111000000110011;
    rom[51034] = 25'b0000000001110111111111010;
    rom[51035] = 25'b0000000001110111111000000;
    rom[51036] = 25'b0000000001110111110000111;
    rom[51037] = 25'b0000000001110111101001101;
    rom[51038] = 25'b0000000001110111100010100;
    rom[51039] = 25'b0000000001110111011011010;
    rom[51040] = 25'b0000000001110111010100001;
    rom[51041] = 25'b0000000001110111001100111;
    rom[51042] = 25'b0000000001110111000101101;
    rom[51043] = 25'b0000000001110110111110011;
    rom[51044] = 25'b0000000001110110110111001;
    rom[51045] = 25'b0000000001110110101111111;
    rom[51046] = 25'b0000000001110110101000101;
    rom[51047] = 25'b0000000001110110100001011;
    rom[51048] = 25'b0000000001110110011010001;
    rom[51049] = 25'b0000000001110110010010111;
    rom[51050] = 25'b0000000001110110001011100;
    rom[51051] = 25'b0000000001110110000100010;
    rom[51052] = 25'b0000000001110101111101000;
    rom[51053] = 25'b0000000001110101110101101;
    rom[51054] = 25'b0000000001110101101110011;
    rom[51055] = 25'b0000000001110101100111001;
    rom[51056] = 25'b0000000001110101011111110;
    rom[51057] = 25'b0000000001110101011000100;
    rom[51058] = 25'b0000000001110101010001001;
    rom[51059] = 25'b0000000001110101001001110;
    rom[51060] = 25'b0000000001110101000010011;
    rom[51061] = 25'b0000000001110100111011001;
    rom[51062] = 25'b0000000001110100110011110;
    rom[51063] = 25'b0000000001110100101100011;
    rom[51064] = 25'b0000000001110100100101000;
    rom[51065] = 25'b0000000001110100011101101;
    rom[51066] = 25'b0000000001110100010110010;
    rom[51067] = 25'b0000000001110100001110111;
    rom[51068] = 25'b0000000001110100000111100;
    rom[51069] = 25'b0000000001110100000000001;
    rom[51070] = 25'b0000000001110011111000101;
    rom[51071] = 25'b0000000001110011110001010;
    rom[51072] = 25'b0000000001110011101001111;
    rom[51073] = 25'b0000000001110011100010011;
    rom[51074] = 25'b0000000001110011011011000;
    rom[51075] = 25'b0000000001110011010011101;
    rom[51076] = 25'b0000000001110011001100001;
    rom[51077] = 25'b0000000001110011000100110;
    rom[51078] = 25'b0000000001110010111101010;
    rom[51079] = 25'b0000000001110010110101110;
    rom[51080] = 25'b0000000001110010101110010;
    rom[51081] = 25'b0000000001110010100110111;
    rom[51082] = 25'b0000000001110010011111011;
    rom[51083] = 25'b0000000001110010010111111;
    rom[51084] = 25'b0000000001110010010000011;
    rom[51085] = 25'b0000000001110010001000111;
    rom[51086] = 25'b0000000001110010000001011;
    rom[51087] = 25'b0000000001110001111001111;
    rom[51088] = 25'b0000000001110001110010011;
    rom[51089] = 25'b0000000001110001101010111;
    rom[51090] = 25'b0000000001110001100011011;
    rom[51091] = 25'b0000000001110001011011110;
    rom[51092] = 25'b0000000001110001010100010;
    rom[51093] = 25'b0000000001110001001100110;
    rom[51094] = 25'b0000000001110001000101001;
    rom[51095] = 25'b0000000001110000111101101;
    rom[51096] = 25'b0000000001110000110110000;
    rom[51097] = 25'b0000000001110000101110100;
    rom[51098] = 25'b0000000001110000100110111;
    rom[51099] = 25'b0000000001110000011111011;
    rom[51100] = 25'b0000000001110000010111110;
    rom[51101] = 25'b0000000001110000010000010;
    rom[51102] = 25'b0000000001110000001000100;
    rom[51103] = 25'b0000000001110000000001000;
    rom[51104] = 25'b0000000001101111111001011;
    rom[51105] = 25'b0000000001101111110001110;
    rom[51106] = 25'b0000000001101111101010001;
    rom[51107] = 25'b0000000001101111100010100;
    rom[51108] = 25'b0000000001101111011010111;
    rom[51109] = 25'b0000000001101111010011010;
    rom[51110] = 25'b0000000001101111001011100;
    rom[51111] = 25'b0000000001101111000100000;
    rom[51112] = 25'b0000000001101110111100011;
    rom[51113] = 25'b0000000001101110110100101;
    rom[51114] = 25'b0000000001101110101101000;
    rom[51115] = 25'b0000000001101110100101011;
    rom[51116] = 25'b0000000001101110011101101;
    rom[51117] = 25'b0000000001101110010110000;
    rom[51118] = 25'b0000000001101110001110010;
    rom[51119] = 25'b0000000001101110000110101;
    rom[51120] = 25'b0000000001101101111110111;
    rom[51121] = 25'b0000000001101101110111010;
    rom[51122] = 25'b0000000001101101101111100;
    rom[51123] = 25'b0000000001101101100111111;
    rom[51124] = 25'b0000000001101101100000001;
    rom[51125] = 25'b0000000001101101011000011;
    rom[51126] = 25'b0000000001101101010000101;
    rom[51127] = 25'b0000000001101101001000111;
    rom[51128] = 25'b0000000001101101000001001;
    rom[51129] = 25'b0000000001101100111001011;
    rom[51130] = 25'b0000000001101100110001101;
    rom[51131] = 25'b0000000001101100101001111;
    rom[51132] = 25'b0000000001101100100010001;
    rom[51133] = 25'b0000000001101100011010011;
    rom[51134] = 25'b0000000001101100010010101;
    rom[51135] = 25'b0000000001101100001010110;
    rom[51136] = 25'b0000000001101100000011000;
    rom[51137] = 25'b0000000001101011111011010;
    rom[51138] = 25'b0000000001101011110011100;
    rom[51139] = 25'b0000000001101011101011110;
    rom[51140] = 25'b0000000001101011100011111;
    rom[51141] = 25'b0000000001101011011100001;
    rom[51142] = 25'b0000000001101011010100010;
    rom[51143] = 25'b0000000001101011001100011;
    rom[51144] = 25'b0000000001101011000100101;
    rom[51145] = 25'b0000000001101010111100111;
    rom[51146] = 25'b0000000001101010110101000;
    rom[51147] = 25'b0000000001101010101101001;
    rom[51148] = 25'b0000000001101010100101010;
    rom[51149] = 25'b0000000001101010011101100;
    rom[51150] = 25'b0000000001101010010101101;
    rom[51151] = 25'b0000000001101010001101110;
    rom[51152] = 25'b0000000001101010000101111;
    rom[51153] = 25'b0000000001101001111110000;
    rom[51154] = 25'b0000000001101001110110001;
    rom[51155] = 25'b0000000001101001101110010;
    rom[51156] = 25'b0000000001101001100110011;
    rom[51157] = 25'b0000000001101001011110100;
    rom[51158] = 25'b0000000001101001010110101;
    rom[51159] = 25'b0000000001101001001110110;
    rom[51160] = 25'b0000000001101001000110110;
    rom[51161] = 25'b0000000001101000111110111;
    rom[51162] = 25'b0000000001101000110111000;
    rom[51163] = 25'b0000000001101000101111001;
    rom[51164] = 25'b0000000001101000100111001;
    rom[51165] = 25'b0000000001101000011111010;
    rom[51166] = 25'b0000000001101000010111010;
    rom[51167] = 25'b0000000001101000001111011;
    rom[51168] = 25'b0000000001101000000111011;
    rom[51169] = 25'b0000000001100111111111100;
    rom[51170] = 25'b0000000001100111110111100;
    rom[51171] = 25'b0000000001100111101111101;
    rom[51172] = 25'b0000000001100111100111101;
    rom[51173] = 25'b0000000001100111011111101;
    rom[51174] = 25'b0000000001100111010111101;
    rom[51175] = 25'b0000000001100111001111110;
    rom[51176] = 25'b0000000001100111000111110;
    rom[51177] = 25'b0000000001100110111111110;
    rom[51178] = 25'b0000000001100110110111110;
    rom[51179] = 25'b0000000001100110101111110;
    rom[51180] = 25'b0000000001100110100111110;
    rom[51181] = 25'b0000000001100110011111110;
    rom[51182] = 25'b0000000001100110010111110;
    rom[51183] = 25'b0000000001100110001111110;
    rom[51184] = 25'b0000000001100110000111110;
    rom[51185] = 25'b0000000001100101111111110;
    rom[51186] = 25'b0000000001100101110111101;
    rom[51187] = 25'b0000000001100101101111101;
    rom[51188] = 25'b0000000001100101100111101;
    rom[51189] = 25'b0000000001100101011111101;
    rom[51190] = 25'b0000000001100101010111100;
    rom[51191] = 25'b0000000001100101001111100;
    rom[51192] = 25'b0000000001100101000111100;
    rom[51193] = 25'b0000000001100100111111100;
    rom[51194] = 25'b0000000001100100110111011;
    rom[51195] = 25'b0000000001100100101111010;
    rom[51196] = 25'b0000000001100100100111001;
    rom[51197] = 25'b0000000001100100011111001;
    rom[51198] = 25'b0000000001100100010111001;
    rom[51199] = 25'b0000000001100100001111000;
    rom[51200] = 25'b0000000001100100000110111;
    rom[51201] = 25'b0000000001100011111110111;
    rom[51202] = 25'b0000000001100011110110110;
    rom[51203] = 25'b0000000001100011101110101;
    rom[51204] = 25'b0000000001100011100110100;
    rom[51205] = 25'b0000000001100011011110011;
    rom[51206] = 25'b0000000001100011010110010;
    rom[51207] = 25'b0000000001100011001110001;
    rom[51208] = 25'b0000000001100011000110000;
    rom[51209] = 25'b0000000001100010111101111;
    rom[51210] = 25'b0000000001100010110101110;
    rom[51211] = 25'b0000000001100010101101101;
    rom[51212] = 25'b0000000001100010100101100;
    rom[51213] = 25'b0000000001100010011101011;
    rom[51214] = 25'b0000000001100010010101010;
    rom[51215] = 25'b0000000001100010001101001;
    rom[51216] = 25'b0000000001100010000101000;
    rom[51217] = 25'b0000000001100001111100111;
    rom[51218] = 25'b0000000001100001110100101;
    rom[51219] = 25'b0000000001100001101100100;
    rom[51220] = 25'b0000000001100001100100010;
    rom[51221] = 25'b0000000001100001011100001;
    rom[51222] = 25'b0000000001100001010011111;
    rom[51223] = 25'b0000000001100001001011110;
    rom[51224] = 25'b0000000001100001000011101;
    rom[51225] = 25'b0000000001100000111011011;
    rom[51226] = 25'b0000000001100000110011001;
    rom[51227] = 25'b0000000001100000101011000;
    rom[51228] = 25'b0000000001100000100010110;
    rom[51229] = 25'b0000000001100000011010101;
    rom[51230] = 25'b0000000001100000010010011;
    rom[51231] = 25'b0000000001100000001010001;
    rom[51232] = 25'b0000000001100000000001111;
    rom[51233] = 25'b0000000001011111111001110;
    rom[51234] = 25'b0000000001011111110001100;
    rom[51235] = 25'b0000000001011111101001010;
    rom[51236] = 25'b0000000001011111100001000;
    rom[51237] = 25'b0000000001011111011000111;
    rom[51238] = 25'b0000000001011111010000100;
    rom[51239] = 25'b0000000001011111001000010;
    rom[51240] = 25'b0000000001011111000000001;
    rom[51241] = 25'b0000000001011110110111110;
    rom[51242] = 25'b0000000001011110101111100;
    rom[51243] = 25'b0000000001011110100111011;
    rom[51244] = 25'b0000000001011110011111000;
    rom[51245] = 25'b0000000001011110010110110;
    rom[51246] = 25'b0000000001011110001110100;
    rom[51247] = 25'b0000000001011110000110001;
    rom[51248] = 25'b0000000001011101111110000;
    rom[51249] = 25'b0000000001011101110101101;
    rom[51250] = 25'b0000000001011101101101011;
    rom[51251] = 25'b0000000001011101100101001;
    rom[51252] = 25'b0000000001011101011100111;
    rom[51253] = 25'b0000000001011101010100100;
    rom[51254] = 25'b0000000001011101001100010;
    rom[51255] = 25'b0000000001011101000011111;
    rom[51256] = 25'b0000000001011100111011101;
    rom[51257] = 25'b0000000001011100110011010;
    rom[51258] = 25'b0000000001011100101011000;
    rom[51259] = 25'b0000000001011100100010101;
    rom[51260] = 25'b0000000001011100011010011;
    rom[51261] = 25'b0000000001011100010010000;
    rom[51262] = 25'b0000000001011100001001110;
    rom[51263] = 25'b0000000001011100000001011;
    rom[51264] = 25'b0000000001011011111001000;
    rom[51265] = 25'b0000000001011011110000101;
    rom[51266] = 25'b0000000001011011101000011;
    rom[51267] = 25'b0000000001011011100000000;
    rom[51268] = 25'b0000000001011011010111101;
    rom[51269] = 25'b0000000001011011001111011;
    rom[51270] = 25'b0000000001011011000110111;
    rom[51271] = 25'b0000000001011010111110101;
    rom[51272] = 25'b0000000001011010110110010;
    rom[51273] = 25'b0000000001011010101101111;
    rom[51274] = 25'b0000000001011010100101100;
    rom[51275] = 25'b0000000001011010011101001;
    rom[51276] = 25'b0000000001011010010100110;
    rom[51277] = 25'b0000000001011010001100011;
    rom[51278] = 25'b0000000001011010000100000;
    rom[51279] = 25'b0000000001011001111011101;
    rom[51280] = 25'b0000000001011001110011010;
    rom[51281] = 25'b0000000001011001101010111;
    rom[51282] = 25'b0000000001011001100010100;
    rom[51283] = 25'b0000000001011001011010000;
    rom[51284] = 25'b0000000001011001010001101;
    rom[51285] = 25'b0000000001011001001001010;
    rom[51286] = 25'b0000000001011001000000111;
    rom[51287] = 25'b0000000001011000111000011;
    rom[51288] = 25'b0000000001011000110000000;
    rom[51289] = 25'b0000000001011000100111101;
    rom[51290] = 25'b0000000001011000011111010;
    rom[51291] = 25'b0000000001011000010110110;
    rom[51292] = 25'b0000000001011000001110010;
    rom[51293] = 25'b0000000001011000000101111;
    rom[51294] = 25'b0000000001010111111101100;
    rom[51295] = 25'b0000000001010111110101000;
    rom[51296] = 25'b0000000001010111101100101;
    rom[51297] = 25'b0000000001010111100100001;
    rom[51298] = 25'b0000000001010111011011110;
    rom[51299] = 25'b0000000001010111010011010;
    rom[51300] = 25'b0000000001010111001010110;
    rom[51301] = 25'b0000000001010111000010011;
    rom[51302] = 25'b0000000001010110111001111;
    rom[51303] = 25'b0000000001010110110001100;
    rom[51304] = 25'b0000000001010110101001000;
    rom[51305] = 25'b0000000001010110100000101;
    rom[51306] = 25'b0000000001010110011000001;
    rom[51307] = 25'b0000000001010110001111101;
    rom[51308] = 25'b0000000001010110000111001;
    rom[51309] = 25'b0000000001010101111110101;
    rom[51310] = 25'b0000000001010101110110001;
    rom[51311] = 25'b0000000001010101101101101;
    rom[51312] = 25'b0000000001010101100101001;
    rom[51313] = 25'b0000000001010101011100110;
    rom[51314] = 25'b0000000001010101010100010;
    rom[51315] = 25'b0000000001010101001011110;
    rom[51316] = 25'b0000000001010101000011010;
    rom[51317] = 25'b0000000001010100111010110;
    rom[51318] = 25'b0000000001010100110010010;
    rom[51319] = 25'b0000000001010100101001110;
    rom[51320] = 25'b0000000001010100100001010;
    rom[51321] = 25'b0000000001010100011000110;
    rom[51322] = 25'b0000000001010100010000010;
    rom[51323] = 25'b0000000001010100000111110;
    rom[51324] = 25'b0000000001010011111111010;
    rom[51325] = 25'b0000000001010011110110110;
    rom[51326] = 25'b0000000001010011101110010;
    rom[51327] = 25'b0000000001010011100101101;
    rom[51328] = 25'b0000000001010011011101001;
    rom[51329] = 25'b0000000001010011010100101;
    rom[51330] = 25'b0000000001010011001100000;
    rom[51331] = 25'b0000000001010011000011100;
    rom[51332] = 25'b0000000001010010111011000;
    rom[51333] = 25'b0000000001010010110010011;
    rom[51334] = 25'b0000000001010010101010000;
    rom[51335] = 25'b0000000001010010100001011;
    rom[51336] = 25'b0000000001010010011000111;
    rom[51337] = 25'b0000000001010010010000010;
    rom[51338] = 25'b0000000001010010000111110;
    rom[51339] = 25'b0000000001010001111111001;
    rom[51340] = 25'b0000000001010001110110101;
    rom[51341] = 25'b0000000001010001101110001;
    rom[51342] = 25'b0000000001010001100101100;
    rom[51343] = 25'b0000000001010001011101000;
    rom[51344] = 25'b0000000001010001010100011;
    rom[51345] = 25'b0000000001010001001011110;
    rom[51346] = 25'b0000000001010001000011010;
    rom[51347] = 25'b0000000001010000111010110;
    rom[51348] = 25'b0000000001010000110010001;
    rom[51349] = 25'b0000000001010000101001100;
    rom[51350] = 25'b0000000001010000100001000;
    rom[51351] = 25'b0000000001010000011000011;
    rom[51352] = 25'b0000000001010000001111110;
    rom[51353] = 25'b0000000001010000000111001;
    rom[51354] = 25'b0000000001001111111110101;
    rom[51355] = 25'b0000000001001111110110000;
    rom[51356] = 25'b0000000001001111101101011;
    rom[51357] = 25'b0000000001001111100100110;
    rom[51358] = 25'b0000000001001111011100010;
    rom[51359] = 25'b0000000001001111010011101;
    rom[51360] = 25'b0000000001001111001011000;
    rom[51361] = 25'b0000000001001111000010011;
    rom[51362] = 25'b0000000001001110111001111;
    rom[51363] = 25'b0000000001001110110001010;
    rom[51364] = 25'b0000000001001110101000101;
    rom[51365] = 25'b0000000001001110100000000;
    rom[51366] = 25'b0000000001001110010111011;
    rom[51367] = 25'b0000000001001110001110110;
    rom[51368] = 25'b0000000001001110000110010;
    rom[51369] = 25'b0000000001001101111101100;
    rom[51370] = 25'b0000000001001101110100111;
    rom[51371] = 25'b0000000001001101101100011;
    rom[51372] = 25'b0000000001001101100011101;
    rom[51373] = 25'b0000000001001101011011000;
    rom[51374] = 25'b0000000001001101010010100;
    rom[51375] = 25'b0000000001001101001001110;
    rom[51376] = 25'b0000000001001101000001001;
    rom[51377] = 25'b0000000001001100111000100;
    rom[51378] = 25'b0000000001001100101111111;
    rom[51379] = 25'b0000000001001100100111010;
    rom[51380] = 25'b0000000001001100011110101;
    rom[51381] = 25'b0000000001001100010110000;
    rom[51382] = 25'b0000000001001100001101011;
    rom[51383] = 25'b0000000001001100000100101;
    rom[51384] = 25'b0000000001001011111100001;
    rom[51385] = 25'b0000000001001011110011011;
    rom[51386] = 25'b0000000001001011101010110;
    rom[51387] = 25'b0000000001001011100010001;
    rom[51388] = 25'b0000000001001011011001011;
    rom[51389] = 25'b0000000001001011010000110;
    rom[51390] = 25'b0000000001001011001000001;
    rom[51391] = 25'b0000000001001010111111100;
    rom[51392] = 25'b0000000001001010110110110;
    rom[51393] = 25'b0000000001001010101110001;
    rom[51394] = 25'b0000000001001010100101100;
    rom[51395] = 25'b0000000001001010011100111;
    rom[51396] = 25'b0000000001001010010100001;
    rom[51397] = 25'b0000000001001010001011100;
    rom[51398] = 25'b0000000001001010000010110;
    rom[51399] = 25'b0000000001001001111010001;
    rom[51400] = 25'b0000000001001001110001011;
    rom[51401] = 25'b0000000001001001101000110;
    rom[51402] = 25'b0000000001001001100000001;
    rom[51403] = 25'b0000000001001001010111011;
    rom[51404] = 25'b0000000001001001001110110;
    rom[51405] = 25'b0000000001001001000110001;
    rom[51406] = 25'b0000000001001000111101011;
    rom[51407] = 25'b0000000001001000110100110;
    rom[51408] = 25'b0000000001001000101100000;
    rom[51409] = 25'b0000000001001000100011011;
    rom[51410] = 25'b0000000001001000011010101;
    rom[51411] = 25'b0000000001001000010010000;
    rom[51412] = 25'b0000000001001000001001010;
    rom[51413] = 25'b0000000001001000000000101;
    rom[51414] = 25'b0000000001000111110111110;
    rom[51415] = 25'b0000000001000111101111001;
    rom[51416] = 25'b0000000001000111100110100;
    rom[51417] = 25'b0000000001000111011101110;
    rom[51418] = 25'b0000000001000111010101001;
    rom[51419] = 25'b0000000001000111001100011;
    rom[51420] = 25'b0000000001000111000011101;
    rom[51421] = 25'b0000000001000110111010111;
    rom[51422] = 25'b0000000001000110110010010;
    rom[51423] = 25'b0000000001000110101001100;
    rom[51424] = 25'b0000000001000110100000111;
    rom[51425] = 25'b0000000001000110011000001;
    rom[51426] = 25'b0000000001000110001111011;
    rom[51427] = 25'b0000000001000110000110110;
    rom[51428] = 25'b0000000001000101111110000;
    rom[51429] = 25'b0000000001000101110101010;
    rom[51430] = 25'b0000000001000101101100101;
    rom[51431] = 25'b0000000001000101100011110;
    rom[51432] = 25'b0000000001000101011011001;
    rom[51433] = 25'b0000000001000101010010011;
    rom[51434] = 25'b0000000001000101001001101;
    rom[51435] = 25'b0000000001000101000001000;
    rom[51436] = 25'b0000000001000100111000010;
    rom[51437] = 25'b0000000001000100101111100;
    rom[51438] = 25'b0000000001000100100110110;
    rom[51439] = 25'b0000000001000100011110000;
    rom[51440] = 25'b0000000001000100010101011;
    rom[51441] = 25'b0000000001000100001100101;
    rom[51442] = 25'b0000000001000100000011111;
    rom[51443] = 25'b0000000001000011111011001;
    rom[51444] = 25'b0000000001000011110010011;
    rom[51445] = 25'b0000000001000011101001101;
    rom[51446] = 25'b0000000001000011100001000;
    rom[51447] = 25'b0000000001000011011000001;
    rom[51448] = 25'b0000000001000011001111100;
    rom[51449] = 25'b0000000001000011000110110;
    rom[51450] = 25'b0000000001000010111110000;
    rom[51451] = 25'b0000000001000010110101010;
    rom[51452] = 25'b0000000001000010101100101;
    rom[51453] = 25'b0000000001000010100011110;
    rom[51454] = 25'b0000000001000010011011000;
    rom[51455] = 25'b0000000001000010010010011;
    rom[51456] = 25'b0000000001000010001001100;
    rom[51457] = 25'b0000000001000010000000111;
    rom[51458] = 25'b0000000001000001111000001;
    rom[51459] = 25'b0000000001000001101111010;
    rom[51460] = 25'b0000000001000001100110101;
    rom[51461] = 25'b0000000001000001011101111;
    rom[51462] = 25'b0000000001000001010101000;
    rom[51463] = 25'b0000000001000001001100011;
    rom[51464] = 25'b0000000001000001000011101;
    rom[51465] = 25'b0000000001000000111010111;
    rom[51466] = 25'b0000000001000000110010001;
    rom[51467] = 25'b0000000001000000101001011;
    rom[51468] = 25'b0000000001000000100000101;
    rom[51469] = 25'b0000000001000000010111110;
    rom[51470] = 25'b0000000001000000001111001;
    rom[51471] = 25'b0000000001000000000110011;
    rom[51472] = 25'b0000000000111111111101100;
    rom[51473] = 25'b0000000000111111110100111;
    rom[51474] = 25'b0000000000111111101100001;
    rom[51475] = 25'b0000000000111111100011011;
    rom[51476] = 25'b0000000000111111011010100;
    rom[51477] = 25'b0000000000111111010001110;
    rom[51478] = 25'b0000000000111111001001001;
    rom[51479] = 25'b0000000000111111000000010;
    rom[51480] = 25'b0000000000111110110111100;
    rom[51481] = 25'b0000000000111110101110110;
    rom[51482] = 25'b0000000000111110100110000;
    rom[51483] = 25'b0000000000111110011101010;
    rom[51484] = 25'b0000000000111110010100100;
    rom[51485] = 25'b0000000000111110001011110;
    rom[51486] = 25'b0000000000111110000011000;
    rom[51487] = 25'b0000000000111101111010001;
    rom[51488] = 25'b0000000000111101110001100;
    rom[51489] = 25'b0000000000111101101000110;
    rom[51490] = 25'b0000000000111101011111111;
    rom[51491] = 25'b0000000000111101010111001;
    rom[51492] = 25'b0000000000111101001110011;
    rom[51493] = 25'b0000000000111101000101101;
    rom[51494] = 25'b0000000000111100111100111;
    rom[51495] = 25'b0000000000111100110100001;
    rom[51496] = 25'b0000000000111100101011011;
    rom[51497] = 25'b0000000000111100100010101;
    rom[51498] = 25'b0000000000111100011001110;
    rom[51499] = 25'b0000000000111100010001000;
    rom[51500] = 25'b0000000000111100001000010;
    rom[51501] = 25'b0000000000111011111111100;
    rom[51502] = 25'b0000000000111011110110110;
    rom[51503] = 25'b0000000000111011101110000;
    rom[51504] = 25'b0000000000111011100101010;
    rom[51505] = 25'b0000000000111011011100011;
    rom[51506] = 25'b0000000000111011010011101;
    rom[51507] = 25'b0000000000111011001010111;
    rom[51508] = 25'b0000000000111011000010001;
    rom[51509] = 25'b0000000000111010111001011;
    rom[51510] = 25'b0000000000111010110000100;
    rom[51511] = 25'b0000000000111010100111110;
    rom[51512] = 25'b0000000000111010011111001;
    rom[51513] = 25'b0000000000111010010110010;
    rom[51514] = 25'b0000000000111010001101100;
    rom[51515] = 25'b0000000000111010000100110;
    rom[51516] = 25'b0000000000111001111100000;
    rom[51517] = 25'b0000000000111001110011001;
    rom[51518] = 25'b0000000000111001101010011;
    rom[51519] = 25'b0000000000111001100001101;
    rom[51520] = 25'b0000000000111001011000111;
    rom[51521] = 25'b0000000000111001010000001;
    rom[51522] = 25'b0000000000111001000111010;
    rom[51523] = 25'b0000000000111000111110101;
    rom[51524] = 25'b0000000000111000110101111;
    rom[51525] = 25'b0000000000111000101101000;
    rom[51526] = 25'b0000000000111000100100010;
    rom[51527] = 25'b0000000000111000011011100;
    rom[51528] = 25'b0000000000111000010010110;
    rom[51529] = 25'b0000000000111000001001111;
    rom[51530] = 25'b0000000000111000000001001;
    rom[51531] = 25'b0000000000110111111000011;
    rom[51532] = 25'b0000000000110111101111101;
    rom[51533] = 25'b0000000000110111100110111;
    rom[51534] = 25'b0000000000110111011110001;
    rom[51535] = 25'b0000000000110111010101011;
    rom[51536] = 25'b0000000000110111001100101;
    rom[51537] = 25'b0000000000110111000011110;
    rom[51538] = 25'b0000000000110110111011000;
    rom[51539] = 25'b0000000000110110110010010;
    rom[51540] = 25'b0000000000110110101001100;
    rom[51541] = 25'b0000000000110110100000110;
    rom[51542] = 25'b0000000000110110010111111;
    rom[51543] = 25'b0000000000110110001111010;
    rom[51544] = 25'b0000000000110110000110100;
    rom[51545] = 25'b0000000000110101111101101;
    rom[51546] = 25'b0000000000110101110100111;
    rom[51547] = 25'b0000000000110101101100001;
    rom[51548] = 25'b0000000000110101100011011;
    rom[51549] = 25'b0000000000110101011010100;
    rom[51550] = 25'b0000000000110101010001110;
    rom[51551] = 25'b0000000000110101001001001;
    rom[51552] = 25'b0000000000110101000000011;
    rom[51553] = 25'b0000000000110100110111100;
    rom[51554] = 25'b0000000000110100101110110;
    rom[51555] = 25'b0000000000110100100110000;
    rom[51556] = 25'b0000000000110100011101010;
    rom[51557] = 25'b0000000000110100010100100;
    rom[51558] = 25'b0000000000110100001011110;
    rom[51559] = 25'b0000000000110100000011000;
    rom[51560] = 25'b0000000000110011111010001;
    rom[51561] = 25'b0000000000110011110001011;
    rom[51562] = 25'b0000000000110011101000101;
    rom[51563] = 25'b0000000000110011100000000;
    rom[51564] = 25'b0000000000110011010111001;
    rom[51565] = 25'b0000000000110011001110011;
    rom[51566] = 25'b0000000000110011000101101;
    rom[51567] = 25'b0000000000110010111100111;
    rom[51568] = 25'b0000000000110010110100001;
    rom[51569] = 25'b0000000000110010101011011;
    rom[51570] = 25'b0000000000110010100010101;
    rom[51571] = 25'b0000000000110010011001110;
    rom[51572] = 25'b0000000000110010010001001;
    rom[51573] = 25'b0000000000110010001000011;
    rom[51574] = 25'b0000000000110001111111101;
    rom[51575] = 25'b0000000000110001110110110;
    rom[51576] = 25'b0000000000110001101110001;
    rom[51577] = 25'b0000000000110001100101011;
    rom[51578] = 25'b0000000000110001011100100;
    rom[51579] = 25'b0000000000110001010011111;
    rom[51580] = 25'b0000000000110001001011001;
    rom[51581] = 25'b0000000000110001000010010;
    rom[51582] = 25'b0000000000110000111001101;
    rom[51583] = 25'b0000000000110000110000111;
    rom[51584] = 25'b0000000000110000101000000;
    rom[51585] = 25'b0000000000110000011111011;
    rom[51586] = 25'b0000000000110000010110101;
    rom[51587] = 25'b0000000000110000001101111;
    rom[51588] = 25'b0000000000110000000101001;
    rom[51589] = 25'b0000000000101111111100011;
    rom[51590] = 25'b0000000000101111110011101;
    rom[51591] = 25'b0000000000101111101010111;
    rom[51592] = 25'b0000000000101111100010001;
    rom[51593] = 25'b0000000000101111011001011;
    rom[51594] = 25'b0000000000101111010000101;
    rom[51595] = 25'b0000000000101111001000000;
    rom[51596] = 25'b0000000000101110111111001;
    rom[51597] = 25'b0000000000101110110110011;
    rom[51598] = 25'b0000000000101110101101110;
    rom[51599] = 25'b0000000000101110100101000;
    rom[51600] = 25'b0000000000101110011100010;
    rom[51601] = 25'b0000000000101110010011100;
    rom[51602] = 25'b0000000000101110001010110;
    rom[51603] = 25'b0000000000101110000010000;
    rom[51604] = 25'b0000000000101101111001011;
    rom[51605] = 25'b0000000000101101110000100;
    rom[51606] = 25'b0000000000101101100111111;
    rom[51607] = 25'b0000000000101101011111001;
    rom[51608] = 25'b0000000000101101010110011;
    rom[51609] = 25'b0000000000101101001101110;
    rom[51610] = 25'b0000000000101101000101000;
    rom[51611] = 25'b0000000000101100111100010;
    rom[51612] = 25'b0000000000101100110011100;
    rom[51613] = 25'b0000000000101100101010110;
    rom[51614] = 25'b0000000000101100100010001;
    rom[51615] = 25'b0000000000101100011001011;
    rom[51616] = 25'b0000000000101100010000101;
    rom[51617] = 25'b0000000000101100001000000;
    rom[51618] = 25'b0000000000101011111111001;
    rom[51619] = 25'b0000000000101011110110100;
    rom[51620] = 25'b0000000000101011101101111;
    rom[51621] = 25'b0000000000101011100101001;
    rom[51622] = 25'b0000000000101011011100011;
    rom[51623] = 25'b0000000000101011010011101;
    rom[51624] = 25'b0000000000101011001011000;
    rom[51625] = 25'b0000000000101011000010010;
    rom[51626] = 25'b0000000000101010111001100;
    rom[51627] = 25'b0000000000101010110000111;
    rom[51628] = 25'b0000000000101010101000001;
    rom[51629] = 25'b0000000000101010011111100;
    rom[51630] = 25'b0000000000101010010110110;
    rom[51631] = 25'b0000000000101010001110001;
    rom[51632] = 25'b0000000000101010000101011;
    rom[51633] = 25'b0000000000101001111100101;
    rom[51634] = 25'b0000000000101001110100000;
    rom[51635] = 25'b0000000000101001101011010;
    rom[51636] = 25'b0000000000101001100010101;
    rom[51637] = 25'b0000000000101001011001111;
    rom[51638] = 25'b0000000000101001010001010;
    rom[51639] = 25'b0000000000101001001000100;
    rom[51640] = 25'b0000000000101000111111111;
    rom[51641] = 25'b0000000000101000110111001;
    rom[51642] = 25'b0000000000101000101110100;
    rom[51643] = 25'b0000000000101000100101110;
    rom[51644] = 25'b0000000000101000011101001;
    rom[51645] = 25'b0000000000101000010100011;
    rom[51646] = 25'b0000000000101000001011110;
    rom[51647] = 25'b0000000000101000000011000;
    rom[51648] = 25'b0000000000100111111010011;
    rom[51649] = 25'b0000000000100111110001110;
    rom[51650] = 25'b0000000000100111101001001;
    rom[51651] = 25'b0000000000100111100000011;
    rom[51652] = 25'b0000000000100111010111110;
    rom[51653] = 25'b0000000000100111001111000;
    rom[51654] = 25'b0000000000100111000110011;
    rom[51655] = 25'b0000000000100110111101110;
    rom[51656] = 25'b0000000000100110110101000;
    rom[51657] = 25'b0000000000100110101100011;
    rom[51658] = 25'b0000000000100110100011110;
    rom[51659] = 25'b0000000000100110011011001;
    rom[51660] = 25'b0000000000100110010010011;
    rom[51661] = 25'b0000000000100110001001110;
    rom[51662] = 25'b0000000000100110000001001;
    rom[51663] = 25'b0000000000100101111000100;
    rom[51664] = 25'b0000000000100101101111111;
    rom[51665] = 25'b0000000000100101100111001;
    rom[51666] = 25'b0000000000100101011110100;
    rom[51667] = 25'b0000000000100101010101111;
    rom[51668] = 25'b0000000000100101001101010;
    rom[51669] = 25'b0000000000100101000100101;
    rom[51670] = 25'b0000000000100100111011111;
    rom[51671] = 25'b0000000000100100110011011;
    rom[51672] = 25'b0000000000100100101010101;
    rom[51673] = 25'b0000000000100100100010001;
    rom[51674] = 25'b0000000000100100011001100;
    rom[51675] = 25'b0000000000100100010000110;
    rom[51676] = 25'b0000000000100100001000010;
    rom[51677] = 25'b0000000000100011111111100;
    rom[51678] = 25'b0000000000100011110110111;
    rom[51679] = 25'b0000000000100011101110011;
    rom[51680] = 25'b0000000000100011100101101;
    rom[51681] = 25'b0000000000100011011101000;
    rom[51682] = 25'b0000000000100011010100100;
    rom[51683] = 25'b0000000000100011001011111;
    rom[51684] = 25'b0000000000100011000011001;
    rom[51685] = 25'b0000000000100010111010101;
    rom[51686] = 25'b0000000000100010110010000;
    rom[51687] = 25'b0000000000100010101001011;
    rom[51688] = 25'b0000000000100010100000111;
    rom[51689] = 25'b0000000000100010011000010;
    rom[51690] = 25'b0000000000100010001111100;
    rom[51691] = 25'b0000000000100010000111000;
    rom[51692] = 25'b0000000000100001111110011;
    rom[51693] = 25'b0000000000100001110101110;
    rom[51694] = 25'b0000000000100001101101001;
    rom[51695] = 25'b0000000000100001100100101;
    rom[51696] = 25'b0000000000100001011100000;
    rom[51697] = 25'b0000000000100001010011011;
    rom[51698] = 25'b0000000000100001001010110;
    rom[51699] = 25'b0000000000100001000010011;
    rom[51700] = 25'b0000000000100000111001110;
    rom[51701] = 25'b0000000000100000110001001;
    rom[51702] = 25'b0000000000100000101000100;
    rom[51703] = 25'b0000000000100000100000000;
    rom[51704] = 25'b0000000000100000010111011;
    rom[51705] = 25'b0000000000100000001110111;
    rom[51706] = 25'b0000000000100000000110010;
    rom[51707] = 25'b0000000000011111111101101;
    rom[51708] = 25'b0000000000011111110101001;
    rom[51709] = 25'b0000000000011111101100101;
    rom[51710] = 25'b0000000000011111100100000;
    rom[51711] = 25'b0000000000011111011011100;
    rom[51712] = 25'b0000000000011111010010111;
    rom[51713] = 25'b0000000000011111001010010;
    rom[51714] = 25'b0000000000011111000001110;
    rom[51715] = 25'b0000000000011110111001010;
    rom[51716] = 25'b0000000000011110110000110;
    rom[51717] = 25'b0000000000011110101000001;
    rom[51718] = 25'b0000000000011110011111101;
    rom[51719] = 25'b0000000000011110010111000;
    rom[51720] = 25'b0000000000011110001110100;
    rom[51721] = 25'b0000000000011110000110000;
    rom[51722] = 25'b0000000000011101111101100;
    rom[51723] = 25'b0000000000011101110101000;
    rom[51724] = 25'b0000000000011101101100100;
    rom[51725] = 25'b0000000000011101100011111;
    rom[51726] = 25'b0000000000011101011011011;
    rom[51727] = 25'b0000000000011101010010111;
    rom[51728] = 25'b0000000000011101001010011;
    rom[51729] = 25'b0000000000011101000001111;
    rom[51730] = 25'b0000000000011100111001010;
    rom[51731] = 25'b0000000000011100110000110;
    rom[51732] = 25'b0000000000011100101000010;
    rom[51733] = 25'b0000000000011100011111110;
    rom[51734] = 25'b0000000000011100010111010;
    rom[51735] = 25'b0000000000011100001110110;
    rom[51736] = 25'b0000000000011100000110010;
    rom[51737] = 25'b0000000000011011111101110;
    rom[51738] = 25'b0000000000011011110101010;
    rom[51739] = 25'b0000000000011011101100110;
    rom[51740] = 25'b0000000000011011100100010;
    rom[51741] = 25'b0000000000011011011011110;
    rom[51742] = 25'b0000000000011011010011011;
    rom[51743] = 25'b0000000000011011001010111;
    rom[51744] = 25'b0000000000011011000010011;
    rom[51745] = 25'b0000000000011010111001111;
    rom[51746] = 25'b0000000000011010110001100;
    rom[51747] = 25'b0000000000011010101001000;
    rom[51748] = 25'b0000000000011010100000100;
    rom[51749] = 25'b0000000000011010011000001;
    rom[51750] = 25'b0000000000011010001111101;
    rom[51751] = 25'b0000000000011010000111001;
    rom[51752] = 25'b0000000000011001111110110;
    rom[51753] = 25'b0000000000011001110110010;
    rom[51754] = 25'b0000000000011001101101110;
    rom[51755] = 25'b0000000000011001100101010;
    rom[51756] = 25'b0000000000011001011100111;
    rom[51757] = 25'b0000000000011001010100011;
    rom[51758] = 25'b0000000000011001001100000;
    rom[51759] = 25'b0000000000011001000011101;
    rom[51760] = 25'b0000000000011000111011001;
    rom[51761] = 25'b0000000000011000110010101;
    rom[51762] = 25'b0000000000011000101010010;
    rom[51763] = 25'b0000000000011000100001111;
    rom[51764] = 25'b0000000000011000011001011;
    rom[51765] = 25'b0000000000011000010001000;
    rom[51766] = 25'b0000000000011000001000100;
    rom[51767] = 25'b0000000000011000000000001;
    rom[51768] = 25'b0000000000010111110111110;
    rom[51769] = 25'b0000000000010111101111011;
    rom[51770] = 25'b0000000000010111100111000;
    rom[51771] = 25'b0000000000010111011110100;
    rom[51772] = 25'b0000000000010111010110001;
    rom[51773] = 25'b0000000000010111001101110;
    rom[51774] = 25'b0000000000010111000101011;
    rom[51775] = 25'b0000000000010110111100111;
    rom[51776] = 25'b0000000000010110110100100;
    rom[51777] = 25'b0000000000010110101100001;
    rom[51778] = 25'b0000000000010110100011110;
    rom[51779] = 25'b0000000000010110011011011;
    rom[51780] = 25'b0000000000010110010011000;
    rom[51781] = 25'b0000000000010110001010101;
    rom[51782] = 25'b0000000000010110000010010;
    rom[51783] = 25'b0000000000010101111001111;
    rom[51784] = 25'b0000000000010101110001100;
    rom[51785] = 25'b0000000000010101101001001;
    rom[51786] = 25'b0000000000010101100000111;
    rom[51787] = 25'b0000000000010101011000011;
    rom[51788] = 25'b0000000000010101010000001;
    rom[51789] = 25'b0000000000010101000111110;
    rom[51790] = 25'b0000000000010100111111011;
    rom[51791] = 25'b0000000000010100110111000;
    rom[51792] = 25'b0000000000010100101110101;
    rom[51793] = 25'b0000000000010100100110011;
    rom[51794] = 25'b0000000000010100011110001;
    rom[51795] = 25'b0000000000010100010101101;
    rom[51796] = 25'b0000000000010100001101011;
    rom[51797] = 25'b0000000000010100000101000;
    rom[51798] = 25'b0000000000010011111100110;
    rom[51799] = 25'b0000000000010011110100011;
    rom[51800] = 25'b0000000000010011101100001;
    rom[51801] = 25'b0000000000010011100011110;
    rom[51802] = 25'b0000000000010011011011100;
    rom[51803] = 25'b0000000000010011010011001;
    rom[51804] = 25'b0000000000010011001010111;
    rom[51805] = 25'b0000000000010011000010100;
    rom[51806] = 25'b0000000000010010111010010;
    rom[51807] = 25'b0000000000010010110001111;
    rom[51808] = 25'b0000000000010010101001101;
    rom[51809] = 25'b0000000000010010100001011;
    rom[51810] = 25'b0000000000010010011001001;
    rom[51811] = 25'b0000000000010010010000110;
    rom[51812] = 25'b0000000000010010001000100;
    rom[51813] = 25'b0000000000010010000000010;
    rom[51814] = 25'b0000000000010001110111111;
    rom[51815] = 25'b0000000000010001101111110;
    rom[51816] = 25'b0000000000010001100111011;
    rom[51817] = 25'b0000000000010001011111001;
    rom[51818] = 25'b0000000000010001010110111;
    rom[51819] = 25'b0000000000010001001110101;
    rom[51820] = 25'b0000000000010001000110011;
    rom[51821] = 25'b0000000000010000111110001;
    rom[51822] = 25'b0000000000010000110101111;
    rom[51823] = 25'b0000000000010000101101101;
    rom[51824] = 25'b0000000000010000100101100;
    rom[51825] = 25'b0000000000010000011101001;
    rom[51826] = 25'b0000000000010000010101000;
    rom[51827] = 25'b0000000000010000001100110;
    rom[51828] = 25'b0000000000010000000100100;
    rom[51829] = 25'b0000000000001111111100010;
    rom[51830] = 25'b0000000000001111110100001;
    rom[51831] = 25'b0000000000001111101011111;
    rom[51832] = 25'b0000000000001111100011101;
    rom[51833] = 25'b0000000000001111011011011;
    rom[51834] = 25'b0000000000001111010011010;
    rom[51835] = 25'b0000000000001111001011001;
    rom[51836] = 25'b0000000000001111000010111;
    rom[51837] = 25'b0000000000001110111010101;
    rom[51838] = 25'b0000000000001110110010011;
    rom[51839] = 25'b0000000000001110101010010;
    rom[51840] = 25'b0000000000001110100010001;
    rom[51841] = 25'b0000000000001110011001111;
    rom[51842] = 25'b0000000000001110010001110;
    rom[51843] = 25'b0000000000001110001001100;
    rom[51844] = 25'b0000000000001110000001011;
    rom[51845] = 25'b0000000000001101111001001;
    rom[51846] = 25'b0000000000001101110001000;
    rom[51847] = 25'b0000000000001101101000111;
    rom[51848] = 25'b0000000000001101100000110;
    rom[51849] = 25'b0000000000001101011000101;
    rom[51850] = 25'b0000000000001101010000100;
    rom[51851] = 25'b0000000000001101001000011;
    rom[51852] = 25'b0000000000001101000000010;
    rom[51853] = 25'b0000000000001100111000000;
    rom[51854] = 25'b0000000000001100101111111;
    rom[51855] = 25'b0000000000001100100111110;
    rom[51856] = 25'b0000000000001100011111101;
    rom[51857] = 25'b0000000000001100010111100;
    rom[51858] = 25'b0000000000001100001111011;
    rom[51859] = 25'b0000000000001100000111010;
    rom[51860] = 25'b0000000000001011111111010;
    rom[51861] = 25'b0000000000001011110111001;
    rom[51862] = 25'b0000000000001011101111000;
    rom[51863] = 25'b0000000000001011100110111;
    rom[51864] = 25'b0000000000001011011110110;
    rom[51865] = 25'b0000000000001011010110101;
    rom[51866] = 25'b0000000000001011001110100;
    rom[51867] = 25'b0000000000001011000110100;
    rom[51868] = 25'b0000000000001010111110011;
    rom[51869] = 25'b0000000000001010110110011;
    rom[51870] = 25'b0000000000001010101110010;
    rom[51871] = 25'b0000000000001010100110010;
    rom[51872] = 25'b0000000000001010011110001;
    rom[51873] = 25'b0000000000001010010110000;
    rom[51874] = 25'b0000000000001010001110000;
    rom[51875] = 25'b0000000000001010000110000;
    rom[51876] = 25'b0000000000001001111110000;
    rom[51877] = 25'b0000000000001001110101111;
    rom[51878] = 25'b0000000000001001101101110;
    rom[51879] = 25'b0000000000001001100101110;
    rom[51880] = 25'b0000000000001001011101110;
    rom[51881] = 25'b0000000000001001010101110;
    rom[51882] = 25'b0000000000001001001101101;
    rom[51883] = 25'b0000000000001001000101101;
    rom[51884] = 25'b0000000000001000111101101;
    rom[51885] = 25'b0000000000001000110101101;
    rom[51886] = 25'b0000000000001000101101101;
    rom[51887] = 25'b0000000000001000100101101;
    rom[51888] = 25'b0000000000001000011101101;
    rom[51889] = 25'b0000000000001000010101101;
    rom[51890] = 25'b0000000000001000001101101;
    rom[51891] = 25'b0000000000001000000101101;
    rom[51892] = 25'b0000000000000111111101101;
    rom[51893] = 25'b0000000000000111110101110;
    rom[51894] = 25'b0000000000000111101101101;
    rom[51895] = 25'b0000000000000111100101110;
    rom[51896] = 25'b0000000000000111011101110;
    rom[51897] = 25'b0000000000000111010101110;
    rom[51898] = 25'b0000000000000111001101111;
    rom[51899] = 25'b0000000000000111000101111;
    rom[51900] = 25'b0000000000000110111110000;
    rom[51901] = 25'b0000000000000110110101111;
    rom[51902] = 25'b0000000000000110101110000;
    rom[51903] = 25'b0000000000000110100110000;
    rom[51904] = 25'b0000000000000110011110001;
    rom[51905] = 25'b0000000000000110010110001;
    rom[51906] = 25'b0000000000000110001110010;
    rom[51907] = 25'b0000000000000110000110011;
    rom[51908] = 25'b0000000000000101111110100;
    rom[51909] = 25'b0000000000000101110110100;
    rom[51910] = 25'b0000000000000101101110101;
    rom[51911] = 25'b0000000000000101100110110;
    rom[51912] = 25'b0000000000000101011110110;
    rom[51913] = 25'b0000000000000101010110111;
    rom[51914] = 25'b0000000000000101001111000;
    rom[51915] = 25'b0000000000000101000111001;
    rom[51916] = 25'b0000000000000100111111010;
    rom[51917] = 25'b0000000000000100110111010;
    rom[51918] = 25'b0000000000000100101111100;
    rom[51919] = 25'b0000000000000100100111101;
    rom[51920] = 25'b0000000000000100011111101;
    rom[51921] = 25'b0000000000000100010111111;
    rom[51922] = 25'b0000000000000100010000000;
    rom[51923] = 25'b0000000000000100001000001;
    rom[51924] = 25'b0000000000000100000000010;
    rom[51925] = 25'b0000000000000011111000100;
    rom[51926] = 25'b0000000000000011110000101;
    rom[51927] = 25'b0000000000000011101000110;
    rom[51928] = 25'b0000000000000011100000111;
    rom[51929] = 25'b0000000000000011011001000;
    rom[51930] = 25'b0000000000000011010001010;
    rom[51931] = 25'b0000000000000011001001011;
    rom[51932] = 25'b0000000000000011000001101;
    rom[51933] = 25'b0000000000000010111001110;
    rom[51934] = 25'b0000000000000010110001111;
    rom[51935] = 25'b0000000000000010101010001;
    rom[51936] = 25'b0000000000000010100010011;
    rom[51937] = 25'b0000000000000010011010101;
    rom[51938] = 25'b0000000000000010010010110;
    rom[51939] = 25'b0000000000000010001011000;
    rom[51940] = 25'b0000000000000010000011010;
    rom[51941] = 25'b0000000000000001111011011;
    rom[51942] = 25'b0000000000000001110011101;
    rom[51943] = 25'b0000000000000001101011111;
    rom[51944] = 25'b0000000000000001100100001;
    rom[51945] = 25'b0000000000000001011100011;
    rom[51946] = 25'b0000000000000001010100101;
    rom[51947] = 25'b0000000000000001001100111;
    rom[51948] = 25'b0000000000000001000101001;
    rom[51949] = 25'b0000000000000000111101011;
    rom[51950] = 25'b0000000000000000110101101;
    rom[51951] = 25'b0000000000000000101101111;
    rom[51952] = 25'b0000000000000000100110001;
    rom[51953] = 25'b0000000000000000011110100;
    rom[51954] = 25'b0000000000000000010110110;
    rom[51955] = 25'b0000000000000000001111000;
    rom[51956] = 25'b0000000000000000000111011;
    rom[51957] = 25'b1111111111111111111111101;
    rom[51958] = 25'b1111111111111111111000000;
    rom[51959] = 25'b1111111111111111110000010;
    rom[51960] = 25'b1111111111111111101000101;
    rom[51961] = 25'b1111111111111111100000111;
    rom[51962] = 25'b1111111111111111011001001;
    rom[51963] = 25'b1111111111111111010001100;
    rom[51964] = 25'b1111111111111111001001111;
    rom[51965] = 25'b1111111111111111000010010;
    rom[51966] = 25'b1111111111111110111010100;
    rom[51967] = 25'b1111111111111110110010111;
    rom[51968] = 25'b1111111111111110101011010;
    rom[51969] = 25'b1111111111111110100011101;
    rom[51970] = 25'b1111111111111110011011111;
    rom[51971] = 25'b1111111111111110010100010;
    rom[51972] = 25'b1111111111111110001100101;
    rom[51973] = 25'b1111111111111110000101000;
    rom[51974] = 25'b1111111111111101111101011;
    rom[51975] = 25'b1111111111111101110101110;
    rom[51976] = 25'b1111111111111101101110001;
    rom[51977] = 25'b1111111111111101100110100;
    rom[51978] = 25'b1111111111111101011111000;
    rom[51979] = 25'b1111111111111101010111010;
    rom[51980] = 25'b1111111111111101001111110;
    rom[51981] = 25'b1111111111111101001000001;
    rom[51982] = 25'b1111111111111101000000100;
    rom[51983] = 25'b1111111111111100111000111;
    rom[51984] = 25'b1111111111111100110001011;
    rom[51985] = 25'b1111111111111100101001110;
    rom[51986] = 25'b1111111111111100100010010;
    rom[51987] = 25'b1111111111111100011010101;
    rom[51988] = 25'b1111111111111100010011001;
    rom[51989] = 25'b1111111111111100001011100;
    rom[51990] = 25'b1111111111111100000100000;
    rom[51991] = 25'b1111111111111011111100011;
    rom[51992] = 25'b1111111111111011110101000;
    rom[51993] = 25'b1111111111111011101101011;
    rom[51994] = 25'b1111111111111011100101111;
    rom[51995] = 25'b1111111111111011011110011;
    rom[51996] = 25'b1111111111111011010110110;
    rom[51997] = 25'b1111111111111011001111010;
    rom[51998] = 25'b1111111111111011000111110;
    rom[51999] = 25'b1111111111111011000000010;
    rom[52000] = 25'b1111111111111010111000110;
    rom[52001] = 25'b1111111111111010110001010;
    rom[52002] = 25'b1111111111111010101001110;
    rom[52003] = 25'b1111111111111010100010010;
    rom[52004] = 25'b1111111111111010011010111;
    rom[52005] = 25'b1111111111111010010011011;
    rom[52006] = 25'b1111111111111010001011111;
    rom[52007] = 25'b1111111111111010000100011;
    rom[52008] = 25'b1111111111111001111101000;
    rom[52009] = 25'b1111111111111001110101100;
    rom[52010] = 25'b1111111111111001101110000;
    rom[52011] = 25'b1111111111111001100110101;
    rom[52012] = 25'b1111111111111001011111001;
    rom[52013] = 25'b1111111111111001010111101;
    rom[52014] = 25'b1111111111111001010000010;
    rom[52015] = 25'b1111111111111001001000111;
    rom[52016] = 25'b1111111111111001000001100;
    rom[52017] = 25'b1111111111111000111010000;
    rom[52018] = 25'b1111111111111000110010101;
    rom[52019] = 25'b1111111111111000101011010;
    rom[52020] = 25'b1111111111111000100011110;
    rom[52021] = 25'b1111111111111000011100011;
    rom[52022] = 25'b1111111111111000010101000;
    rom[52023] = 25'b1111111111111000001101101;
    rom[52024] = 25'b1111111111111000000110010;
    rom[52025] = 25'b1111111111110111111110111;
    rom[52026] = 25'b1111111111110111110111100;
    rom[52027] = 25'b1111111111110111110000001;
    rom[52028] = 25'b1111111111110111101000110;
    rom[52029] = 25'b1111111111110111100001100;
    rom[52030] = 25'b1111111111110111011010001;
    rom[52031] = 25'b1111111111110111010010110;
    rom[52032] = 25'b1111111111110111001011011;
    rom[52033] = 25'b1111111111110111000100000;
    rom[52034] = 25'b1111111111110110111100110;
    rom[52035] = 25'b1111111111110110110101011;
    rom[52036] = 25'b1111111111110110101110001;
    rom[52037] = 25'b1111111111110110100110110;
    rom[52038] = 25'b1111111111110110011111011;
    rom[52039] = 25'b1111111111110110011000001;
    rom[52040] = 25'b1111111111110110010000111;
    rom[52041] = 25'b1111111111110110001001101;
    rom[52042] = 25'b1111111111110110000010010;
    rom[52043] = 25'b1111111111110101111011000;
    rom[52044] = 25'b1111111111110101110011110;
    rom[52045] = 25'b1111111111110101101100100;
    rom[52046] = 25'b1111111111110101100101001;
    rom[52047] = 25'b1111111111110101011110000;
    rom[52048] = 25'b1111111111110101010110101;
    rom[52049] = 25'b1111111111110101001111011;
    rom[52050] = 25'b1111111111110101001000010;
    rom[52051] = 25'b1111111111110101000000111;
    rom[52052] = 25'b1111111111110100111001110;
    rom[52053] = 25'b1111111111110100110010100;
    rom[52054] = 25'b1111111111110100101011010;
    rom[52055] = 25'b1111111111110100100100001;
    rom[52056] = 25'b1111111111110100011100110;
    rom[52057] = 25'b1111111111110100010101101;
    rom[52058] = 25'b1111111111110100001110011;
    rom[52059] = 25'b1111111111110100000111010;
    rom[52060] = 25'b1111111111110100000000000;
    rom[52061] = 25'b1111111111110011111000111;
    rom[52062] = 25'b1111111111110011110001101;
    rom[52063] = 25'b1111111111110011101010100;
    rom[52064] = 25'b1111111111110011100011011;
    rom[52065] = 25'b1111111111110011011100001;
    rom[52066] = 25'b1111111111110011010101000;
    rom[52067] = 25'b1111111111110011001101111;
    rom[52068] = 25'b1111111111110011000110101;
    rom[52069] = 25'b1111111111110010111111101;
    rom[52070] = 25'b1111111111110010111000011;
    rom[52071] = 25'b1111111111110010110001010;
    rom[52072] = 25'b1111111111110010101010001;
    rom[52073] = 25'b1111111111110010100011000;
    rom[52074] = 25'b1111111111110010011011111;
    rom[52075] = 25'b1111111111110010010100110;
    rom[52076] = 25'b1111111111110010001101110;
    rom[52077] = 25'b1111111111110010000110101;
    rom[52078] = 25'b1111111111110001111111100;
    rom[52079] = 25'b1111111111110001111000011;
    rom[52080] = 25'b1111111111110001110001011;
    rom[52081] = 25'b1111111111110001101010010;
    rom[52082] = 25'b1111111111110001100011010;
    rom[52083] = 25'b1111111111110001011100001;
    rom[52084] = 25'b1111111111110001010101000;
    rom[52085] = 25'b1111111111110001001110000;
    rom[52086] = 25'b1111111111110001000110111;
    rom[52087] = 25'b1111111111110000111111111;
    rom[52088] = 25'b1111111111110000111000111;
    rom[52089] = 25'b1111111111110000110001111;
    rom[52090] = 25'b1111111111110000101010111;
    rom[52091] = 25'b1111111111110000100011110;
    rom[52092] = 25'b1111111111110000011100110;
    rom[52093] = 25'b1111111111110000010101110;
    rom[52094] = 25'b1111111111110000001110110;
    rom[52095] = 25'b1111111111110000000111110;
    rom[52096] = 25'b1111111111110000000000110;
    rom[52097] = 25'b1111111111101111111001110;
    rom[52098] = 25'b1111111111101111110010110;
    rom[52099] = 25'b1111111111101111101011110;
    rom[52100] = 25'b1111111111101111100100111;
    rom[52101] = 25'b1111111111101111011101111;
    rom[52102] = 25'b1111111111101111010111000;
    rom[52103] = 25'b1111111111101111010000000;
    rom[52104] = 25'b1111111111101111001001000;
    rom[52105] = 25'b1111111111101111000010000;
    rom[52106] = 25'b1111111111101110111011001;
    rom[52107] = 25'b1111111111101110110100010;
    rom[52108] = 25'b1111111111101110101101010;
    rom[52109] = 25'b1111111111101110100110011;
    rom[52110] = 25'b1111111111101110011111100;
    rom[52111] = 25'b1111111111101110011000101;
    rom[52112] = 25'b1111111111101110010001101;
    rom[52113] = 25'b1111111111101110001010110;
    rom[52114] = 25'b1111111111101110000011111;
    rom[52115] = 25'b1111111111101101111100111;
    rom[52116] = 25'b1111111111101101110110001;
    rom[52117] = 25'b1111111111101101101111010;
    rom[52118] = 25'b1111111111101101101000011;
    rom[52119] = 25'b1111111111101101100001100;
    rom[52120] = 25'b1111111111101101011010101;
    rom[52121] = 25'b1111111111101101010011110;
    rom[52122] = 25'b1111111111101101001100111;
    rom[52123] = 25'b1111111111101101000110001;
    rom[52124] = 25'b1111111111101100111111010;
    rom[52125] = 25'b1111111111101100111000100;
    rom[52126] = 25'b1111111111101100110001101;
    rom[52127] = 25'b1111111111101100101010111;
    rom[52128] = 25'b1111111111101100100100000;
    rom[52129] = 25'b1111111111101100011101010;
    rom[52130] = 25'b1111111111101100010110011;
    rom[52131] = 25'b1111111111101100001111101;
    rom[52132] = 25'b1111111111101100001000111;
    rom[52133] = 25'b1111111111101100000010000;
    rom[52134] = 25'b1111111111101011111011010;
    rom[52135] = 25'b1111111111101011110100100;
    rom[52136] = 25'b1111111111101011101101110;
    rom[52137] = 25'b1111111111101011100111000;
    rom[52138] = 25'b1111111111101011100000010;
    rom[52139] = 25'b1111111111101011011001100;
    rom[52140] = 25'b1111111111101011010010110;
    rom[52141] = 25'b1111111111101011001100000;
    rom[52142] = 25'b1111111111101011000101010;
    rom[52143] = 25'b1111111111101010111110100;
    rom[52144] = 25'b1111111111101010110111111;
    rom[52145] = 25'b1111111111101010110001001;
    rom[52146] = 25'b1111111111101010101010011;
    rom[52147] = 25'b1111111111101010100011110;
    rom[52148] = 25'b1111111111101010011101001;
    rom[52149] = 25'b1111111111101010010110011;
    rom[52150] = 25'b1111111111101010001111101;
    rom[52151] = 25'b1111111111101010001001000;
    rom[52152] = 25'b1111111111101010000010011;
    rom[52153] = 25'b1111111111101001111011101;
    rom[52154] = 25'b1111111111101001110101000;
    rom[52155] = 25'b1111111111101001101110011;
    rom[52156] = 25'b1111111111101001100111110;
    rom[52157] = 25'b1111111111101001100001001;
    rom[52158] = 25'b1111111111101001011010100;
    rom[52159] = 25'b1111111111101001010011111;
    rom[52160] = 25'b1111111111101001001101010;
    rom[52161] = 25'b1111111111101001000110101;
    rom[52162] = 25'b1111111111101001000000000;
    rom[52163] = 25'b1111111111101000111001011;
    rom[52164] = 25'b1111111111101000110010110;
    rom[52165] = 25'b1111111111101000101100001;
    rom[52166] = 25'b1111111111101000100101101;
    rom[52167] = 25'b1111111111101000011111000;
    rom[52168] = 25'b1111111111101000011000100;
    rom[52169] = 25'b1111111111101000010001111;
    rom[52170] = 25'b1111111111101000001011010;
    rom[52171] = 25'b1111111111101000000100110;
    rom[52172] = 25'b1111111111100111111110010;
    rom[52173] = 25'b1111111111100111110111110;
    rom[52174] = 25'b1111111111100111110001001;
    rom[52175] = 25'b1111111111100111101010101;
    rom[52176] = 25'b1111111111100111100100001;
    rom[52177] = 25'b1111111111100111011101101;
    rom[52178] = 25'b1111111111100111010111001;
    rom[52179] = 25'b1111111111100111010000100;
    rom[52180] = 25'b1111111111100111001010001;
    rom[52181] = 25'b1111111111100111000011101;
    rom[52182] = 25'b1111111111100110111101001;
    rom[52183] = 25'b1111111111100110110110101;
    rom[52184] = 25'b1111111111100110110000001;
    rom[52185] = 25'b1111111111100110101001110;
    rom[52186] = 25'b1111111111100110100011010;
    rom[52187] = 25'b1111111111100110011100110;
    rom[52188] = 25'b1111111111100110010110010;
    rom[52189] = 25'b1111111111100110001111111;
    rom[52190] = 25'b1111111111100110001001100;
    rom[52191] = 25'b1111111111100110000011000;
    rom[52192] = 25'b1111111111100101111100101;
    rom[52193] = 25'b1111111111100101110110001;
    rom[52194] = 25'b1111111111100101101111110;
    rom[52195] = 25'b1111111111100101101001011;
    rom[52196] = 25'b1111111111100101100010111;
    rom[52197] = 25'b1111111111100101011100101;
    rom[52198] = 25'b1111111111100101010110010;
    rom[52199] = 25'b1111111111100101001111110;
    rom[52200] = 25'b1111111111100101001001011;
    rom[52201] = 25'b1111111111100101000011001;
    rom[52202] = 25'b1111111111100100111100110;
    rom[52203] = 25'b1111111111100100110110011;
    rom[52204] = 25'b1111111111100100110000000;
    rom[52205] = 25'b1111111111100100101001101;
    rom[52206] = 25'b1111111111100100100011011;
    rom[52207] = 25'b1111111111100100011101000;
    rom[52208] = 25'b1111111111100100010110101;
    rom[52209] = 25'b1111111111100100010000011;
    rom[52210] = 25'b1111111111100100001010000;
    rom[52211] = 25'b1111111111100100000011110;
    rom[52212] = 25'b1111111111100011111101011;
    rom[52213] = 25'b1111111111100011110111001;
    rom[52214] = 25'b1111111111100011110000111;
    rom[52215] = 25'b1111111111100011101010100;
    rom[52216] = 25'b1111111111100011100100010;
    rom[52217] = 25'b1111111111100011011110000;
    rom[52218] = 25'b1111111111100011010111110;
    rom[52219] = 25'b1111111111100011010001100;
    rom[52220] = 25'b1111111111100011001011010;
    rom[52221] = 25'b1111111111100011000101000;
    rom[52222] = 25'b1111111111100010111110111;
    rom[52223] = 25'b1111111111100010111000101;
    rom[52224] = 25'b1111111111100010110010011;
    rom[52225] = 25'b1111111111100010101100001;
    rom[52226] = 25'b1111111111100010100101111;
    rom[52227] = 25'b1111111111100010011111110;
    rom[52228] = 25'b1111111111100010011001100;
    rom[52229] = 25'b1111111111100010010011011;
    rom[52230] = 25'b1111111111100010001101001;
    rom[52231] = 25'b1111111111100010000111000;
    rom[52232] = 25'b1111111111100010000000111;
    rom[52233] = 25'b1111111111100001111010101;
    rom[52234] = 25'b1111111111100001110100100;
    rom[52235] = 25'b1111111111100001101110011;
    rom[52236] = 25'b1111111111100001101000001;
    rom[52237] = 25'b1111111111100001100010000;
    rom[52238] = 25'b1111111111100001011100000;
    rom[52239] = 25'b1111111111100001010101110;
    rom[52240] = 25'b1111111111100001001111110;
    rom[52241] = 25'b1111111111100001001001100;
    rom[52242] = 25'b1111111111100001000011100;
    rom[52243] = 25'b1111111111100000111101011;
    rom[52244] = 25'b1111111111100000110111010;
    rom[52245] = 25'b1111111111100000110001001;
    rom[52246] = 25'b1111111111100000101011001;
    rom[52247] = 25'b1111111111100000100101000;
    rom[52248] = 25'b1111111111100000011111000;
    rom[52249] = 25'b1111111111100000011000111;
    rom[52250] = 25'b1111111111100000010010111;
    rom[52251] = 25'b1111111111100000001100110;
    rom[52252] = 25'b1111111111100000000110110;
    rom[52253] = 25'b1111111111100000000000110;
    rom[52254] = 25'b1111111111011111111010101;
    rom[52255] = 25'b1111111111011111110100101;
    rom[52256] = 25'b1111111111011111101110101;
    rom[52257] = 25'b1111111111011111101000101;
    rom[52258] = 25'b1111111111011111100010101;
    rom[52259] = 25'b1111111111011111011100101;
    rom[52260] = 25'b1111111111011111010110101;
    rom[52261] = 25'b1111111111011111010000110;
    rom[52262] = 25'b1111111111011111001010110;
    rom[52263] = 25'b1111111111011111000100110;
    rom[52264] = 25'b1111111111011110111110110;
    rom[52265] = 25'b1111111111011110111000110;
    rom[52266] = 25'b1111111111011110110010111;
    rom[52267] = 25'b1111111111011110101101000;
    rom[52268] = 25'b1111111111011110100111000;
    rom[52269] = 25'b1111111111011110100001001;
    rom[52270] = 25'b1111111111011110011011001;
    rom[52271] = 25'b1111111111011110010101010;
    rom[52272] = 25'b1111111111011110001111011;
    rom[52273] = 25'b1111111111011110001001011;
    rom[52274] = 25'b1111111111011110000011100;
    rom[52275] = 25'b1111111111011101111101101;
    rom[52276] = 25'b1111111111011101110111110;
    rom[52277] = 25'b1111111111011101110001111;
    rom[52278] = 25'b1111111111011101101100000;
    rom[52279] = 25'b1111111111011101100110001;
    rom[52280] = 25'b1111111111011101100000010;
    rom[52281] = 25'b1111111111011101011010011;
    rom[52282] = 25'b1111111111011101010100101;
    rom[52283] = 25'b1111111111011101001110110;
    rom[52284] = 25'b1111111111011101001000111;
    rom[52285] = 25'b1111111111011101000011000;
    rom[52286] = 25'b1111111111011100111101010;
    rom[52287] = 25'b1111111111011100110111100;
    rom[52288] = 25'b1111111111011100110001101;
    rom[52289] = 25'b1111111111011100101011111;
    rom[52290] = 25'b1111111111011100100110001;
    rom[52291] = 25'b1111111111011100100000010;
    rom[52292] = 25'b1111111111011100011010100;
    rom[52293] = 25'b1111111111011100010100110;
    rom[52294] = 25'b1111111111011100001110111;
    rom[52295] = 25'b1111111111011100001001010;
    rom[52296] = 25'b1111111111011100000011100;
    rom[52297] = 25'b1111111111011011111101110;
    rom[52298] = 25'b1111111111011011111000000;
    rom[52299] = 25'b1111111111011011110010010;
    rom[52300] = 25'b1111111111011011101100100;
    rom[52301] = 25'b1111111111011011100110110;
    rom[52302] = 25'b1111111111011011100001001;
    rom[52303] = 25'b1111111111011011011011011;
    rom[52304] = 25'b1111111111011011010101101;
    rom[52305] = 25'b1111111111011011010000000;
    rom[52306] = 25'b1111111111011011001010010;
    rom[52307] = 25'b1111111111011011000100101;
    rom[52308] = 25'b1111111111011010111111000;
    rom[52309] = 25'b1111111111011010111001010;
    rom[52310] = 25'b1111111111011010110011110;
    rom[52311] = 25'b1111111111011010101110000;
    rom[52312] = 25'b1111111111011010101000011;
    rom[52313] = 25'b1111111111011010100010110;
    rom[52314] = 25'b1111111111011010011101001;
    rom[52315] = 25'b1111111111011010010111100;
    rom[52316] = 25'b1111111111011010010001111;
    rom[52317] = 25'b1111111111011010001100010;
    rom[52318] = 25'b1111111111011010000110101;
    rom[52319] = 25'b1111111111011010000001001;
    rom[52320] = 25'b1111111111011001111011100;
    rom[52321] = 25'b1111111111011001110101111;
    rom[52322] = 25'b1111111111011001110000011;
    rom[52323] = 25'b1111111111011001101010110;
    rom[52324] = 25'b1111111111011001100101001;
    rom[52325] = 25'b1111111111011001011111101;
    rom[52326] = 25'b1111111111011001011010001;
    rom[52327] = 25'b1111111111011001010100100;
    rom[52328] = 25'b1111111111011001001111000;
    rom[52329] = 25'b1111111111011001001001100;
    rom[52330] = 25'b1111111111011001000100000;
    rom[52331] = 25'b1111111111011000111110100;
    rom[52332] = 25'b1111111111011000111001000;
    rom[52333] = 25'b1111111111011000110011100;
    rom[52334] = 25'b1111111111011000101110000;
    rom[52335] = 25'b1111111111011000101000100;
    rom[52336] = 25'b1111111111011000100011000;
    rom[52337] = 25'b1111111111011000011101100;
    rom[52338] = 25'b1111111111011000011000001;
    rom[52339] = 25'b1111111111011000010010101;
    rom[52340] = 25'b1111111111011000001101001;
    rom[52341] = 25'b1111111111011000000111110;
    rom[52342] = 25'b1111111111011000000010010;
    rom[52343] = 25'b1111111111010111111100111;
    rom[52344] = 25'b1111111111010111110111011;
    rom[52345] = 25'b1111111111010111110010000;
    rom[52346] = 25'b1111111111010111101100101;
    rom[52347] = 25'b1111111111010111100111001;
    rom[52348] = 25'b1111111111010111100001111;
    rom[52349] = 25'b1111111111010111011100011;
    rom[52350] = 25'b1111111111010111010111000;
    rom[52351] = 25'b1111111111010111010001110;
    rom[52352] = 25'b1111111111010111001100010;
    rom[52353] = 25'b1111111111010111000111000;
    rom[52354] = 25'b1111111111010111000001100;
    rom[52355] = 25'b1111111111010110111100010;
    rom[52356] = 25'b1111111111010110110110111;
    rom[52357] = 25'b1111111111010110110001101;
    rom[52358] = 25'b1111111111010110101100010;
    rom[52359] = 25'b1111111111010110100110111;
    rom[52360] = 25'b1111111111010110100001101;
    rom[52361] = 25'b1111111111010110011100010;
    rom[52362] = 25'b1111111111010110010111000;
    rom[52363] = 25'b1111111111010110010001110;
    rom[52364] = 25'b1111111111010110001100011;
    rom[52365] = 25'b1111111111010110000111001;
    rom[52366] = 25'b1111111111010110000001111;
    rom[52367] = 25'b1111111111010101111100101;
    rom[52368] = 25'b1111111111010101110111011;
    rom[52369] = 25'b1111111111010101110010001;
    rom[52370] = 25'b1111111111010101101100111;
    rom[52371] = 25'b1111111111010101100111101;
    rom[52372] = 25'b1111111111010101100010011;
    rom[52373] = 25'b1111111111010101011101001;
    rom[52374] = 25'b1111111111010101011000000;
    rom[52375] = 25'b1111111111010101010010110;
    rom[52376] = 25'b1111111111010101001101100;
    rom[52377] = 25'b1111111111010101001000011;
    rom[52378] = 25'b1111111111010101000011001;
    rom[52379] = 25'b1111111111010100111110000;
    rom[52380] = 25'b1111111111010100111000111;
    rom[52381] = 25'b1111111111010100110011101;
    rom[52382] = 25'b1111111111010100101110100;
    rom[52383] = 25'b1111111111010100101001011;
    rom[52384] = 25'b1111111111010100100100001;
    rom[52385] = 25'b1111111111010100011111000;
    rom[52386] = 25'b1111111111010100011001111;
    rom[52387] = 25'b1111111111010100010100111;
    rom[52388] = 25'b1111111111010100001111110;
    rom[52389] = 25'b1111111111010100001010101;
    rom[52390] = 25'b1111111111010100000101100;
    rom[52391] = 25'b1111111111010100000000011;
    rom[52392] = 25'b1111111111010011111011010;
    rom[52393] = 25'b1111111111010011110110010;
    rom[52394] = 25'b1111111111010011110001010;
    rom[52395] = 25'b1111111111010011101100000;
    rom[52396] = 25'b1111111111010011100111000;
    rom[52397] = 25'b1111111111010011100010000;
    rom[52398] = 25'b1111111111010011011100111;
    rom[52399] = 25'b1111111111010011010111111;
    rom[52400] = 25'b1111111111010011010010111;
    rom[52401] = 25'b1111111111010011001101111;
    rom[52402] = 25'b1111111111010011001000111;
    rom[52403] = 25'b1111111111010011000011110;
    rom[52404] = 25'b1111111111010010111110111;
    rom[52405] = 25'b1111111111010010111001110;
    rom[52406] = 25'b1111111111010010110100111;
    rom[52407] = 25'b1111111111010010101111111;
    rom[52408] = 25'b1111111111010010101010111;
    rom[52409] = 25'b1111111111010010100101111;
    rom[52410] = 25'b1111111111010010100001000;
    rom[52411] = 25'b1111111111010010011100000;
    rom[52412] = 25'b1111111111010010010111001;
    rom[52413] = 25'b1111111111010010010010001;
    rom[52414] = 25'b1111111111010010001101001;
    rom[52415] = 25'b1111111111010010001000010;
    rom[52416] = 25'b1111111111010010000011011;
    rom[52417] = 25'b1111111111010001111110011;
    rom[52418] = 25'b1111111111010001111001100;
    rom[52419] = 25'b1111111111010001110100101;
    rom[52420] = 25'b1111111111010001101111110;
    rom[52421] = 25'b1111111111010001101010111;
    rom[52422] = 25'b1111111111010001100110000;
    rom[52423] = 25'b1111111111010001100001001;
    rom[52424] = 25'b1111111111010001011100010;
    rom[52425] = 25'b1111111111010001010111011;
    rom[52426] = 25'b1111111111010001010010101;
    rom[52427] = 25'b1111111111010001001101110;
    rom[52428] = 25'b1111111111010001001000111;
    rom[52429] = 25'b1111111111010001000100000;
    rom[52430] = 25'b1111111111010000111111010;
    rom[52431] = 25'b1111111111010000111010011;
    rom[52432] = 25'b1111111111010000110101101;
    rom[52433] = 25'b1111111111010000110000111;
    rom[52434] = 25'b1111111111010000101100000;
    rom[52435] = 25'b1111111111010000100111010;
    rom[52436] = 25'b1111111111010000100010100;
    rom[52437] = 25'b1111111111010000011101110;
    rom[52438] = 25'b1111111111010000011001000;
    rom[52439] = 25'b1111111111010000010100010;
    rom[52440] = 25'b1111111111010000001111100;
    rom[52441] = 25'b1111111111010000001010110;
    rom[52442] = 25'b1111111111010000000110000;
    rom[52443] = 25'b1111111111010000000001010;
    rom[52444] = 25'b1111111111001111111100101;
    rom[52445] = 25'b1111111111001111110111111;
    rom[52446] = 25'b1111111111001111110011001;
    rom[52447] = 25'b1111111111001111101110100;
    rom[52448] = 25'b1111111111001111101001110;
    rom[52449] = 25'b1111111111001111100101001;
    rom[52450] = 25'b1111111111001111100000011;
    rom[52451] = 25'b1111111111001111011011110;
    rom[52452] = 25'b1111111111001111010111001;
    rom[52453] = 25'b1111111111001111010010100;
    rom[52454] = 25'b1111111111001111001101111;
    rom[52455] = 25'b1111111111001111001001001;
    rom[52456] = 25'b1111111111001111000100101;
    rom[52457] = 25'b1111111111001110111111111;
    rom[52458] = 25'b1111111111001110111011011;
    rom[52459] = 25'b1111111111001110110110101;
    rom[52460] = 25'b1111111111001110110010001;
    rom[52461] = 25'b1111111111001110101101100;
    rom[52462] = 25'b1111111111001110101000111;
    rom[52463] = 25'b1111111111001110100100011;
    rom[52464] = 25'b1111111111001110011111110;
    rom[52465] = 25'b1111111111001110011011010;
    rom[52466] = 25'b1111111111001110010110101;
    rom[52467] = 25'b1111111111001110010010001;
    rom[52468] = 25'b1111111111001110001101101;
    rom[52469] = 25'b1111111111001110001001000;
    rom[52470] = 25'b1111111111001110000100100;
    rom[52471] = 25'b1111111111001110000000000;
    rom[52472] = 25'b1111111111001101111011100;
    rom[52473] = 25'b1111111111001101110111000;
    rom[52474] = 25'b1111111111001101110010100;
    rom[52475] = 25'b1111111111001101101110000;
    rom[52476] = 25'b1111111111001101101001100;
    rom[52477] = 25'b1111111111001101100101000;
    rom[52478] = 25'b1111111111001101100000100;
    rom[52479] = 25'b1111111111001101011100001;
    rom[52480] = 25'b1111111111001101010111101;
    rom[52481] = 25'b1111111111001101010011010;
    rom[52482] = 25'b1111111111001101001110110;
    rom[52483] = 25'b1111111111001101001010011;
    rom[52484] = 25'b1111111111001101000101111;
    rom[52485] = 25'b1111111111001101000001100;
    rom[52486] = 25'b1111111111001100111101001;
    rom[52487] = 25'b1111111111001100111000101;
    rom[52488] = 25'b1111111111001100110100010;
    rom[52489] = 25'b1111111111001100101111110;
    rom[52490] = 25'b1111111111001100101011100;
    rom[52491] = 25'b1111111111001100100111001;
    rom[52492] = 25'b1111111111001100100010110;
    rom[52493] = 25'b1111111111001100011110011;
    rom[52494] = 25'b1111111111001100011010000;
    rom[52495] = 25'b1111111111001100010101101;
    rom[52496] = 25'b1111111111001100010001011;
    rom[52497] = 25'b1111111111001100001101000;
    rom[52498] = 25'b1111111111001100001000101;
    rom[52499] = 25'b1111111111001100000100011;
    rom[52500] = 25'b1111111111001100000000001;
    rom[52501] = 25'b1111111111001011111011110;
    rom[52502] = 25'b1111111111001011110111100;
    rom[52503] = 25'b1111111111001011110011010;
    rom[52504] = 25'b1111111111001011101110111;
    rom[52505] = 25'b1111111111001011101010101;
    rom[52506] = 25'b1111111111001011100110011;
    rom[52507] = 25'b1111111111001011100010001;
    rom[52508] = 25'b1111111111001011011101111;
    rom[52509] = 25'b1111111111001011011001101;
    rom[52510] = 25'b1111111111001011010101011;
    rom[52511] = 25'b1111111111001011010001001;
    rom[52512] = 25'b1111111111001011001100111;
    rom[52513] = 25'b1111111111001011001000110;
    rom[52514] = 25'b1111111111001011000100100;
    rom[52515] = 25'b1111111111001011000000010;
    rom[52516] = 25'b1111111111001010111100001;
    rom[52517] = 25'b1111111111001010110111111;
    rom[52518] = 25'b1111111111001010110011110;
    rom[52519] = 25'b1111111111001010101111101;
    rom[52520] = 25'b1111111111001010101011011;
    rom[52521] = 25'b1111111111001010100111010;
    rom[52522] = 25'b1111111111001010100011001;
    rom[52523] = 25'b1111111111001010011111000;
    rom[52524] = 25'b1111111111001010011010111;
    rom[52525] = 25'b1111111111001010010110110;
    rom[52526] = 25'b1111111111001010010010101;
    rom[52527] = 25'b1111111111001010001110100;
    rom[52528] = 25'b1111111111001010001010011;
    rom[52529] = 25'b1111111111001010000110011;
    rom[52530] = 25'b1111111111001010000010010;
    rom[52531] = 25'b1111111111001001111110001;
    rom[52532] = 25'b1111111111001001111010001;
    rom[52533] = 25'b1111111111001001110110000;
    rom[52534] = 25'b1111111111001001110010000;
    rom[52535] = 25'b1111111111001001101101111;
    rom[52536] = 25'b1111111111001001101001111;
    rom[52537] = 25'b1111111111001001100101111;
    rom[52538] = 25'b1111111111001001100001110;
    rom[52539] = 25'b1111111111001001011101110;
    rom[52540] = 25'b1111111111001001011001110;
    rom[52541] = 25'b1111111111001001010101110;
    rom[52542] = 25'b1111111111001001010001110;
    rom[52543] = 25'b1111111111001001001101110;
    rom[52544] = 25'b1111111111001001001001110;
    rom[52545] = 25'b1111111111001001000101110;
    rom[52546] = 25'b1111111111001001000001110;
    rom[52547] = 25'b1111111111001000111101111;
    rom[52548] = 25'b1111111111001000111001111;
    rom[52549] = 25'b1111111111001000110101111;
    rom[52550] = 25'b1111111111001000110010000;
    rom[52551] = 25'b1111111111001000101110001;
    rom[52552] = 25'b1111111111001000101010001;
    rom[52553] = 25'b1111111111001000100110010;
    rom[52554] = 25'b1111111111001000100010010;
    rom[52555] = 25'b1111111111001000011110011;
    rom[52556] = 25'b1111111111001000011010100;
    rom[52557] = 25'b1111111111001000010110101;
    rom[52558] = 25'b1111111111001000010010110;
    rom[52559] = 25'b1111111111001000001110111;
    rom[52560] = 25'b1111111111001000001011000;
    rom[52561] = 25'b1111111111001000000111001;
    rom[52562] = 25'b1111111111001000000011010;
    rom[52563] = 25'b1111111111000111111111100;
    rom[52564] = 25'b1111111111000111111011101;
    rom[52565] = 25'b1111111111000111110111110;
    rom[52566] = 25'b1111111111000111110100000;
    rom[52567] = 25'b1111111111000111110000001;
    rom[52568] = 25'b1111111111000111101100011;
    rom[52569] = 25'b1111111111000111101000100;
    rom[52570] = 25'b1111111111000111100100110;
    rom[52571] = 25'b1111111111000111100000111;
    rom[52572] = 25'b1111111111000111011101010;
    rom[52573] = 25'b1111111111000111011001011;
    rom[52574] = 25'b1111111111000111010101101;
    rom[52575] = 25'b1111111111000111010001111;
    rom[52576] = 25'b1111111111000111001110001;
    rom[52577] = 25'b1111111111000111001010011;
    rom[52578] = 25'b1111111111000111000110101;
    rom[52579] = 25'b1111111111000111000011000;
    rom[52580] = 25'b1111111111000110111111010;
    rom[52581] = 25'b1111111111000110111011100;
    rom[52582] = 25'b1111111111000110110111111;
    rom[52583] = 25'b1111111111000110110100001;
    rom[52584] = 25'b1111111111000110110000100;
    rom[52585] = 25'b1111111111000110101100110;
    rom[52586] = 25'b1111111111000110101001001;
    rom[52587] = 25'b1111111111000110100101100;
    rom[52588] = 25'b1111111111000110100001110;
    rom[52589] = 25'b1111111111000110011110000;
    rom[52590] = 25'b1111111111000110011010011;
    rom[52591] = 25'b1111111111000110010110110;
    rom[52592] = 25'b1111111111000110010011001;
    rom[52593] = 25'b1111111111000110001111101;
    rom[52594] = 25'b1111111111000110001100000;
    rom[52595] = 25'b1111111111000110001000010;
    rom[52596] = 25'b1111111111000110000100110;
    rom[52597] = 25'b1111111111000110000001001;
    rom[52598] = 25'b1111111111000101111101100;
    rom[52599] = 25'b1111111111000101111010000;
    rom[52600] = 25'b1111111111000101110110011;
    rom[52601] = 25'b1111111111000101110010111;
    rom[52602] = 25'b1111111111000101101111010;
    rom[52603] = 25'b1111111111000101101011110;
    rom[52604] = 25'b1111111111000101101000001;
    rom[52605] = 25'b1111111111000101100100101;
    rom[52606] = 25'b1111111111000101100001001;
    rom[52607] = 25'b1111111111000101011101101;
    rom[52608] = 25'b1111111111000101011010001;
    rom[52609] = 25'b1111111111000101010110101;
    rom[52610] = 25'b1111111111000101010011001;
    rom[52611] = 25'b1111111111000101001111101;
    rom[52612] = 25'b1111111111000101001100001;
    rom[52613] = 25'b1111111111000101001000110;
    rom[52614] = 25'b1111111111000101000101010;
    rom[52615] = 25'b1111111111000101000001110;
    rom[52616] = 25'b1111111111000100111110011;
    rom[52617] = 25'b1111111111000100111010111;
    rom[52618] = 25'b1111111111000100110111011;
    rom[52619] = 25'b1111111111000100110100000;
    rom[52620] = 25'b1111111111000100110000101;
    rom[52621] = 25'b1111111111000100101101001;
    rom[52622] = 25'b1111111111000100101001110;
    rom[52623] = 25'b1111111111000100100110011;
    rom[52624] = 25'b1111111111000100100011000;
    rom[52625] = 25'b1111111111000100011111101;
    rom[52626] = 25'b1111111111000100011100010;
    rom[52627] = 25'b1111111111000100011000111;
    rom[52628] = 25'b1111111111000100010101100;
    rom[52629] = 25'b1111111111000100010010001;
    rom[52630] = 25'b1111111111000100001110110;
    rom[52631] = 25'b1111111111000100001011100;
    rom[52632] = 25'b1111111111000100001000001;
    rom[52633] = 25'b1111111111000100000100111;
    rom[52634] = 25'b1111111111000100000001100;
    rom[52635] = 25'b1111111111000011111110001;
    rom[52636] = 25'b1111111111000011111010111;
    rom[52637] = 25'b1111111111000011110111100;
    rom[52638] = 25'b1111111111000011110100010;
    rom[52639] = 25'b1111111111000011110001000;
    rom[52640] = 25'b1111111111000011101101110;
    rom[52641] = 25'b1111111111000011101010100;
    rom[52642] = 25'b1111111111000011100111010;
    rom[52643] = 25'b1111111111000011100100000;
    rom[52644] = 25'b1111111111000011100000110;
    rom[52645] = 25'b1111111111000011011101100;
    rom[52646] = 25'b1111111111000011011010010;
    rom[52647] = 25'b1111111111000011010111000;
    rom[52648] = 25'b1111111111000011010011111;
    rom[52649] = 25'b1111111111000011010000101;
    rom[52650] = 25'b1111111111000011001101011;
    rom[52651] = 25'b1111111111000011001010010;
    rom[52652] = 25'b1111111111000011000111001;
    rom[52653] = 25'b1111111111000011000011111;
    rom[52654] = 25'b1111111111000011000000110;
    rom[52655] = 25'b1111111111000010111101100;
    rom[52656] = 25'b1111111111000010111010011;
    rom[52657] = 25'b1111111111000010110111010;
    rom[52658] = 25'b1111111111000010110100001;
    rom[52659] = 25'b1111111111000010110001000;
    rom[52660] = 25'b1111111111000010101101111;
    rom[52661] = 25'b1111111111000010101010110;
    rom[52662] = 25'b1111111111000010100111110;
    rom[52663] = 25'b1111111111000010100100100;
    rom[52664] = 25'b1111111111000010100001100;
    rom[52665] = 25'b1111111111000010011110011;
    rom[52666] = 25'b1111111111000010011011010;
    rom[52667] = 25'b1111111111000010011000010;
    rom[52668] = 25'b1111111111000010010101010;
    rom[52669] = 25'b1111111111000010010010001;
    rom[52670] = 25'b1111111111000010001111000;
    rom[52671] = 25'b1111111111000010001100001;
    rom[52672] = 25'b1111111111000010001001000;
    rom[52673] = 25'b1111111111000010000110000;
    rom[52674] = 25'b1111111111000010000010111;
    rom[52675] = 25'b1111111111000001111111111;
    rom[52676] = 25'b1111111111000001111100111;
    rom[52677] = 25'b1111111111000001111010000;
    rom[52678] = 25'b1111111111000001110111000;
    rom[52679] = 25'b1111111111000001110100000;
    rom[52680] = 25'b1111111111000001110001000;
    rom[52681] = 25'b1111111111000001101110001;
    rom[52682] = 25'b1111111111000001101011001;
    rom[52683] = 25'b1111111111000001101000001;
    rom[52684] = 25'b1111111111000001100101010;
    rom[52685] = 25'b1111111111000001100010010;
    rom[52686] = 25'b1111111111000001011111011;
    rom[52687] = 25'b1111111111000001011100011;
    rom[52688] = 25'b1111111111000001011001100;
    rom[52689] = 25'b1111111111000001010110100;
    rom[52690] = 25'b1111111111000001010011101;
    rom[52691] = 25'b1111111111000001010000110;
    rom[52692] = 25'b1111111111000001001110000;
    rom[52693] = 25'b1111111111000001001011001;
    rom[52694] = 25'b1111111111000001001000001;
    rom[52695] = 25'b1111111111000001000101010;
    rom[52696] = 25'b1111111111000001000010100;
    rom[52697] = 25'b1111111111000000111111101;
    rom[52698] = 25'b1111111111000000111100110;
    rom[52699] = 25'b1111111111000000111010000;
    rom[52700] = 25'b1111111111000000110111001;
    rom[52701] = 25'b1111111111000000110100010;
    rom[52702] = 25'b1111111111000000110001100;
    rom[52703] = 25'b1111111111000000101110101;
    rom[52704] = 25'b1111111111000000101011111;
    rom[52705] = 25'b1111111111000000101001001;
    rom[52706] = 25'b1111111111000000100110011;
    rom[52707] = 25'b1111111111000000100011101;
    rom[52708] = 25'b1111111111000000100000110;
    rom[52709] = 25'b1111111111000000011110000;
    rom[52710] = 25'b1111111111000000011011010;
    rom[52711] = 25'b1111111111000000011000100;
    rom[52712] = 25'b1111111111000000010101111;
    rom[52713] = 25'b1111111111000000010011001;
    rom[52714] = 25'b1111111111000000010000011;
    rom[52715] = 25'b1111111111000000001101101;
    rom[52716] = 25'b1111111111000000001010111;
    rom[52717] = 25'b1111111111000000001000010;
    rom[52718] = 25'b1111111111000000000101101;
    rom[52719] = 25'b1111111111000000000010111;
    rom[52720] = 25'b1111111111000000000000001;
    rom[52721] = 25'b1111111110111111111101100;
    rom[52722] = 25'b1111111110111111111010111;
    rom[52723] = 25'b1111111110111111111000010;
    rom[52724] = 25'b1111111110111111110101101;
    rom[52725] = 25'b1111111110111111110010111;
    rom[52726] = 25'b1111111110111111110000010;
    rom[52727] = 25'b1111111110111111101101101;
    rom[52728] = 25'b1111111110111111101011001;
    rom[52729] = 25'b1111111110111111101000100;
    rom[52730] = 25'b1111111110111111100101111;
    rom[52731] = 25'b1111111110111111100011011;
    rom[52732] = 25'b1111111110111111100000110;
    rom[52733] = 25'b1111111110111111011110001;
    rom[52734] = 25'b1111111110111111011011100;
    rom[52735] = 25'b1111111110111111011001000;
    rom[52736] = 25'b1111111110111111010110011;
    rom[52737] = 25'b1111111110111111010011111;
    rom[52738] = 25'b1111111110111111010001010;
    rom[52739] = 25'b1111111110111111001110110;
    rom[52740] = 25'b1111111110111111001100010;
    rom[52741] = 25'b1111111110111111001001110;
    rom[52742] = 25'b1111111110111111000111010;
    rom[52743] = 25'b1111111110111111000100110;
    rom[52744] = 25'b1111111110111111000010010;
    rom[52745] = 25'b1111111110111110111111110;
    rom[52746] = 25'b1111111110111110111101010;
    rom[52747] = 25'b1111111110111110111010110;
    rom[52748] = 25'b1111111110111110111000011;
    rom[52749] = 25'b1111111110111110110101111;
    rom[52750] = 25'b1111111110111110110011011;
    rom[52751] = 25'b1111111110111110110001000;
    rom[52752] = 25'b1111111110111110101110100;
    rom[52753] = 25'b1111111110111110101100001;
    rom[52754] = 25'b1111111110111110101001110;
    rom[52755] = 25'b1111111110111110100111010;
    rom[52756] = 25'b1111111110111110100100111;
    rom[52757] = 25'b1111111110111110100010100;
    rom[52758] = 25'b1111111110111110100000001;
    rom[52759] = 25'b1111111110111110011101101;
    rom[52760] = 25'b1111111110111110011011010;
    rom[52761] = 25'b1111111110111110011001000;
    rom[52762] = 25'b1111111110111110010110100;
    rom[52763] = 25'b1111111110111110010100010;
    rom[52764] = 25'b1111111110111110010001111;
    rom[52765] = 25'b1111111110111110001111100;
    rom[52766] = 25'b1111111110111110001101010;
    rom[52767] = 25'b1111111110111110001010111;
    rom[52768] = 25'b1111111110111110001000100;
    rom[52769] = 25'b1111111110111110000110010;
    rom[52770] = 25'b1111111110111110000100000;
    rom[52771] = 25'b1111111110111110000001101;
    rom[52772] = 25'b1111111110111101111111011;
    rom[52773] = 25'b1111111110111101111101000;
    rom[52774] = 25'b1111111110111101111010111;
    rom[52775] = 25'b1111111110111101111000101;
    rom[52776] = 25'b1111111110111101110110010;
    rom[52777] = 25'b1111111110111101110100000;
    rom[52778] = 25'b1111111110111101110001110;
    rom[52779] = 25'b1111111110111101101111100;
    rom[52780] = 25'b1111111110111101101101010;
    rom[52781] = 25'b1111111110111101101011001;
    rom[52782] = 25'b1111111110111101101000111;
    rom[52783] = 25'b1111111110111101100110101;
    rom[52784] = 25'b1111111110111101100100100;
    rom[52785] = 25'b1111111110111101100010010;
    rom[52786] = 25'b1111111110111101100000001;
    rom[52787] = 25'b1111111110111101011101111;
    rom[52788] = 25'b1111111110111101011011110;
    rom[52789] = 25'b1111111110111101011001101;
    rom[52790] = 25'b1111111110111101010111011;
    rom[52791] = 25'b1111111110111101010101010;
    rom[52792] = 25'b1111111110111101010011001;
    rom[52793] = 25'b1111111110111101010001000;
    rom[52794] = 25'b1111111110111101001110111;
    rom[52795] = 25'b1111111110111101001100110;
    rom[52796] = 25'b1111111110111101001010101;
    rom[52797] = 25'b1111111110111101001000100;
    rom[52798] = 25'b1111111110111101000110011;
    rom[52799] = 25'b1111111110111101000100011;
    rom[52800] = 25'b1111111110111101000010010;
    rom[52801] = 25'b1111111110111101000000001;
    rom[52802] = 25'b1111111110111100111110001;
    rom[52803] = 25'b1111111110111100111100000;
    rom[52804] = 25'b1111111110111100111010000;
    rom[52805] = 25'b1111111110111100111000000;
    rom[52806] = 25'b1111111110111100110101111;
    rom[52807] = 25'b1111111110111100110011111;
    rom[52808] = 25'b1111111110111100110001111;
    rom[52809] = 25'b1111111110111100101111111;
    rom[52810] = 25'b1111111110111100101101111;
    rom[52811] = 25'b1111111110111100101011110;
    rom[52812] = 25'b1111111110111100101001111;
    rom[52813] = 25'b1111111110111100100111111;
    rom[52814] = 25'b1111111110111100100101111;
    rom[52815] = 25'b1111111110111100100011111;
    rom[52816] = 25'b1111111110111100100001111;
    rom[52817] = 25'b1111111110111100100000000;
    rom[52818] = 25'b1111111110111100011110000;
    rom[52819] = 25'b1111111110111100011100001;
    rom[52820] = 25'b1111111110111100011010001;
    rom[52821] = 25'b1111111110111100011000010;
    rom[52822] = 25'b1111111110111100010110011;
    rom[52823] = 25'b1111111110111100010100011;
    rom[52824] = 25'b1111111110111100010010100;
    rom[52825] = 25'b1111111110111100010000100;
    rom[52826] = 25'b1111111110111100001110101;
    rom[52827] = 25'b1111111110111100001100110;
    rom[52828] = 25'b1111111110111100001010111;
    rom[52829] = 25'b1111111110111100001001001;
    rom[52830] = 25'b1111111110111100000111010;
    rom[52831] = 25'b1111111110111100000101011;
    rom[52832] = 25'b1111111110111100000011100;
    rom[52833] = 25'b1111111110111100000001101;
    rom[52834] = 25'b1111111110111011111111111;
    rom[52835] = 25'b1111111110111011111110000;
    rom[52836] = 25'b1111111110111011111100001;
    rom[52837] = 25'b1111111110111011111010010;
    rom[52838] = 25'b1111111110111011111000100;
    rom[52839] = 25'b1111111110111011110110110;
    rom[52840] = 25'b1111111110111011110101000;
    rom[52841] = 25'b1111111110111011110011010;
    rom[52842] = 25'b1111111110111011110001100;
    rom[52843] = 25'b1111111110111011101111101;
    rom[52844] = 25'b1111111110111011101101111;
    rom[52845] = 25'b1111111110111011101100001;
    rom[52846] = 25'b1111111110111011101010011;
    rom[52847] = 25'b1111111110111011101000101;
    rom[52848] = 25'b1111111110111011100110111;
    rom[52849] = 25'b1111111110111011100101010;
    rom[52850] = 25'b1111111110111011100011011;
    rom[52851] = 25'b1111111110111011100001110;
    rom[52852] = 25'b1111111110111011100000001;
    rom[52853] = 25'b1111111110111011011110011;
    rom[52854] = 25'b1111111110111011011100101;
    rom[52855] = 25'b1111111110111011011010111;
    rom[52856] = 25'b1111111110111011011001011;
    rom[52857] = 25'b1111111110111011010111101;
    rom[52858] = 25'b1111111110111011010110000;
    rom[52859] = 25'b1111111110111011010100010;
    rom[52860] = 25'b1111111110111011010010110;
    rom[52861] = 25'b1111111110111011010001000;
    rom[52862] = 25'b1111111110111011001111100;
    rom[52863] = 25'b1111111110111011001101110;
    rom[52864] = 25'b1111111110111011001100001;
    rom[52865] = 25'b1111111110111011001010101;
    rom[52866] = 25'b1111111110111011001001000;
    rom[52867] = 25'b1111111110111011000111011;
    rom[52868] = 25'b1111111110111011000101111;
    rom[52869] = 25'b1111111110111011000100010;
    rom[52870] = 25'b1111111110111011000010101;
    rom[52871] = 25'b1111111110111011000001001;
    rom[52872] = 25'b1111111110111010111111100;
    rom[52873] = 25'b1111111110111010111110000;
    rom[52874] = 25'b1111111110111010111100011;
    rom[52875] = 25'b1111111110111010111010111;
    rom[52876] = 25'b1111111110111010111001011;
    rom[52877] = 25'b1111111110111010110111111;
    rom[52878] = 25'b1111111110111010110110011;
    rom[52879] = 25'b1111111110111010110100111;
    rom[52880] = 25'b1111111110111010110011011;
    rom[52881] = 25'b1111111110111010110001111;
    rom[52882] = 25'b1111111110111010110000011;
    rom[52883] = 25'b1111111110111010101110111;
    rom[52884] = 25'b1111111110111010101101011;
    rom[52885] = 25'b1111111110111010101100000;
    rom[52886] = 25'b1111111110111010101010100;
    rom[52887] = 25'b1111111110111010101001000;
    rom[52888] = 25'b1111111110111010100111101;
    rom[52889] = 25'b1111111110111010100110001;
    rom[52890] = 25'b1111111110111010100100101;
    rom[52891] = 25'b1111111110111010100011010;
    rom[52892] = 25'b1111111110111010100001111;
    rom[52893] = 25'b1111111110111010100000100;
    rom[52894] = 25'b1111111110111010011111001;
    rom[52895] = 25'b1111111110111010011101101;
    rom[52896] = 25'b1111111110111010011100010;
    rom[52897] = 25'b1111111110111010011010111;
    rom[52898] = 25'b1111111110111010011001101;
    rom[52899] = 25'b1111111110111010011000001;
    rom[52900] = 25'b1111111110111010010110111;
    rom[52901] = 25'b1111111110111010010101100;
    rom[52902] = 25'b1111111110111010010100001;
    rom[52903] = 25'b1111111110111010010010111;
    rom[52904] = 25'b1111111110111010010001100;
    rom[52905] = 25'b1111111110111010010000001;
    rom[52906] = 25'b1111111110111010001110111;
    rom[52907] = 25'b1111111110111010001101100;
    rom[52908] = 25'b1111111110111010001100010;
    rom[52909] = 25'b1111111110111010001010111;
    rom[52910] = 25'b1111111110111010001001110;
    rom[52911] = 25'b1111111110111010001000011;
    rom[52912] = 25'b1111111110111010000111001;
    rom[52913] = 25'b1111111110111010000101111;
    rom[52914] = 25'b1111111110111010000100100;
    rom[52915] = 25'b1111111110111010000011011;
    rom[52916] = 25'b1111111110111010000010001;
    rom[52917] = 25'b1111111110111010000000111;
    rom[52918] = 25'b1111111110111001111111101;
    rom[52919] = 25'b1111111110111001111110011;
    rom[52920] = 25'b1111111110111001111101001;
    rom[52921] = 25'b1111111110111001111100000;
    rom[52922] = 25'b1111111110111001111010110;
    rom[52923] = 25'b1111111110111001111001101;
    rom[52924] = 25'b1111111110111001111000011;
    rom[52925] = 25'b1111111110111001110111010;
    rom[52926] = 25'b1111111110111001110110001;
    rom[52927] = 25'b1111111110111001110100111;
    rom[52928] = 25'b1111111110111001110011110;
    rom[52929] = 25'b1111111110111001110010101;
    rom[52930] = 25'b1111111110111001110001011;
    rom[52931] = 25'b1111111110111001110000010;
    rom[52932] = 25'b1111111110111001101111001;
    rom[52933] = 25'b1111111110111001101110000;
    rom[52934] = 25'b1111111110111001101100111;
    rom[52935] = 25'b1111111110111001101011110;
    rom[52936] = 25'b1111111110111001101010110;
    rom[52937] = 25'b1111111110111001101001101;
    rom[52938] = 25'b1111111110111001101000100;
    rom[52939] = 25'b1111111110111001100111100;
    rom[52940] = 25'b1111111110111001100110011;
    rom[52941] = 25'b1111111110111001100101011;
    rom[52942] = 25'b1111111110111001100100010;
    rom[52943] = 25'b1111111110111001100011010;
    rom[52944] = 25'b1111111110111001100010001;
    rom[52945] = 25'b1111111110111001100001001;
    rom[52946] = 25'b1111111110111001100000001;
    rom[52947] = 25'b1111111110111001011111001;
    rom[52948] = 25'b1111111110111001011110001;
    rom[52949] = 25'b1111111110111001011101000;
    rom[52950] = 25'b1111111110111001011100000;
    rom[52951] = 25'b1111111110111001011011001;
    rom[52952] = 25'b1111111110111001011010000;
    rom[52953] = 25'b1111111110111001011001001;
    rom[52954] = 25'b1111111110111001011000001;
    rom[52955] = 25'b1111111110111001010111001;
    rom[52956] = 25'b1111111110111001010110010;
    rom[52957] = 25'b1111111110111001010101010;
    rom[52958] = 25'b1111111110111001010100010;
    rom[52959] = 25'b1111111110111001010011011;
    rom[52960] = 25'b1111111110111001010010011;
    rom[52961] = 25'b1111111110111001010001100;
    rom[52962] = 25'b1111111110111001010000101;
    rom[52963] = 25'b1111111110111001001111110;
    rom[52964] = 25'b1111111110111001001110110;
    rom[52965] = 25'b1111111110111001001101111;
    rom[52966] = 25'b1111111110111001001101000;
    rom[52967] = 25'b1111111110111001001100001;
    rom[52968] = 25'b1111111110111001001011010;
    rom[52969] = 25'b1111111110111001001010011;
    rom[52970] = 25'b1111111110111001001001100;
    rom[52971] = 25'b1111111110111001001000110;
    rom[52972] = 25'b1111111110111001000111110;
    rom[52973] = 25'b1111111110111001000110111;
    rom[52974] = 25'b1111111110111001000110001;
    rom[52975] = 25'b1111111110111001000101011;
    rom[52976] = 25'b1111111110111001000100100;
    rom[52977] = 25'b1111111110111001000011101;
    rom[52978] = 25'b1111111110111001000010111;
    rom[52979] = 25'b1111111110111001000010000;
    rom[52980] = 25'b1111111110111001000001010;
    rom[52981] = 25'b1111111110111001000000100;
    rom[52982] = 25'b1111111110111000111111110;
    rom[52983] = 25'b1111111110111000111110111;
    rom[52984] = 25'b1111111110111000111110001;
    rom[52985] = 25'b1111111110111000111101011;
    rom[52986] = 25'b1111111110111000111100101;
    rom[52987] = 25'b1111111110111000111011111;
    rom[52988] = 25'b1111111110111000111011001;
    rom[52989] = 25'b1111111110111000111010011;
    rom[52990] = 25'b1111111110111000111001110;
    rom[52991] = 25'b1111111110111000111001000;
    rom[52992] = 25'b1111111110111000111000010;
    rom[52993] = 25'b1111111110111000110111101;
    rom[52994] = 25'b1111111110111000110110111;
    rom[52995] = 25'b1111111110111000110110010;
    rom[52996] = 25'b1111111110111000110101100;
    rom[52997] = 25'b1111111110111000110100111;
    rom[52998] = 25'b1111111110111000110100001;
    rom[52999] = 25'b1111111110111000110011100;
    rom[53000] = 25'b1111111110111000110010111;
    rom[53001] = 25'b1111111110111000110010001;
    rom[53002] = 25'b1111111110111000110001101;
    rom[53003] = 25'b1111111110111000110001000;
    rom[53004] = 25'b1111111110111000110000011;
    rom[53005] = 25'b1111111110111000101111101;
    rom[53006] = 25'b1111111110111000101111001;
    rom[53007] = 25'b1111111110111000101110100;
    rom[53008] = 25'b1111111110111000101101111;
    rom[53009] = 25'b1111111110111000101101011;
    rom[53010] = 25'b1111111110111000101100101;
    rom[53011] = 25'b1111111110111000101100001;
    rom[53012] = 25'b1111111110111000101011100;
    rom[53013] = 25'b1111111110111000101011000;
    rom[53014] = 25'b1111111110111000101010011;
    rom[53015] = 25'b1111111110111000101001111;
    rom[53016] = 25'b1111111110111000101001010;
    rom[53017] = 25'b1111111110111000101000110;
    rom[53018] = 25'b1111111110111000101000010;
    rom[53019] = 25'b1111111110111000100111110;
    rom[53020] = 25'b1111111110111000100111010;
    rom[53021] = 25'b1111111110111000100110110;
    rom[53022] = 25'b1111111110111000100110010;
    rom[53023] = 25'b1111111110111000100101101;
    rom[53024] = 25'b1111111110111000100101010;
    rom[53025] = 25'b1111111110111000100100110;
    rom[53026] = 25'b1111111110111000100100010;
    rom[53027] = 25'b1111111110111000100011110;
    rom[53028] = 25'b1111111110111000100011011;
    rom[53029] = 25'b1111111110111000100010111;
    rom[53030] = 25'b1111111110111000100010011;
    rom[53031] = 25'b1111111110111000100001111;
    rom[53032] = 25'b1111111110111000100001100;
    rom[53033] = 25'b1111111110111000100001001;
    rom[53034] = 25'b1111111110111000100000110;
    rom[53035] = 25'b1111111110111000100000010;
    rom[53036] = 25'b1111111110111000011111111;
    rom[53037] = 25'b1111111110111000011111011;
    rom[53038] = 25'b1111111110111000011111000;
    rom[53039] = 25'b1111111110111000011110101;
    rom[53040] = 25'b1111111110111000011110010;
    rom[53041] = 25'b1111111110111000011101111;
    rom[53042] = 25'b1111111110111000011101100;
    rom[53043] = 25'b1111111110111000011101001;
    rom[53044] = 25'b1111111110111000011100110;
    rom[53045] = 25'b1111111110111000011100100;
    rom[53046] = 25'b1111111110111000011100001;
    rom[53047] = 25'b1111111110111000011011110;
    rom[53048] = 25'b1111111110111000011011100;
    rom[53049] = 25'b1111111110111000011011001;
    rom[53050] = 25'b1111111110111000011010111;
    rom[53051] = 25'b1111111110111000011010100;
    rom[53052] = 25'b1111111110111000011010010;
    rom[53053] = 25'b1111111110111000011001111;
    rom[53054] = 25'b1111111110111000011001101;
    rom[53055] = 25'b1111111110111000011001011;
    rom[53056] = 25'b1111111110111000011001001;
    rom[53057] = 25'b1111111110111000011000110;
    rom[53058] = 25'b1111111110111000011000101;
    rom[53059] = 25'b1111111110111000011000011;
    rom[53060] = 25'b1111111110111000011000000;
    rom[53061] = 25'b1111111110111000010111111;
    rom[53062] = 25'b1111111110111000010111101;
    rom[53063] = 25'b1111111110111000010111011;
    rom[53064] = 25'b1111111110111000010111001;
    rom[53065] = 25'b1111111110111000010110111;
    rom[53066] = 25'b1111111110111000010110110;
    rom[53067] = 25'b1111111110111000010110100;
    rom[53068] = 25'b1111111110111000010110011;
    rom[53069] = 25'b1111111110111000010110001;
    rom[53070] = 25'b1111111110111000010110000;
    rom[53071] = 25'b1111111110111000010101110;
    rom[53072] = 25'b1111111110111000010101101;
    rom[53073] = 25'b1111111110111000010101011;
    rom[53074] = 25'b1111111110111000010101010;
    rom[53075] = 25'b1111111110111000010101001;
    rom[53076] = 25'b1111111110111000010101000;
    rom[53077] = 25'b1111111110111000010100111;
    rom[53078] = 25'b1111111110111000010100110;
    rom[53079] = 25'b1111111110111000010100101;
    rom[53080] = 25'b1111111110111000010100100;
    rom[53081] = 25'b1111111110111000010100011;
    rom[53082] = 25'b1111111110111000010100010;
    rom[53083] = 25'b1111111110111000010100010;
    rom[53084] = 25'b1111111110111000010100001;
    rom[53085] = 25'b1111111110111000010100000;
    rom[53086] = 25'b1111111110111000010011111;
    rom[53087] = 25'b1111111110111000010011111;
    rom[53088] = 25'b1111111110111000010011111;
    rom[53089] = 25'b1111111110111000010011110;
    rom[53090] = 25'b1111111110111000010011101;
    rom[53091] = 25'b1111111110111000010011101;
    rom[53092] = 25'b1111111110111000010011101;
    rom[53093] = 25'b1111111110111000010011100;
    rom[53094] = 25'b1111111110111000010011100;
    rom[53095] = 25'b1111111110111000010011100;
    rom[53096] = 25'b1111111110111000010011100;
    rom[53097] = 25'b1111111110111000010011100;
    rom[53098] = 25'b1111111110111000010011100;
    rom[53099] = 25'b1111111110111000010011100;
    rom[53100] = 25'b1111111110111000010011100;
    rom[53101] = 25'b1111111110111000010011100;
    rom[53102] = 25'b1111111110111000010011100;
    rom[53103] = 25'b1111111110111000010011101;
    rom[53104] = 25'b1111111110111000010011101;
    rom[53105] = 25'b1111111110111000010011110;
    rom[53106] = 25'b1111111110111000010011110;
    rom[53107] = 25'b1111111110111000010011111;
    rom[53108] = 25'b1111111110111000010011111;
    rom[53109] = 25'b1111111110111000010100000;
    rom[53110] = 25'b1111111110111000010100000;
    rom[53111] = 25'b1111111110111000010100001;
    rom[53112] = 25'b1111111110111000010100010;
    rom[53113] = 25'b1111111110111000010100010;
    rom[53114] = 25'b1111111110111000010100011;
    rom[53115] = 25'b1111111110111000010100101;
    rom[53116] = 25'b1111111110111000010100101;
    rom[53117] = 25'b1111111110111000010100110;
    rom[53118] = 25'b1111111110111000010101000;
    rom[53119] = 25'b1111111110111000010101000;
    rom[53120] = 25'b1111111110111000010101010;
    rom[53121] = 25'b1111111110111000010101011;
    rom[53122] = 25'b1111111110111000010101100;
    rom[53123] = 25'b1111111110111000010101110;
    rom[53124] = 25'b1111111110111000010101111;
    rom[53125] = 25'b1111111110111000010110000;
    rom[53126] = 25'b1111111110111000010110001;
    rom[53127] = 25'b1111111110111000010110011;
    rom[53128] = 25'b1111111110111000010110101;
    rom[53129] = 25'b1111111110111000010110111;
    rom[53130] = 25'b1111111110111000010111000;
    rom[53131] = 25'b1111111110111000010111010;
    rom[53132] = 25'b1111111110111000010111100;
    rom[53133] = 25'b1111111110111000010111101;
    rom[53134] = 25'b1111111110111000011000000;
    rom[53135] = 25'b1111111110111000011000001;
    rom[53136] = 25'b1111111110111000011000011;
    rom[53137] = 25'b1111111110111000011000110;
    rom[53138] = 25'b1111111110111000011000111;
    rom[53139] = 25'b1111111110111000011001001;
    rom[53140] = 25'b1111111110111000011001011;
    rom[53141] = 25'b1111111110111000011001110;
    rom[53142] = 25'b1111111110111000011010000;
    rom[53143] = 25'b1111111110111000011010010;
    rom[53144] = 25'b1111111110111000011010100;
    rom[53145] = 25'b1111111110111000011010111;
    rom[53146] = 25'b1111111110111000011011010;
    rom[53147] = 25'b1111111110111000011011100;
    rom[53148] = 25'b1111111110111000011011111;
    rom[53149] = 25'b1111111110111000011100001;
    rom[53150] = 25'b1111111110111000011100100;
    rom[53151] = 25'b1111111110111000011100111;
    rom[53152] = 25'b1111111110111000011101001;
    rom[53153] = 25'b1111111110111000011101100;
    rom[53154] = 25'b1111111110111000011101111;
    rom[53155] = 25'b1111111110111000011110010;
    rom[53156] = 25'b1111111110111000011110101;
    rom[53157] = 25'b1111111110111000011111000;
    rom[53158] = 25'b1111111110111000011111011;
    rom[53159] = 25'b1111111110111000011111110;
    rom[53160] = 25'b1111111110111000100000001;
    rom[53161] = 25'b1111111110111000100000101;
    rom[53162] = 25'b1111111110111000100001000;
    rom[53163] = 25'b1111111110111000100001100;
    rom[53164] = 25'b1111111110111000100001111;
    rom[53165] = 25'b1111111110111000100010010;
    rom[53166] = 25'b1111111110111000100010101;
    rom[53167] = 25'b1111111110111000100011001;
    rom[53168] = 25'b1111111110111000100011101;
    rom[53169] = 25'b1111111110111000100100001;
    rom[53170] = 25'b1111111110111000100100100;
    rom[53171] = 25'b1111111110111000100101000;
    rom[53172] = 25'b1111111110111000100101100;
    rom[53173] = 25'b1111111110111000100110000;
    rom[53174] = 25'b1111111110111000100110011;
    rom[53175] = 25'b1111111110111000100110111;
    rom[53176] = 25'b1111111110111000100111100;
    rom[53177] = 25'b1111111110111000100111111;
    rom[53178] = 25'b1111111110111000101000100;
    rom[53179] = 25'b1111111110111000101001000;
    rom[53180] = 25'b1111111110111000101001100;
    rom[53181] = 25'b1111111110111000101010000;
    rom[53182] = 25'b1111111110111000101010100;
    rom[53183] = 25'b1111111110111000101011001;
    rom[53184] = 25'b1111111110111000101011101;
    rom[53185] = 25'b1111111110111000101100010;
    rom[53186] = 25'b1111111110111000101100110;
    rom[53187] = 25'b1111111110111000101101011;
    rom[53188] = 25'b1111111110111000101101111;
    rom[53189] = 25'b1111111110111000101110100;
    rom[53190] = 25'b1111111110111000101111000;
    rom[53191] = 25'b1111111110111000101111101;
    rom[53192] = 25'b1111111110111000110000010;
    rom[53193] = 25'b1111111110111000110000110;
    rom[53194] = 25'b1111111110111000110001011;
    rom[53195] = 25'b1111111110111000110010000;
    rom[53196] = 25'b1111111110111000110010101;
    rom[53197] = 25'b1111111110111000110011010;
    rom[53198] = 25'b1111111110111000110100000;
    rom[53199] = 25'b1111111110111000110100100;
    rom[53200] = 25'b1111111110111000110101001;
    rom[53201] = 25'b1111111110111000110101111;
    rom[53202] = 25'b1111111110111000110110100;
    rom[53203] = 25'b1111111110111000110111001;
    rom[53204] = 25'b1111111110111000110111111;
    rom[53205] = 25'b1111111110111000111000100;
    rom[53206] = 25'b1111111110111000111001010;
    rom[53207] = 25'b1111111110111000111001111;
    rom[53208] = 25'b1111111110111000111010101;
    rom[53209] = 25'b1111111110111000111011010;
    rom[53210] = 25'b1111111110111000111100000;
    rom[53211] = 25'b1111111110111000111100101;
    rom[53212] = 25'b1111111110111000111101011;
    rom[53213] = 25'b1111111110111000111110001;
    rom[53214] = 25'b1111111110111000111110111;
    rom[53215] = 25'b1111111110111000111111101;
    rom[53216] = 25'b1111111110111001000000011;
    rom[53217] = 25'b1111111110111001000001000;
    rom[53218] = 25'b1111111110111001000001111;
    rom[53219] = 25'b1111111110111001000010101;
    rom[53220] = 25'b1111111110111001000011011;
    rom[53221] = 25'b1111111110111001000100001;
    rom[53222] = 25'b1111111110111001000100111;
    rom[53223] = 25'b1111111110111001000101110;
    rom[53224] = 25'b1111111110111001000110100;
    rom[53225] = 25'b1111111110111001000111010;
    rom[53226] = 25'b1111111110111001001000000;
    rom[53227] = 25'b1111111110111001001000111;
    rom[53228] = 25'b1111111110111001001001110;
    rom[53229] = 25'b1111111110111001001010100;
    rom[53230] = 25'b1111111110111001001011010;
    rom[53231] = 25'b1111111110111001001100001;
    rom[53232] = 25'b1111111110111001001101000;
    rom[53233] = 25'b1111111110111001001101111;
    rom[53234] = 25'b1111111110111001001110101;
    rom[53235] = 25'b1111111110111001001111100;
    rom[53236] = 25'b1111111110111001010000100;
    rom[53237] = 25'b1111111110111001010001010;
    rom[53238] = 25'b1111111110111001010010001;
    rom[53239] = 25'b1111111110111001010011000;
    rom[53240] = 25'b1111111110111001010011111;
    rom[53241] = 25'b1111111110111001010100111;
    rom[53242] = 25'b1111111110111001010101101;
    rom[53243] = 25'b1111111110111001010110101;
    rom[53244] = 25'b1111111110111001010111100;
    rom[53245] = 25'b1111111110111001011000011;
    rom[53246] = 25'b1111111110111001011001011;
    rom[53247] = 25'b1111111110111001011010010;
    rom[53248] = 25'b1111111110111001011011001;
    rom[53249] = 25'b1111111110111001011100001;
    rom[53250] = 25'b1111111110111001011101000;
    rom[53251] = 25'b1111111110111001011110000;
    rom[53252] = 25'b1111111110111001011110111;
    rom[53253] = 25'b1111111110111001100000000;
    rom[53254] = 25'b1111111110111001100000111;
    rom[53255] = 25'b1111111110111001100001110;
    rom[53256] = 25'b1111111110111001100010111;
    rom[53257] = 25'b1111111110111001100011110;
    rom[53258] = 25'b1111111110111001100100110;
    rom[53259] = 25'b1111111110111001100101111;
    rom[53260] = 25'b1111111110111001100110110;
    rom[53261] = 25'b1111111110111001100111110;
    rom[53262] = 25'b1111111110111001101000111;
    rom[53263] = 25'b1111111110111001101001111;
    rom[53264] = 25'b1111111110111001101010111;
    rom[53265] = 25'b1111111110111001101011111;
    rom[53266] = 25'b1111111110111001101100111;
    rom[53267] = 25'b1111111110111001101110000;
    rom[53268] = 25'b1111111110111001101111000;
    rom[53269] = 25'b1111111110111001110000001;
    rom[53270] = 25'b1111111110111001110001001;
    rom[53271] = 25'b1111111110111001110010001;
    rom[53272] = 25'b1111111110111001110011010;
    rom[53273] = 25'b1111111110111001110100010;
    rom[53274] = 25'b1111111110111001110101011;
    rom[53275] = 25'b1111111110111001110110100;
    rom[53276] = 25'b1111111110111001110111101;
    rom[53277] = 25'b1111111110111001111000110;
    rom[53278] = 25'b1111111110111001111001110;
    rom[53279] = 25'b1111111110111001111010111;
    rom[53280] = 25'b1111111110111001111100000;
    rom[53281] = 25'b1111111110111001111101001;
    rom[53282] = 25'b1111111110111001111110010;
    rom[53283] = 25'b1111111110111001111111011;
    rom[53284] = 25'b1111111110111010000000100;
    rom[53285] = 25'b1111111110111010000001101;
    rom[53286] = 25'b1111111110111010000010110;
    rom[53287] = 25'b1111111110111010000100000;
    rom[53288] = 25'b1111111110111010000101001;
    rom[53289] = 25'b1111111110111010000110011;
    rom[53290] = 25'b1111111110111010000111100;
    rom[53291] = 25'b1111111110111010001000101;
    rom[53292] = 25'b1111111110111010001001110;
    rom[53293] = 25'b1111111110111010001011000;
    rom[53294] = 25'b1111111110111010001100010;
    rom[53295] = 25'b1111111110111010001101011;
    rom[53296] = 25'b1111111110111010001110101;
    rom[53297] = 25'b1111111110111010001111111;
    rom[53298] = 25'b1111111110111010010001001;
    rom[53299] = 25'b1111111110111010010010010;
    rom[53300] = 25'b1111111110111010010011100;
    rom[53301] = 25'b1111111110111010010100110;
    rom[53302] = 25'b1111111110111010010101111;
    rom[53303] = 25'b1111111110111010010111010;
    rom[53304] = 25'b1111111110111010011000100;
    rom[53305] = 25'b1111111110111010011001101;
    rom[53306] = 25'b1111111110111010011011000;
    rom[53307] = 25'b1111111110111010011100001;
    rom[53308] = 25'b1111111110111010011101100;
    rom[53309] = 25'b1111111110111010011110110;
    rom[53310] = 25'b1111111110111010100000000;
    rom[53311] = 25'b1111111110111010100001011;
    rom[53312] = 25'b1111111110111010100010101;
    rom[53313] = 25'b1111111110111010100011111;
    rom[53314] = 25'b1111111110111010100101010;
    rom[53315] = 25'b1111111110111010100110100;
    rom[53316] = 25'b1111111110111010100111111;
    rom[53317] = 25'b1111111110111010101001001;
    rom[53318] = 25'b1111111110111010101010100;
    rom[53319] = 25'b1111111110111010101011111;
    rom[53320] = 25'b1111111110111010101101001;
    rom[53321] = 25'b1111111110111010101110100;
    rom[53322] = 25'b1111111110111010101111111;
    rom[53323] = 25'b1111111110111010110001010;
    rom[53324] = 25'b1111111110111010110010101;
    rom[53325] = 25'b1111111110111010110100000;
    rom[53326] = 25'b1111111110111010110101010;
    rom[53327] = 25'b1111111110111010110110110;
    rom[53328] = 25'b1111111110111010111000001;
    rom[53329] = 25'b1111111110111010111001100;
    rom[53330] = 25'b1111111110111010111010111;
    rom[53331] = 25'b1111111110111010111100010;
    rom[53332] = 25'b1111111110111010111101101;
    rom[53333] = 25'b1111111110111010111111001;
    rom[53334] = 25'b1111111110111011000000100;
    rom[53335] = 25'b1111111110111011000001111;
    rom[53336] = 25'b1111111110111011000011010;
    rom[53337] = 25'b1111111110111011000100110;
    rom[53338] = 25'b1111111110111011000110010;
    rom[53339] = 25'b1111111110111011000111101;
    rom[53340] = 25'b1111111110111011001001001;
    rom[53341] = 25'b1111111110111011001010100;
    rom[53342] = 25'b1111111110111011001100000;
    rom[53343] = 25'b1111111110111011001101100;
    rom[53344] = 25'b1111111110111011001110111;
    rom[53345] = 25'b1111111110111011010000011;
    rom[53346] = 25'b1111111110111011010001111;
    rom[53347] = 25'b1111111110111011010011011;
    rom[53348] = 25'b1111111110111011010100111;
    rom[53349] = 25'b1111111110111011010110011;
    rom[53350] = 25'b1111111110111011010111111;
    rom[53351] = 25'b1111111110111011011001011;
    rom[53352] = 25'b1111111110111011011010111;
    rom[53353] = 25'b1111111110111011011100011;
    rom[53354] = 25'b1111111110111011011101111;
    rom[53355] = 25'b1111111110111011011111011;
    rom[53356] = 25'b1111111110111011100000111;
    rom[53357] = 25'b1111111110111011100010100;
    rom[53358] = 25'b1111111110111011100100000;
    rom[53359] = 25'b1111111110111011100101101;
    rom[53360] = 25'b1111111110111011100111001;
    rom[53361] = 25'b1111111110111011101000101;
    rom[53362] = 25'b1111111110111011101010010;
    rom[53363] = 25'b1111111110111011101011111;
    rom[53364] = 25'b1111111110111011101101011;
    rom[53365] = 25'b1111111110111011101110111;
    rom[53366] = 25'b1111111110111011110000100;
    rom[53367] = 25'b1111111110111011110010001;
    rom[53368] = 25'b1111111110111011110011101;
    rom[53369] = 25'b1111111110111011110101010;
    rom[53370] = 25'b1111111110111011110111000;
    rom[53371] = 25'b1111111110111011111000100;
    rom[53372] = 25'b1111111110111011111010001;
    rom[53373] = 25'b1111111110111011111011110;
    rom[53374] = 25'b1111111110111011111101011;
    rom[53375] = 25'b1111111110111011111111000;
    rom[53376] = 25'b1111111110111100000000101;
    rom[53377] = 25'b1111111110111100000010010;
    rom[53378] = 25'b1111111110111100000011111;
    rom[53379] = 25'b1111111110111100000101101;
    rom[53380] = 25'b1111111110111100000111010;
    rom[53381] = 25'b1111111110111100001000111;
    rom[53382] = 25'b1111111110111100001010100;
    rom[53383] = 25'b1111111110111100001100010;
    rom[53384] = 25'b1111111110111100001101111;
    rom[53385] = 25'b1111111110111100001111101;
    rom[53386] = 25'b1111111110111100010001010;
    rom[53387] = 25'b1111111110111100010011000;
    rom[53388] = 25'b1111111110111100010100101;
    rom[53389] = 25'b1111111110111100010110011;
    rom[53390] = 25'b1111111110111100011000001;
    rom[53391] = 25'b1111111110111100011001110;
    rom[53392] = 25'b1111111110111100011011100;
    rom[53393] = 25'b1111111110111100011101010;
    rom[53394] = 25'b1111111110111100011110111;
    rom[53395] = 25'b1111111110111100100000110;
    rom[53396] = 25'b1111111110111100100010100;
    rom[53397] = 25'b1111111110111100100100001;
    rom[53398] = 25'b1111111110111100100101111;
    rom[53399] = 25'b1111111110111100100111110;
    rom[53400] = 25'b1111111110111100101001100;
    rom[53401] = 25'b1111111110111100101011001;
    rom[53402] = 25'b1111111110111100101100111;
    rom[53403] = 25'b1111111110111100101110110;
    rom[53404] = 25'b1111111110111100110000100;
    rom[53405] = 25'b1111111110111100110010010;
    rom[53406] = 25'b1111111110111100110100001;
    rom[53407] = 25'b1111111110111100110101111;
    rom[53408] = 25'b1111111110111100110111101;
    rom[53409] = 25'b1111111110111100111001100;
    rom[53410] = 25'b1111111110111100111011010;
    rom[53411] = 25'b1111111110111100111101001;
    rom[53412] = 25'b1111111110111100111111000;
    rom[53413] = 25'b1111111110111101000000110;
    rom[53414] = 25'b1111111110111101000010101;
    rom[53415] = 25'b1111111110111101000100011;
    rom[53416] = 25'b1111111110111101000110010;
    rom[53417] = 25'b1111111110111101001000001;
    rom[53418] = 25'b1111111110111101001001111;
    rom[53419] = 25'b1111111110111101001011110;
    rom[53420] = 25'b1111111110111101001101101;
    rom[53421] = 25'b1111111110111101001111100;
    rom[53422] = 25'b1111111110111101010001011;
    rom[53423] = 25'b1111111110111101010011010;
    rom[53424] = 25'b1111111110111101010101001;
    rom[53425] = 25'b1111111110111101010111000;
    rom[53426] = 25'b1111111110111101011000111;
    rom[53427] = 25'b1111111110111101011010110;
    rom[53428] = 25'b1111111110111101011100101;
    rom[53429] = 25'b1111111110111101011110101;
    rom[53430] = 25'b1111111110111101100000100;
    rom[53431] = 25'b1111111110111101100010011;
    rom[53432] = 25'b1111111110111101100100010;
    rom[53433] = 25'b1111111110111101100110001;
    rom[53434] = 25'b1111111110111101101000001;
    rom[53435] = 25'b1111111110111101101010001;
    rom[53436] = 25'b1111111110111101101100000;
    rom[53437] = 25'b1111111110111101101101111;
    rom[53438] = 25'b1111111110111101101111111;
    rom[53439] = 25'b1111111110111101110001111;
    rom[53440] = 25'b1111111110111101110011110;
    rom[53441] = 25'b1111111110111101110101110;
    rom[53442] = 25'b1111111110111101110111110;
    rom[53443] = 25'b1111111110111101111001110;
    rom[53444] = 25'b1111111110111101111011101;
    rom[53445] = 25'b1111111110111101111101101;
    rom[53446] = 25'b1111111110111101111111101;
    rom[53447] = 25'b1111111110111110000001101;
    rom[53448] = 25'b1111111110111110000011101;
    rom[53449] = 25'b1111111110111110000101101;
    rom[53450] = 25'b1111111110111110000111101;
    rom[53451] = 25'b1111111110111110001001101;
    rom[53452] = 25'b1111111110111110001011101;
    rom[53453] = 25'b1111111110111110001101101;
    rom[53454] = 25'b1111111110111110001111101;
    rom[53455] = 25'b1111111110111110010001110;
    rom[53456] = 25'b1111111110111110010011110;
    rom[53457] = 25'b1111111110111110010101110;
    rom[53458] = 25'b1111111110111110010111110;
    rom[53459] = 25'b1111111110111110011001111;
    rom[53460] = 25'b1111111110111110011011111;
    rom[53461] = 25'b1111111110111110011101111;
    rom[53462] = 25'b1111111110111110100000000;
    rom[53463] = 25'b1111111110111110100010000;
    rom[53464] = 25'b1111111110111110100100001;
    rom[53465] = 25'b1111111110111110100110010;
    rom[53466] = 25'b1111111110111110101000010;
    rom[53467] = 25'b1111111110111110101010011;
    rom[53468] = 25'b1111111110111110101100011;
    rom[53469] = 25'b1111111110111110101110100;
    rom[53470] = 25'b1111111110111110110000101;
    rom[53471] = 25'b1111111110111110110010110;
    rom[53472] = 25'b1111111110111110110100110;
    rom[53473] = 25'b1111111110111110110111000;
    rom[53474] = 25'b1111111110111110111001001;
    rom[53475] = 25'b1111111110111110111011001;
    rom[53476] = 25'b1111111110111110111101010;
    rom[53477] = 25'b1111111110111110111111100;
    rom[53478] = 25'b1111111110111111000001101;
    rom[53479] = 25'b1111111110111111000011101;
    rom[53480] = 25'b1111111110111111000101110;
    rom[53481] = 25'b1111111110111111001000000;
    rom[53482] = 25'b1111111110111111001010001;
    rom[53483] = 25'b1111111110111111001100011;
    rom[53484] = 25'b1111111110111111001110100;
    rom[53485] = 25'b1111111110111111010000101;
    rom[53486] = 25'b1111111110111111010010110;
    rom[53487] = 25'b1111111110111111010100111;
    rom[53488] = 25'b1111111110111111010111001;
    rom[53489] = 25'b1111111110111111011001011;
    rom[53490] = 25'b1111111110111111011011100;
    rom[53491] = 25'b1111111110111111011101110;
    rom[53492] = 25'b1111111110111111011111111;
    rom[53493] = 25'b1111111110111111100010001;
    rom[53494] = 25'b1111111110111111100100011;
    rom[53495] = 25'b1111111110111111100110100;
    rom[53496] = 25'b1111111110111111101000110;
    rom[53497] = 25'b1111111110111111101011000;
    rom[53498] = 25'b1111111110111111101101010;
    rom[53499] = 25'b1111111110111111101111011;
    rom[53500] = 25'b1111111110111111110001101;
    rom[53501] = 25'b1111111110111111110011111;
    rom[53502] = 25'b1111111110111111110110001;
    rom[53503] = 25'b1111111110111111111000011;
    rom[53504] = 25'b1111111110111111111010101;
    rom[53505] = 25'b1111111110111111111100110;
    rom[53506] = 25'b1111111110111111111111001;
    rom[53507] = 25'b1111111111000000000001011;
    rom[53508] = 25'b1111111111000000000011101;
    rom[53509] = 25'b1111111111000000000101111;
    rom[53510] = 25'b1111111111000000001000010;
    rom[53511] = 25'b1111111111000000001010100;
    rom[53512] = 25'b1111111111000000001100110;
    rom[53513] = 25'b1111111111000000001111000;
    rom[53514] = 25'b1111111111000000010001011;
    rom[53515] = 25'b1111111111000000010011101;
    rom[53516] = 25'b1111111111000000010101111;
    rom[53517] = 25'b1111111111000000011000010;
    rom[53518] = 25'b1111111111000000011010100;
    rom[53519] = 25'b1111111111000000011100111;
    rom[53520] = 25'b1111111111000000011111001;
    rom[53521] = 25'b1111111111000000100001100;
    rom[53522] = 25'b1111111111000000100011111;
    rom[53523] = 25'b1111111111000000100110001;
    rom[53524] = 25'b1111111111000000101000100;
    rom[53525] = 25'b1111111111000000101010111;
    rom[53526] = 25'b1111111111000000101101001;
    rom[53527] = 25'b1111111111000000101111100;
    rom[53528] = 25'b1111111111000000110001111;
    rom[53529] = 25'b1111111111000000110100010;
    rom[53530] = 25'b1111111111000000110110101;
    rom[53531] = 25'b1111111111000000111001000;
    rom[53532] = 25'b1111111111000000111011011;
    rom[53533] = 25'b1111111111000000111101110;
    rom[53534] = 25'b1111111111000001000000001;
    rom[53535] = 25'b1111111111000001000010100;
    rom[53536] = 25'b1111111111000001000100111;
    rom[53537] = 25'b1111111111000001000111010;
    rom[53538] = 25'b1111111111000001001001101;
    rom[53539] = 25'b1111111111000001001100001;
    rom[53540] = 25'b1111111111000001001110011;
    rom[53541] = 25'b1111111111000001010000111;
    rom[53542] = 25'b1111111111000001010011010;
    rom[53543] = 25'b1111111111000001010101110;
    rom[53544] = 25'b1111111111000001011000001;
    rom[53545] = 25'b1111111111000001011010101;
    rom[53546] = 25'b1111111111000001011101000;
    rom[53547] = 25'b1111111111000001011111011;
    rom[53548] = 25'b1111111111000001100001111;
    rom[53549] = 25'b1111111111000001100100010;
    rom[53550] = 25'b1111111111000001100110110;
    rom[53551] = 25'b1111111111000001101001010;
    rom[53552] = 25'b1111111111000001101011101;
    rom[53553] = 25'b1111111111000001101110001;
    rom[53554] = 25'b1111111111000001110000101;
    rom[53555] = 25'b1111111111000001110011000;
    rom[53556] = 25'b1111111111000001110101100;
    rom[53557] = 25'b1111111111000001111000000;
    rom[53558] = 25'b1111111111000001111010100;
    rom[53559] = 25'b1111111111000001111100111;
    rom[53560] = 25'b1111111111000001111111100;
    rom[53561] = 25'b1111111111000010000010000;
    rom[53562] = 25'b1111111111000010000100011;
    rom[53563] = 25'b1111111111000010000110111;
    rom[53564] = 25'b1111111111000010001001100;
    rom[53565] = 25'b1111111111000010001100000;
    rom[53566] = 25'b1111111111000010001110100;
    rom[53567] = 25'b1111111111000010010001000;
    rom[53568] = 25'b1111111111000010010011100;
    rom[53569] = 25'b1111111111000010010110000;
    rom[53570] = 25'b1111111111000010011000101;
    rom[53571] = 25'b1111111111000010011011001;
    rom[53572] = 25'b1111111111000010011101101;
    rom[53573] = 25'b1111111111000010100000001;
    rom[53574] = 25'b1111111111000010100010101;
    rom[53575] = 25'b1111111111000010100101010;
    rom[53576] = 25'b1111111111000010100111110;
    rom[53577] = 25'b1111111111000010101010011;
    rom[53578] = 25'b1111111111000010101100111;
    rom[53579] = 25'b1111111111000010101111100;
    rom[53580] = 25'b1111111111000010110010001;
    rom[53581] = 25'b1111111111000010110100101;
    rom[53582] = 25'b1111111111000010110111010;
    rom[53583] = 25'b1111111111000010111001110;
    rom[53584] = 25'b1111111111000010111100011;
    rom[53585] = 25'b1111111111000010111111000;
    rom[53586] = 25'b1111111111000011000001101;
    rom[53587] = 25'b1111111111000011000100001;
    rom[53588] = 25'b1111111111000011000110110;
    rom[53589] = 25'b1111111111000011001001011;
    rom[53590] = 25'b1111111111000011001100000;
    rom[53591] = 25'b1111111111000011001110100;
    rom[53592] = 25'b1111111111000011010001001;
    rom[53593] = 25'b1111111111000011010011110;
    rom[53594] = 25'b1111111111000011010110011;
    rom[53595] = 25'b1111111111000011011001000;
    rom[53596] = 25'b1111111111000011011011101;
    rom[53597] = 25'b1111111111000011011110011;
    rom[53598] = 25'b1111111111000011100001000;
    rom[53599] = 25'b1111111111000011100011101;
    rom[53600] = 25'b1111111111000011100110010;
    rom[53601] = 25'b1111111111000011101000111;
    rom[53602] = 25'b1111111111000011101011100;
    rom[53603] = 25'b1111111111000011101110010;
    rom[53604] = 25'b1111111111000011110000111;
    rom[53605] = 25'b1111111111000011110011100;
    rom[53606] = 25'b1111111111000011110110001;
    rom[53607] = 25'b1111111111000011111000111;
    rom[53608] = 25'b1111111111000011111011101;
    rom[53609] = 25'b1111111111000011111110001;
    rom[53610] = 25'b1111111111000100000000111;
    rom[53611] = 25'b1111111111000100000011101;
    rom[53612] = 25'b1111111111000100000110010;
    rom[53613] = 25'b1111111111000100001001000;
    rom[53614] = 25'b1111111111000100001011101;
    rom[53615] = 25'b1111111111000100001110011;
    rom[53616] = 25'b1111111111000100010001000;
    rom[53617] = 25'b1111111111000100010011110;
    rom[53618] = 25'b1111111111000100010110100;
    rom[53619] = 25'b1111111111000100011001010;
    rom[53620] = 25'b1111111111000100011100000;
    rom[53621] = 25'b1111111111000100011110101;
    rom[53622] = 25'b1111111111000100100001011;
    rom[53623] = 25'b1111111111000100100100001;
    rom[53624] = 25'b1111111111000100100110111;
    rom[53625] = 25'b1111111111000100101001101;
    rom[53626] = 25'b1111111111000100101100011;
    rom[53627] = 25'b1111111111000100101111001;
    rom[53628] = 25'b1111111111000100110001111;
    rom[53629] = 25'b1111111111000100110100101;
    rom[53630] = 25'b1111111111000100110111011;
    rom[53631] = 25'b1111111111000100111010001;
    rom[53632] = 25'b1111111111000100111101000;
    rom[53633] = 25'b1111111111000100111111101;
    rom[53634] = 25'b1111111111000101000010100;
    rom[53635] = 25'b1111111111000101000101010;
    rom[53636] = 25'b1111111111000101001000000;
    rom[53637] = 25'b1111111111000101001010110;
    rom[53638] = 25'b1111111111000101001101100;
    rom[53639] = 25'b1111111111000101010000011;
    rom[53640] = 25'b1111111111000101010011001;
    rom[53641] = 25'b1111111111000101010110000;
    rom[53642] = 25'b1111111111000101011000110;
    rom[53643] = 25'b1111111111000101011011101;
    rom[53644] = 25'b1111111111000101011110011;
    rom[53645] = 25'b1111111111000101100001001;
    rom[53646] = 25'b1111111111000101100100000;
    rom[53647] = 25'b1111111111000101100110110;
    rom[53648] = 25'b1111111111000101101001101;
    rom[53649] = 25'b1111111111000101101100100;
    rom[53650] = 25'b1111111111000101101111010;
    rom[53651] = 25'b1111111111000101110010001;
    rom[53652] = 25'b1111111111000101110101000;
    rom[53653] = 25'b1111111111000101110111110;
    rom[53654] = 25'b1111111111000101111010101;
    rom[53655] = 25'b1111111111000101111101100;
    rom[53656] = 25'b1111111111000110000000011;
    rom[53657] = 25'b1111111111000110000011001;
    rom[53658] = 25'b1111111111000110000110000;
    rom[53659] = 25'b1111111111000110001001000;
    rom[53660] = 25'b1111111111000110001011110;
    rom[53661] = 25'b1111111111000110001110101;
    rom[53662] = 25'b1111111111000110010001100;
    rom[53663] = 25'b1111111111000110010100100;
    rom[53664] = 25'b1111111111000110010111010;
    rom[53665] = 25'b1111111111000110011010001;
    rom[53666] = 25'b1111111111000110011101000;
    rom[53667] = 25'b1111111111000110011111111;
    rom[53668] = 25'b1111111111000110100010111;
    rom[53669] = 25'b1111111111000110100101110;
    rom[53670] = 25'b1111111111000110101000101;
    rom[53671] = 25'b1111111111000110101011100;
    rom[53672] = 25'b1111111111000110101110011;
    rom[53673] = 25'b1111111111000110110001010;
    rom[53674] = 25'b1111111111000110110100010;
    rom[53675] = 25'b1111111111000110110111001;
    rom[53676] = 25'b1111111111000110111010001;
    rom[53677] = 25'b1111111111000110111101000;
    rom[53678] = 25'b1111111111000111000000000;
    rom[53679] = 25'b1111111111000111000010111;
    rom[53680] = 25'b1111111111000111000101111;
    rom[53681] = 25'b1111111111000111001000110;
    rom[53682] = 25'b1111111111000111001011101;
    rom[53683] = 25'b1111111111000111001110101;
    rom[53684] = 25'b1111111111000111010001101;
    rom[53685] = 25'b1111111111000111010100100;
    rom[53686] = 25'b1111111111000111010111100;
    rom[53687] = 25'b1111111111000111011010011;
    rom[53688] = 25'b1111111111000111011101011;
    rom[53689] = 25'b1111111111000111100000011;
    rom[53690] = 25'b1111111111000111100011011;
    rom[53691] = 25'b1111111111000111100110010;
    rom[53692] = 25'b1111111111000111101001010;
    rom[53693] = 25'b1111111111000111101100010;
    rom[53694] = 25'b1111111111000111101111010;
    rom[53695] = 25'b1111111111000111110010010;
    rom[53696] = 25'b1111111111000111110101010;
    rom[53697] = 25'b1111111111000111111000001;
    rom[53698] = 25'b1111111111000111111011001;
    rom[53699] = 25'b1111111111000111111110001;
    rom[53700] = 25'b1111111111001000000001001;
    rom[53701] = 25'b1111111111001000000100001;
    rom[53702] = 25'b1111111111001000000111001;
    rom[53703] = 25'b1111111111001000001010010;
    rom[53704] = 25'b1111111111001000001101010;
    rom[53705] = 25'b1111111111001000010000001;
    rom[53706] = 25'b1111111111001000010011001;
    rom[53707] = 25'b1111111111001000010110010;
    rom[53708] = 25'b1111111111001000011001010;
    rom[53709] = 25'b1111111111001000011100011;
    rom[53710] = 25'b1111111111001000011111010;
    rom[53711] = 25'b1111111111001000100010011;
    rom[53712] = 25'b1111111111001000100101011;
    rom[53713] = 25'b1111111111001000101000100;
    rom[53714] = 25'b1111111111001000101011100;
    rom[53715] = 25'b1111111111001000101110100;
    rom[53716] = 25'b1111111111001000110001100;
    rom[53717] = 25'b1111111111001000110100101;
    rom[53718] = 25'b1111111111001000110111101;
    rom[53719] = 25'b1111111111001000111010110;
    rom[53720] = 25'b1111111111001000111101110;
    rom[53721] = 25'b1111111111001001000000111;
    rom[53722] = 25'b1111111111001001000011111;
    rom[53723] = 25'b1111111111001001000111000;
    rom[53724] = 25'b1111111111001001001010001;
    rom[53725] = 25'b1111111111001001001101001;
    rom[53726] = 25'b1111111111001001010000010;
    rom[53727] = 25'b1111111111001001010011011;
    rom[53728] = 25'b1111111111001001010110011;
    rom[53729] = 25'b1111111111001001011001100;
    rom[53730] = 25'b1111111111001001011100101;
    rom[53731] = 25'b1111111111001001011111101;
    rom[53732] = 25'b1111111111001001100010110;
    rom[53733] = 25'b1111111111001001100101111;
    rom[53734] = 25'b1111111111001001101001000;
    rom[53735] = 25'b1111111111001001101100001;
    rom[53736] = 25'b1111111111001001101111001;
    rom[53737] = 25'b1111111111001001110010011;
    rom[53738] = 25'b1111111111001001110101011;
    rom[53739] = 25'b1111111111001001111000100;
    rom[53740] = 25'b1111111111001001111011101;
    rom[53741] = 25'b1111111111001001111110110;
    rom[53742] = 25'b1111111111001010000001111;
    rom[53743] = 25'b1111111111001010000101000;
    rom[53744] = 25'b1111111111001010001000001;
    rom[53745] = 25'b1111111111001010001011010;
    rom[53746] = 25'b1111111111001010001110100;
    rom[53747] = 25'b1111111111001010010001101;
    rom[53748] = 25'b1111111111001010010100110;
    rom[53749] = 25'b1111111111001010010111111;
    rom[53750] = 25'b1111111111001010011011000;
    rom[53751] = 25'b1111111111001010011110010;
    rom[53752] = 25'b1111111111001010100001010;
    rom[53753] = 25'b1111111111001010100100100;
    rom[53754] = 25'b1111111111001010100111101;
    rom[53755] = 25'b1111111111001010101010111;
    rom[53756] = 25'b1111111111001010101110000;
    rom[53757] = 25'b1111111111001010110001001;
    rom[53758] = 25'b1111111111001010110100011;
    rom[53759] = 25'b1111111111001010110111100;
    rom[53760] = 25'b1111111111001010111010110;
    rom[53761] = 25'b1111111111001010111101111;
    rom[53762] = 25'b1111111111001011000001000;
    rom[53763] = 25'b1111111111001011000100010;
    rom[53764] = 25'b1111111111001011000111011;
    rom[53765] = 25'b1111111111001011001010101;
    rom[53766] = 25'b1111111111001011001101111;
    rom[53767] = 25'b1111111111001011010001000;
    rom[53768] = 25'b1111111111001011010100010;
    rom[53769] = 25'b1111111111001011010111100;
    rom[53770] = 25'b1111111111001011011010101;
    rom[53771] = 25'b1111111111001011011101111;
    rom[53772] = 25'b1111111111001011100001001;
    rom[53773] = 25'b1111111111001011100100010;
    rom[53774] = 25'b1111111111001011100111100;
    rom[53775] = 25'b1111111111001011101010110;
    rom[53776] = 25'b1111111111001011101110000;
    rom[53777] = 25'b1111111111001011110001001;
    rom[53778] = 25'b1111111111001011110100011;
    rom[53779] = 25'b1111111111001011110111101;
    rom[53780] = 25'b1111111111001011111010111;
    rom[53781] = 25'b1111111111001011111110001;
    rom[53782] = 25'b1111111111001100000001010;
    rom[53783] = 25'b1111111111001100000100101;
    rom[53784] = 25'b1111111111001100000111111;
    rom[53785] = 25'b1111111111001100001011001;
    rom[53786] = 25'b1111111111001100001110010;
    rom[53787] = 25'b1111111111001100010001100;
    rom[53788] = 25'b1111111111001100010100111;
    rom[53789] = 25'b1111111111001100011000001;
    rom[53790] = 25'b1111111111001100011011011;
    rom[53791] = 25'b1111111111001100011110101;
    rom[53792] = 25'b1111111111001100100001111;
    rom[53793] = 25'b1111111111001100100101001;
    rom[53794] = 25'b1111111111001100101000011;
    rom[53795] = 25'b1111111111001100101011110;
    rom[53796] = 25'b1111111111001100101111000;
    rom[53797] = 25'b1111111111001100110010010;
    rom[53798] = 25'b1111111111001100110101100;
    rom[53799] = 25'b1111111111001100111000111;
    rom[53800] = 25'b1111111111001100111100001;
    rom[53801] = 25'b1111111111001100111111011;
    rom[53802] = 25'b1111111111001101000010101;
    rom[53803] = 25'b1111111111001101000110000;
    rom[53804] = 25'b1111111111001101001001010;
    rom[53805] = 25'b1111111111001101001100101;
    rom[53806] = 25'b1111111111001101001111111;
    rom[53807] = 25'b1111111111001101010011010;
    rom[53808] = 25'b1111111111001101010110100;
    rom[53809] = 25'b1111111111001101011001111;
    rom[53810] = 25'b1111111111001101011101001;
    rom[53811] = 25'b1111111111001101100000100;
    rom[53812] = 25'b1111111111001101100011110;
    rom[53813] = 25'b1111111111001101100111001;
    rom[53814] = 25'b1111111111001101101010011;
    rom[53815] = 25'b1111111111001101101101110;
    rom[53816] = 25'b1111111111001101110001001;
    rom[53817] = 25'b1111111111001101110100011;
    rom[53818] = 25'b1111111111001101110111110;
    rom[53819] = 25'b1111111111001101111011001;
    rom[53820] = 25'b1111111111001101111110011;
    rom[53821] = 25'b1111111111001110000001110;
    rom[53822] = 25'b1111111111001110000101001;
    rom[53823] = 25'b1111111111001110001000011;
    rom[53824] = 25'b1111111111001110001011110;
    rom[53825] = 25'b1111111111001110001111001;
    rom[53826] = 25'b1111111111001110010010011;
    rom[53827] = 25'b1111111111001110010101110;
    rom[53828] = 25'b1111111111001110011001001;
    rom[53829] = 25'b1111111111001110011100100;
    rom[53830] = 25'b1111111111001110011111111;
    rom[53831] = 25'b1111111111001110100011010;
    rom[53832] = 25'b1111111111001110100110101;
    rom[53833] = 25'b1111111111001110101010000;
    rom[53834] = 25'b1111111111001110101101011;
    rom[53835] = 25'b1111111111001110110000110;
    rom[53836] = 25'b1111111111001110110100001;
    rom[53837] = 25'b1111111111001110110111100;
    rom[53838] = 25'b1111111111001110111010111;
    rom[53839] = 25'b1111111111001110111110010;
    rom[53840] = 25'b1111111111001111000001101;
    rom[53841] = 25'b1111111111001111000101000;
    rom[53842] = 25'b1111111111001111001000011;
    rom[53843] = 25'b1111111111001111001011111;
    rom[53844] = 25'b1111111111001111001111010;
    rom[53845] = 25'b1111111111001111010010101;
    rom[53846] = 25'b1111111111001111010110000;
    rom[53847] = 25'b1111111111001111011001011;
    rom[53848] = 25'b1111111111001111011100110;
    rom[53849] = 25'b1111111111001111100000010;
    rom[53850] = 25'b1111111111001111100011101;
    rom[53851] = 25'b1111111111001111100111000;
    rom[53852] = 25'b1111111111001111101010100;
    rom[53853] = 25'b1111111111001111101101111;
    rom[53854] = 25'b1111111111001111110001010;
    rom[53855] = 25'b1111111111001111110100101;
    rom[53856] = 25'b1111111111001111111000001;
    rom[53857] = 25'b1111111111001111111011101;
    rom[53858] = 25'b1111111111001111111111000;
    rom[53859] = 25'b1111111111010000000010011;
    rom[53860] = 25'b1111111111010000000101111;
    rom[53861] = 25'b1111111111010000001001010;
    rom[53862] = 25'b1111111111010000001100101;
    rom[53863] = 25'b1111111111010000010000001;
    rom[53864] = 25'b1111111111010000010011101;
    rom[53865] = 25'b1111111111010000010111000;
    rom[53866] = 25'b1111111111010000011010100;
    rom[53867] = 25'b1111111111010000011101111;
    rom[53868] = 25'b1111111111010000100001010;
    rom[53869] = 25'b1111111111010000100100110;
    rom[53870] = 25'b1111111111010000101000010;
    rom[53871] = 25'b1111111111010000101011101;
    rom[53872] = 25'b1111111111010000101111001;
    rom[53873] = 25'b1111111111010000110010101;
    rom[53874] = 25'b1111111111010000110110000;
    rom[53875] = 25'b1111111111010000111001100;
    rom[53876] = 25'b1111111111010000111101000;
    rom[53877] = 25'b1111111111010001000000100;
    rom[53878] = 25'b1111111111010001000100000;
    rom[53879] = 25'b1111111111010001000111011;
    rom[53880] = 25'b1111111111010001001010111;
    rom[53881] = 25'b1111111111010001001110011;
    rom[53882] = 25'b1111111111010001010001111;
    rom[53883] = 25'b1111111111010001010101011;
    rom[53884] = 25'b1111111111010001011000110;
    rom[53885] = 25'b1111111111010001011100010;
    rom[53886] = 25'b1111111111010001011111110;
    rom[53887] = 25'b1111111111010001100011010;
    rom[53888] = 25'b1111111111010001100110110;
    rom[53889] = 25'b1111111111010001101010010;
    rom[53890] = 25'b1111111111010001101101110;
    rom[53891] = 25'b1111111111010001110001010;
    rom[53892] = 25'b1111111111010001110100110;
    rom[53893] = 25'b1111111111010001111000010;
    rom[53894] = 25'b1111111111010001111011110;
    rom[53895] = 25'b1111111111010001111111010;
    rom[53896] = 25'b1111111111010010000010110;
    rom[53897] = 25'b1111111111010010000110010;
    rom[53898] = 25'b1111111111010010001001110;
    rom[53899] = 25'b1111111111010010001101010;
    rom[53900] = 25'b1111111111010010010000110;
    rom[53901] = 25'b1111111111010010010100010;
    rom[53902] = 25'b1111111111010010010111111;
    rom[53903] = 25'b1111111111010010011011010;
    rom[53904] = 25'b1111111111010010011110111;
    rom[53905] = 25'b1111111111010010100010011;
    rom[53906] = 25'b1111111111010010100101111;
    rom[53907] = 25'b1111111111010010101001011;
    rom[53908] = 25'b1111111111010010101100111;
    rom[53909] = 25'b1111111111010010110000100;
    rom[53910] = 25'b1111111111010010110100000;
    rom[53911] = 25'b1111111111010010110111101;
    rom[53912] = 25'b1111111111010010111011000;
    rom[53913] = 25'b1111111111010010111110101;
    rom[53914] = 25'b1111111111010011000010001;
    rom[53915] = 25'b1111111111010011000101101;
    rom[53916] = 25'b1111111111010011001001010;
    rom[53917] = 25'b1111111111010011001100110;
    rom[53918] = 25'b1111111111010011010000011;
    rom[53919] = 25'b1111111111010011010011111;
    rom[53920] = 25'b1111111111010011010111011;
    rom[53921] = 25'b1111111111010011011011000;
    rom[53922] = 25'b1111111111010011011110100;
    rom[53923] = 25'b1111111111010011100010000;
    rom[53924] = 25'b1111111111010011100101101;
    rom[53925] = 25'b1111111111010011101001001;
    rom[53926] = 25'b1111111111010011101100110;
    rom[53927] = 25'b1111111111010011110000011;
    rom[53928] = 25'b1111111111010011110011111;
    rom[53929] = 25'b1111111111010011110111100;
    rom[53930] = 25'b1111111111010011111011000;
    rom[53931] = 25'b1111111111010011111110100;
    rom[53932] = 25'b1111111111010100000010001;
    rom[53933] = 25'b1111111111010100000101110;
    rom[53934] = 25'b1111111111010100001001010;
    rom[53935] = 25'b1111111111010100001100111;
    rom[53936] = 25'b1111111111010100010000100;
    rom[53937] = 25'b1111111111010100010100000;
    rom[53938] = 25'b1111111111010100010111101;
    rom[53939] = 25'b1111111111010100011011010;
    rom[53940] = 25'b1111111111010100011110110;
    rom[53941] = 25'b1111111111010100100010011;
    rom[53942] = 25'b1111111111010100100110000;
    rom[53943] = 25'b1111111111010100101001101;
    rom[53944] = 25'b1111111111010100101101001;
    rom[53945] = 25'b1111111111010100110000110;
    rom[53946] = 25'b1111111111010100110100011;
    rom[53947] = 25'b1111111111010100111000000;
    rom[53948] = 25'b1111111111010100111011100;
    rom[53949] = 25'b1111111111010100111111001;
    rom[53950] = 25'b1111111111010101000010110;
    rom[53951] = 25'b1111111111010101000110011;
    rom[53952] = 25'b1111111111010101001001111;
    rom[53953] = 25'b1111111111010101001101100;
    rom[53954] = 25'b1111111111010101010001010;
    rom[53955] = 25'b1111111111010101010100110;
    rom[53956] = 25'b1111111111010101011000011;
    rom[53957] = 25'b1111111111010101011100000;
    rom[53958] = 25'b1111111111010101011111101;
    rom[53959] = 25'b1111111111010101100011010;
    rom[53960] = 25'b1111111111010101100110111;
    rom[53961] = 25'b1111111111010101101010100;
    rom[53962] = 25'b1111111111010101101110000;
    rom[53963] = 25'b1111111111010101110001110;
    rom[53964] = 25'b1111111111010101110101011;
    rom[53965] = 25'b1111111111010101111001000;
    rom[53966] = 25'b1111111111010101111100101;
    rom[53967] = 25'b1111111111010110000000010;
    rom[53968] = 25'b1111111111010110000011110;
    rom[53969] = 25'b1111111111010110000111100;
    rom[53970] = 25'b1111111111010110001011001;
    rom[53971] = 25'b1111111111010110001110110;
    rom[53972] = 25'b1111111111010110010010011;
    rom[53973] = 25'b1111111111010110010110000;
    rom[53974] = 25'b1111111111010110011001101;
    rom[53975] = 25'b1111111111010110011101010;
    rom[53976] = 25'b1111111111010110100001000;
    rom[53977] = 25'b1111111111010110100100101;
    rom[53978] = 25'b1111111111010110101000010;
    rom[53979] = 25'b1111111111010110101011111;
    rom[53980] = 25'b1111111111010110101111100;
    rom[53981] = 25'b1111111111010110110011001;
    rom[53982] = 25'b1111111111010110110110110;
    rom[53983] = 25'b1111111111010110111010100;
    rom[53984] = 25'b1111111111010110111110001;
    rom[53985] = 25'b1111111111010111000001111;
    rom[53986] = 25'b1111111111010111000101100;
    rom[53987] = 25'b1111111111010111001001001;
    rom[53988] = 25'b1111111111010111001100110;
    rom[53989] = 25'b1111111111010111010000011;
    rom[53990] = 25'b1111111111010111010100001;
    rom[53991] = 25'b1111111111010111010111110;
    rom[53992] = 25'b1111111111010111011011011;
    rom[53993] = 25'b1111111111010111011111000;
    rom[53994] = 25'b1111111111010111100010110;
    rom[53995] = 25'b1111111111010111100110011;
    rom[53996] = 25'b1111111111010111101010001;
    rom[53997] = 25'b1111111111010111101101110;
    rom[53998] = 25'b1111111111010111110001100;
    rom[53999] = 25'b1111111111010111110101001;
    rom[54000] = 25'b1111111111010111111000110;
    rom[54001] = 25'b1111111111010111111100100;
    rom[54002] = 25'b1111111111011000000000001;
    rom[54003] = 25'b1111111111011000000011111;
    rom[54004] = 25'b1111111111011000000111100;
    rom[54005] = 25'b1111111111011000001011001;
    rom[54006] = 25'b1111111111011000001110111;
    rom[54007] = 25'b1111111111011000010010100;
    rom[54008] = 25'b1111111111011000010110010;
    rom[54009] = 25'b1111111111011000011001111;
    rom[54010] = 25'b1111111111011000011101101;
    rom[54011] = 25'b1111111111011000100001010;
    rom[54012] = 25'b1111111111011000100101000;
    rom[54013] = 25'b1111111111011000101000101;
    rom[54014] = 25'b1111111111011000101100011;
    rom[54015] = 25'b1111111111011000110000000;
    rom[54016] = 25'b1111111111011000110011110;
    rom[54017] = 25'b1111111111011000110111100;
    rom[54018] = 25'b1111111111011000111011001;
    rom[54019] = 25'b1111111111011000111110111;
    rom[54020] = 25'b1111111111011001000010100;
    rom[54021] = 25'b1111111111011001000110010;
    rom[54022] = 25'b1111111111011001001010000;
    rom[54023] = 25'b1111111111011001001101101;
    rom[54024] = 25'b1111111111011001010001011;
    rom[54025] = 25'b1111111111011001010101001;
    rom[54026] = 25'b1111111111011001011000111;
    rom[54027] = 25'b1111111111011001011100100;
    rom[54028] = 25'b1111111111011001100000010;
    rom[54029] = 25'b1111111111011001100011111;
    rom[54030] = 25'b1111111111011001100111101;
    rom[54031] = 25'b1111111111011001101011011;
    rom[54032] = 25'b1111111111011001101111000;
    rom[54033] = 25'b1111111111011001110010110;
    rom[54034] = 25'b1111111111011001110110100;
    rom[54035] = 25'b1111111111011001111010001;
    rom[54036] = 25'b1111111111011001111101111;
    rom[54037] = 25'b1111111111011010000001101;
    rom[54038] = 25'b1111111111011010000101011;
    rom[54039] = 25'b1111111111011010001001001;
    rom[54040] = 25'b1111111111011010001100111;
    rom[54041] = 25'b1111111111011010010000100;
    rom[54042] = 25'b1111111111011010010100010;
    rom[54043] = 25'b1111111111011010011000000;
    rom[54044] = 25'b1111111111011010011011110;
    rom[54045] = 25'b1111111111011010011111011;
    rom[54046] = 25'b1111111111011010100011001;
    rom[54047] = 25'b1111111111011010100110111;
    rom[54048] = 25'b1111111111011010101010101;
    rom[54049] = 25'b1111111111011010101110011;
    rom[54050] = 25'b1111111111011010110010001;
    rom[54051] = 25'b1111111111011010110101111;
    rom[54052] = 25'b1111111111011010111001101;
    rom[54053] = 25'b1111111111011010111101010;
    rom[54054] = 25'b1111111111011011000001000;
    rom[54055] = 25'b1111111111011011000100110;
    rom[54056] = 25'b1111111111011011001000100;
    rom[54057] = 25'b1111111111011011001100010;
    rom[54058] = 25'b1111111111011011010000000;
    rom[54059] = 25'b1111111111011011010011110;
    rom[54060] = 25'b1111111111011011010111100;
    rom[54061] = 25'b1111111111011011011011010;
    rom[54062] = 25'b1111111111011011011110111;
    rom[54063] = 25'b1111111111011011100010110;
    rom[54064] = 25'b1111111111011011100110100;
    rom[54065] = 25'b1111111111011011101010010;
    rom[54066] = 25'b1111111111011011101110000;
    rom[54067] = 25'b1111111111011011110001110;
    rom[54068] = 25'b1111111111011011110101011;
    rom[54069] = 25'b1111111111011011111001001;
    rom[54070] = 25'b1111111111011011111101000;
    rom[54071] = 25'b1111111111011100000000110;
    rom[54072] = 25'b1111111111011100000100100;
    rom[54073] = 25'b1111111111011100001000010;
    rom[54074] = 25'b1111111111011100001100000;
    rom[54075] = 25'b1111111111011100001111110;
    rom[54076] = 25'b1111111111011100010011100;
    rom[54077] = 25'b1111111111011100010111010;
    rom[54078] = 25'b1111111111011100011011000;
    rom[54079] = 25'b1111111111011100011110110;
    rom[54080] = 25'b1111111111011100100010100;
    rom[54081] = 25'b1111111111011100100110010;
    rom[54082] = 25'b1111111111011100101010001;
    rom[54083] = 25'b1111111111011100101101111;
    rom[54084] = 25'b1111111111011100110001101;
    rom[54085] = 25'b1111111111011100110101011;
    rom[54086] = 25'b1111111111011100111001001;
    rom[54087] = 25'b1111111111011100111100111;
    rom[54088] = 25'b1111111111011101000000110;
    rom[54089] = 25'b1111111111011101000100100;
    rom[54090] = 25'b1111111111011101001000001;
    rom[54091] = 25'b1111111111011101001100000;
    rom[54092] = 25'b1111111111011101001111110;
    rom[54093] = 25'b1111111111011101010011100;
    rom[54094] = 25'b1111111111011101010111010;
    rom[54095] = 25'b1111111111011101011011000;
    rom[54096] = 25'b1111111111011101011110111;
    rom[54097] = 25'b1111111111011101100010101;
    rom[54098] = 25'b1111111111011101100110011;
    rom[54099] = 25'b1111111111011101101010001;
    rom[54100] = 25'b1111111111011101101101111;
    rom[54101] = 25'b1111111111011101110001110;
    rom[54102] = 25'b1111111111011101110101100;
    rom[54103] = 25'b1111111111011101111001010;
    rom[54104] = 25'b1111111111011101111101000;
    rom[54105] = 25'b1111111111011110000000111;
    rom[54106] = 25'b1111111111011110000100101;
    rom[54107] = 25'b1111111111011110001000011;
    rom[54108] = 25'b1111111111011110001100001;
    rom[54109] = 25'b1111111111011110010000000;
    rom[54110] = 25'b1111111111011110010011110;
    rom[54111] = 25'b1111111111011110010111100;
    rom[54112] = 25'b1111111111011110011011010;
    rom[54113] = 25'b1111111111011110011111001;
    rom[54114] = 25'b1111111111011110100010111;
    rom[54115] = 25'b1111111111011110100110101;
    rom[54116] = 25'b1111111111011110101010011;
    rom[54117] = 25'b1111111111011110101110010;
    rom[54118] = 25'b1111111111011110110010000;
    rom[54119] = 25'b1111111111011110110101110;
    rom[54120] = 25'b1111111111011110111001101;
    rom[54121] = 25'b1111111111011110111101011;
    rom[54122] = 25'b1111111111011111000001010;
    rom[54123] = 25'b1111111111011111000101000;
    rom[54124] = 25'b1111111111011111001000110;
    rom[54125] = 25'b1111111111011111001100101;
    rom[54126] = 25'b1111111111011111010000011;
    rom[54127] = 25'b1111111111011111010100001;
    rom[54128] = 25'b1111111111011111010111111;
    rom[54129] = 25'b1111111111011111011011110;
    rom[54130] = 25'b1111111111011111011111100;
    rom[54131] = 25'b1111111111011111100011010;
    rom[54132] = 25'b1111111111011111100111001;
    rom[54133] = 25'b1111111111011111101011000;
    rom[54134] = 25'b1111111111011111101110101;
    rom[54135] = 25'b1111111111011111110010100;
    rom[54136] = 25'b1111111111011111110110011;
    rom[54137] = 25'b1111111111011111111010001;
    rom[54138] = 25'b1111111111011111111101111;
    rom[54139] = 25'b1111111111100000000001110;
    rom[54140] = 25'b1111111111100000000101100;
    rom[54141] = 25'b1111111111100000001001010;
    rom[54142] = 25'b1111111111100000001101001;
    rom[54143] = 25'b1111111111100000010001000;
    rom[54144] = 25'b1111111111100000010100110;
    rom[54145] = 25'b1111111111100000011000100;
    rom[54146] = 25'b1111111111100000011100011;
    rom[54147] = 25'b1111111111100000100000001;
    rom[54148] = 25'b1111111111100000100011111;
    rom[54149] = 25'b1111111111100000100111110;
    rom[54150] = 25'b1111111111100000101011101;
    rom[54151] = 25'b1111111111100000101111010;
    rom[54152] = 25'b1111111111100000110011001;
    rom[54153] = 25'b1111111111100000110111000;
    rom[54154] = 25'b1111111111100000111010110;
    rom[54155] = 25'b1111111111100000111110100;
    rom[54156] = 25'b1111111111100001000010011;
    rom[54157] = 25'b1111111111100001000110001;
    rom[54158] = 25'b1111111111100001001010000;
    rom[54159] = 25'b1111111111100001001101111;
    rom[54160] = 25'b1111111111100001010001101;
    rom[54161] = 25'b1111111111100001010101011;
    rom[54162] = 25'b1111111111100001011001010;
    rom[54163] = 25'b1111111111100001011101001;
    rom[54164] = 25'b1111111111100001100000111;
    rom[54165] = 25'b1111111111100001100100101;
    rom[54166] = 25'b1111111111100001101000100;
    rom[54167] = 25'b1111111111100001101100010;
    rom[54168] = 25'b1111111111100001110000001;
    rom[54169] = 25'b1111111111100001110100000;
    rom[54170] = 25'b1111111111100001110111101;
    rom[54171] = 25'b1111111111100001111011100;
    rom[54172] = 25'b1111111111100001111111011;
    rom[54173] = 25'b1111111111100010000011001;
    rom[54174] = 25'b1111111111100010000111000;
    rom[54175] = 25'b1111111111100010001010111;
    rom[54176] = 25'b1111111111100010001110100;
    rom[54177] = 25'b1111111111100010010010011;
    rom[54178] = 25'b1111111111100010010110010;
    rom[54179] = 25'b1111111111100010011010000;
    rom[54180] = 25'b1111111111100010011101111;
    rom[54181] = 25'b1111111111100010100001110;
    rom[54182] = 25'b1111111111100010100101100;
    rom[54183] = 25'b1111111111100010101001010;
    rom[54184] = 25'b1111111111100010101101001;
    rom[54185] = 25'b1111111111100010110000111;
    rom[54186] = 25'b1111111111100010110100110;
    rom[54187] = 25'b1111111111100010111000101;
    rom[54188] = 25'b1111111111100010111100011;
    rom[54189] = 25'b1111111111100011000000010;
    rom[54190] = 25'b1111111111100011000100000;
    rom[54191] = 25'b1111111111100011000111110;
    rom[54192] = 25'b1111111111100011001011101;
    rom[54193] = 25'b1111111111100011001111100;
    rom[54194] = 25'b1111111111100011010011010;
    rom[54195] = 25'b1111111111100011010111001;
    rom[54196] = 25'b1111111111100011011011000;
    rom[54197] = 25'b1111111111100011011110110;
    rom[54198] = 25'b1111111111100011100010101;
    rom[54199] = 25'b1111111111100011100110011;
    rom[54200] = 25'b1111111111100011101010001;
    rom[54201] = 25'b1111111111100011101110000;
    rom[54202] = 25'b1111111111100011110001111;
    rom[54203] = 25'b1111111111100011110101101;
    rom[54204] = 25'b1111111111100011111001100;
    rom[54205] = 25'b1111111111100011111101011;
    rom[54206] = 25'b1111111111100100000001001;
    rom[54207] = 25'b1111111111100100000101000;
    rom[54208] = 25'b1111111111100100001000110;
    rom[54209] = 25'b1111111111100100001100100;
    rom[54210] = 25'b1111111111100100010000011;
    rom[54211] = 25'b1111111111100100010100010;
    rom[54212] = 25'b1111111111100100011000000;
    rom[54213] = 25'b1111111111100100011011111;
    rom[54214] = 25'b1111111111100100011111101;
    rom[54215] = 25'b1111111111100100100011100;
    rom[54216] = 25'b1111111111100100100111011;
    rom[54217] = 25'b1111111111100100101011001;
    rom[54218] = 25'b1111111111100100101111000;
    rom[54219] = 25'b1111111111100100110010110;
    rom[54220] = 25'b1111111111100100110110101;
    rom[54221] = 25'b1111111111100100111010011;
    rom[54222] = 25'b1111111111100100111110010;
    rom[54223] = 25'b1111111111100101000010000;
    rom[54224] = 25'b1111111111100101000101111;
    rom[54225] = 25'b1111111111100101001001110;
    rom[54226] = 25'b1111111111100101001101100;
    rom[54227] = 25'b1111111111100101010001011;
    rom[54228] = 25'b1111111111100101010101010;
    rom[54229] = 25'b1111111111100101011001000;
    rom[54230] = 25'b1111111111100101011100110;
    rom[54231] = 25'b1111111111100101100000101;
    rom[54232] = 25'b1111111111100101100100011;
    rom[54233] = 25'b1111111111100101101000010;
    rom[54234] = 25'b1111111111100101101100001;
    rom[54235] = 25'b1111111111100101101111111;
    rom[54236] = 25'b1111111111100101110011110;
    rom[54237] = 25'b1111111111100101110111101;
    rom[54238] = 25'b1111111111100101111011011;
    rom[54239] = 25'b1111111111100101111111010;
    rom[54240] = 25'b1111111111100110000011000;
    rom[54241] = 25'b1111111111100110000110110;
    rom[54242] = 25'b1111111111100110001010101;
    rom[54243] = 25'b1111111111100110001110100;
    rom[54244] = 25'b1111111111100110010010010;
    rom[54245] = 25'b1111111111100110010110001;
    rom[54246] = 25'b1111111111100110011001111;
    rom[54247] = 25'b1111111111100110011101110;
    rom[54248] = 25'b1111111111100110100001101;
    rom[54249] = 25'b1111111111100110100101011;
    rom[54250] = 25'b1111111111100110101001010;
    rom[54251] = 25'b1111111111100110101101000;
    rom[54252] = 25'b1111111111100110110000110;
    rom[54253] = 25'b1111111111100110110100101;
    rom[54254] = 25'b1111111111100110111000100;
    rom[54255] = 25'b1111111111100110111100010;
    rom[54256] = 25'b1111111111100111000000001;
    rom[54257] = 25'b1111111111100111000100000;
    rom[54258] = 25'b1111111111100111000111110;
    rom[54259] = 25'b1111111111100111001011100;
    rom[54260] = 25'b1111111111100111001111011;
    rom[54261] = 25'b1111111111100111010011001;
    rom[54262] = 25'b1111111111100111010111000;
    rom[54263] = 25'b1111111111100111011010111;
    rom[54264] = 25'b1111111111100111011110101;
    rom[54265] = 25'b1111111111100111100010100;
    rom[54266] = 25'b1111111111100111100110011;
    rom[54267] = 25'b1111111111100111101010000;
    rom[54268] = 25'b1111111111100111101101111;
    rom[54269] = 25'b1111111111100111110001110;
    rom[54270] = 25'b1111111111100111110101100;
    rom[54271] = 25'b1111111111100111111001011;
    rom[54272] = 25'b1111111111100111111101010;
    rom[54273] = 25'b1111111111101000000000111;
    rom[54274] = 25'b1111111111101000000100110;
    rom[54275] = 25'b1111111111101000001000101;
    rom[54276] = 25'b1111111111101000001100011;
    rom[54277] = 25'b1111111111101000010000010;
    rom[54278] = 25'b1111111111101000010100001;
    rom[54279] = 25'b1111111111101000010111111;
    rom[54280] = 25'b1111111111101000011011101;
    rom[54281] = 25'b1111111111101000011111100;
    rom[54282] = 25'b1111111111101000100011010;
    rom[54283] = 25'b1111111111101000100111001;
    rom[54284] = 25'b1111111111101000101011000;
    rom[54285] = 25'b1111111111101000101110110;
    rom[54286] = 25'b1111111111101000110010100;
    rom[54287] = 25'b1111111111101000110110011;
    rom[54288] = 25'b1111111111101000111010001;
    rom[54289] = 25'b1111111111101000111110000;
    rom[54290] = 25'b1111111111101001000001110;
    rom[54291] = 25'b1111111111101001000101101;
    rom[54292] = 25'b1111111111101001001001011;
    rom[54293] = 25'b1111111111101001001101010;
    rom[54294] = 25'b1111111111101001010001000;
    rom[54295] = 25'b1111111111101001010100110;
    rom[54296] = 25'b1111111111101001011000101;
    rom[54297] = 25'b1111111111101001011100100;
    rom[54298] = 25'b1111111111101001100000010;
    rom[54299] = 25'b1111111111101001100100000;
    rom[54300] = 25'b1111111111101001100111111;
    rom[54301] = 25'b1111111111101001101011101;
    rom[54302] = 25'b1111111111101001101111011;
    rom[54303] = 25'b1111111111101001110011010;
    rom[54304] = 25'b1111111111101001110111001;
    rom[54305] = 25'b1111111111101001111010111;
    rom[54306] = 25'b1111111111101001111110101;
    rom[54307] = 25'b1111111111101010000010100;
    rom[54308] = 25'b1111111111101010000110010;
    rom[54309] = 25'b1111111111101010001010000;
    rom[54310] = 25'b1111111111101010001101111;
    rom[54311] = 25'b1111111111101010010001101;
    rom[54312] = 25'b1111111111101010010101011;
    rom[54313] = 25'b1111111111101010011001010;
    rom[54314] = 25'b1111111111101010011101001;
    rom[54315] = 25'b1111111111101010100000111;
    rom[54316] = 25'b1111111111101010100100101;
    rom[54317] = 25'b1111111111101010101000100;
    rom[54318] = 25'b1111111111101010101100010;
    rom[54319] = 25'b1111111111101010110000000;
    rom[54320] = 25'b1111111111101010110011111;
    rom[54321] = 25'b1111111111101010110111101;
    rom[54322] = 25'b1111111111101010111011011;
    rom[54323] = 25'b1111111111101010111111010;
    rom[54324] = 25'b1111111111101011000011000;
    rom[54325] = 25'b1111111111101011000110111;
    rom[54326] = 25'b1111111111101011001010101;
    rom[54327] = 25'b1111111111101011001110011;
    rom[54328] = 25'b1111111111101011010010010;
    rom[54329] = 25'b1111111111101011010110000;
    rom[54330] = 25'b1111111111101011011001110;
    rom[54331] = 25'b1111111111101011011101101;
    rom[54332] = 25'b1111111111101011100001011;
    rom[54333] = 25'b1111111111101011100101001;
    rom[54334] = 25'b1111111111101011101000111;
    rom[54335] = 25'b1111111111101011101100110;
    rom[54336] = 25'b1111111111101011110000100;
    rom[54337] = 25'b1111111111101011110100010;
    rom[54338] = 25'b1111111111101011111000000;
    rom[54339] = 25'b1111111111101011111011111;
    rom[54340] = 25'b1111111111101011111111110;
    rom[54341] = 25'b1111111111101100000011011;
    rom[54342] = 25'b1111111111101100000111010;
    rom[54343] = 25'b1111111111101100001011000;
    rom[54344] = 25'b1111111111101100001110111;
    rom[54345] = 25'b1111111111101100010010100;
    rom[54346] = 25'b1111111111101100010110011;
    rom[54347] = 25'b1111111111101100011010001;
    rom[54348] = 25'b1111111111101100011101111;
    rom[54349] = 25'b1111111111101100100001110;
    rom[54350] = 25'b1111111111101100100101011;
    rom[54351] = 25'b1111111111101100101001010;
    rom[54352] = 25'b1111111111101100101101000;
    rom[54353] = 25'b1111111111101100110000111;
    rom[54354] = 25'b1111111111101100110100100;
    rom[54355] = 25'b1111111111101100111000011;
    rom[54356] = 25'b1111111111101100111100001;
    rom[54357] = 25'b1111111111101100111111111;
    rom[54358] = 25'b1111111111101101000011101;
    rom[54359] = 25'b1111111111101101000111011;
    rom[54360] = 25'b1111111111101101001011010;
    rom[54361] = 25'b1111111111101101001111000;
    rom[54362] = 25'b1111111111101101010010110;
    rom[54363] = 25'b1111111111101101010110100;
    rom[54364] = 25'b1111111111101101011010010;
    rom[54365] = 25'b1111111111101101011110000;
    rom[54366] = 25'b1111111111101101100001111;
    rom[54367] = 25'b1111111111101101100101101;
    rom[54368] = 25'b1111111111101101101001011;
    rom[54369] = 25'b1111111111101101101101001;
    rom[54370] = 25'b1111111111101101110000111;
    rom[54371] = 25'b1111111111101101110100101;
    rom[54372] = 25'b1111111111101101111000100;
    rom[54373] = 25'b1111111111101101111100001;
    rom[54374] = 25'b1111111111101101111111111;
    rom[54375] = 25'b1111111111101110000011101;
    rom[54376] = 25'b1111111111101110000111100;
    rom[54377] = 25'b1111111111101110001011010;
    rom[54378] = 25'b1111111111101110001111000;
    rom[54379] = 25'b1111111111101110010010101;
    rom[54380] = 25'b1111111111101110010110100;
    rom[54381] = 25'b1111111111101110011010010;
    rom[54382] = 25'b1111111111101110011110000;
    rom[54383] = 25'b1111111111101110100001110;
    rom[54384] = 25'b1111111111101110100101100;
    rom[54385] = 25'b1111111111101110101001010;
    rom[54386] = 25'b1111111111101110101101000;
    rom[54387] = 25'b1111111111101110110000110;
    rom[54388] = 25'b1111111111101110110100100;
    rom[54389] = 25'b1111111111101110111000010;
    rom[54390] = 25'b1111111111101110111100000;
    rom[54391] = 25'b1111111111101110111111110;
    rom[54392] = 25'b1111111111101111000011011;
    rom[54393] = 25'b1111111111101111000111010;
    rom[54394] = 25'b1111111111101111001011000;
    rom[54395] = 25'b1111111111101111001110110;
    rom[54396] = 25'b1111111111101111010010100;
    rom[54397] = 25'b1111111111101111010110010;
    rom[54398] = 25'b1111111111101111011010000;
    rom[54399] = 25'b1111111111101111011101101;
    rom[54400] = 25'b1111111111101111100001011;
    rom[54401] = 25'b1111111111101111100101001;
    rom[54402] = 25'b1111111111101111101000111;
    rom[54403] = 25'b1111111111101111101100101;
    rom[54404] = 25'b1111111111101111110000011;
    rom[54405] = 25'b1111111111101111110100001;
    rom[54406] = 25'b1111111111101111110111111;
    rom[54407] = 25'b1111111111101111111011100;
    rom[54408] = 25'b1111111111101111111111010;
    rom[54409] = 25'b1111111111110000000011000;
    rom[54410] = 25'b1111111111110000000110110;
    rom[54411] = 25'b1111111111110000001010100;
    rom[54412] = 25'b1111111111110000001110010;
    rom[54413] = 25'b1111111111110000010010000;
    rom[54414] = 25'b1111111111110000010101101;
    rom[54415] = 25'b1111111111110000011001011;
    rom[54416] = 25'b1111111111110000011101001;
    rom[54417] = 25'b1111111111110000100000111;
    rom[54418] = 25'b1111111111110000100100100;
    rom[54419] = 25'b1111111111110000101000010;
    rom[54420] = 25'b1111111111110000101100000;
    rom[54421] = 25'b1111111111110000101111101;
    rom[54422] = 25'b1111111111110000110011011;
    rom[54423] = 25'b1111111111110000110111001;
    rom[54424] = 25'b1111111111110000111010111;
    rom[54425] = 25'b1111111111110000111110101;
    rom[54426] = 25'b1111111111110001000010010;
    rom[54427] = 25'b1111111111110001000110000;
    rom[54428] = 25'b1111111111110001001001110;
    rom[54429] = 25'b1111111111110001001101100;
    rom[54430] = 25'b1111111111110001010001001;
    rom[54431] = 25'b1111111111110001010100111;
    rom[54432] = 25'b1111111111110001011000101;
    rom[54433] = 25'b1111111111110001011100010;
    rom[54434] = 25'b1111111111110001100000000;
    rom[54435] = 25'b1111111111110001100011101;
    rom[54436] = 25'b1111111111110001100111011;
    rom[54437] = 25'b1111111111110001101011001;
    rom[54438] = 25'b1111111111110001101110110;
    rom[54439] = 25'b1111111111110001110010100;
    rom[54440] = 25'b1111111111110001110110001;
    rom[54441] = 25'b1111111111110001111001111;
    rom[54442] = 25'b1111111111110001111101100;
    rom[54443] = 25'b1111111111110010000001010;
    rom[54444] = 25'b1111111111110010000100111;
    rom[54445] = 25'b1111111111110010001000101;
    rom[54446] = 25'b1111111111110010001100010;
    rom[54447] = 25'b1111111111110010010000000;
    rom[54448] = 25'b1111111111110010010011101;
    rom[54449] = 25'b1111111111110010010111011;
    rom[54450] = 25'b1111111111110010011011001;
    rom[54451] = 25'b1111111111110010011110110;
    rom[54452] = 25'b1111111111110010100010100;
    rom[54453] = 25'b1111111111110010100110001;
    rom[54454] = 25'b1111111111110010101001111;
    rom[54455] = 25'b1111111111110010101101100;
    rom[54456] = 25'b1111111111110010110001010;
    rom[54457] = 25'b1111111111110010110100111;
    rom[54458] = 25'b1111111111110010111000101;
    rom[54459] = 25'b1111111111110010111100010;
    rom[54460] = 25'b1111111111110010111111111;
    rom[54461] = 25'b1111111111110011000011101;
    rom[54462] = 25'b1111111111110011000111010;
    rom[54463] = 25'b1111111111110011001010111;
    rom[54464] = 25'b1111111111110011001110101;
    rom[54465] = 25'b1111111111110011010010010;
    rom[54466] = 25'b1111111111110011010101111;
    rom[54467] = 25'b1111111111110011011001101;
    rom[54468] = 25'b1111111111110011011101010;
    rom[54469] = 25'b1111111111110011100000111;
    rom[54470] = 25'b1111111111110011100100100;
    rom[54471] = 25'b1111111111110011101000010;
    rom[54472] = 25'b1111111111110011101100000;
    rom[54473] = 25'b1111111111110011101111101;
    rom[54474] = 25'b1111111111110011110011010;
    rom[54475] = 25'b1111111111110011110110111;
    rom[54476] = 25'b1111111111110011111010100;
    rom[54477] = 25'b1111111111110011111110010;
    rom[54478] = 25'b1111111111110100000001111;
    rom[54479] = 25'b1111111111110100000101100;
    rom[54480] = 25'b1111111111110100001001001;
    rom[54481] = 25'b1111111111110100001100110;
    rom[54482] = 25'b1111111111110100010000100;
    rom[54483] = 25'b1111111111110100010100001;
    rom[54484] = 25'b1111111111110100010111110;
    rom[54485] = 25'b1111111111110100011011011;
    rom[54486] = 25'b1111111111110100011111000;
    rom[54487] = 25'b1111111111110100100010101;
    rom[54488] = 25'b1111111111110100100110010;
    rom[54489] = 25'b1111111111110100101010000;
    rom[54490] = 25'b1111111111110100101101101;
    rom[54491] = 25'b1111111111110100110001010;
    rom[54492] = 25'b1111111111110100110100111;
    rom[54493] = 25'b1111111111110100111000100;
    rom[54494] = 25'b1111111111110100111100001;
    rom[54495] = 25'b1111111111110100111111110;
    rom[54496] = 25'b1111111111110101000011011;
    rom[54497] = 25'b1111111111110101000111000;
    rom[54498] = 25'b1111111111110101001010101;
    rom[54499] = 25'b1111111111110101001110010;
    rom[54500] = 25'b1111111111110101010001111;
    rom[54501] = 25'b1111111111110101010101100;
    rom[54502] = 25'b1111111111110101011001001;
    rom[54503] = 25'b1111111111110101011100110;
    rom[54504] = 25'b1111111111110101100000011;
    rom[54505] = 25'b1111111111110101100100000;
    rom[54506] = 25'b1111111111110101100111101;
    rom[54507] = 25'b1111111111110101101011010;
    rom[54508] = 25'b1111111111110101101110111;
    rom[54509] = 25'b1111111111110101110010011;
    rom[54510] = 25'b1111111111110101110110000;
    rom[54511] = 25'b1111111111110101111001110;
    rom[54512] = 25'b1111111111110101111101010;
    rom[54513] = 25'b1111111111110110000000111;
    rom[54514] = 25'b1111111111110110000100100;
    rom[54515] = 25'b1111111111110110001000001;
    rom[54516] = 25'b1111111111110110001011110;
    rom[54517] = 25'b1111111111110110001111010;
    rom[54518] = 25'b1111111111110110010010111;
    rom[54519] = 25'b1111111111110110010110100;
    rom[54520] = 25'b1111111111110110011010001;
    rom[54521] = 25'b1111111111110110011101101;
    rom[54522] = 25'b1111111111110110100001010;
    rom[54523] = 25'b1111111111110110100100111;
    rom[54524] = 25'b1111111111110110101000100;
    rom[54525] = 25'b1111111111110110101100000;
    rom[54526] = 25'b1111111111110110101111101;
    rom[54527] = 25'b1111111111110110110011010;
    rom[54528] = 25'b1111111111110110110110110;
    rom[54529] = 25'b1111111111110110111010011;
    rom[54530] = 25'b1111111111110110111110000;
    rom[54531] = 25'b1111111111110111000001100;
    rom[54532] = 25'b1111111111110111000101001;
    rom[54533] = 25'b1111111111110111001000110;
    rom[54534] = 25'b1111111111110111001100010;
    rom[54535] = 25'b1111111111110111001111111;
    rom[54536] = 25'b1111111111110111010011100;
    rom[54537] = 25'b1111111111110111010111000;
    rom[54538] = 25'b1111111111110111011010100;
    rom[54539] = 25'b1111111111110111011110001;
    rom[54540] = 25'b1111111111110111100001110;
    rom[54541] = 25'b1111111111110111100101010;
    rom[54542] = 25'b1111111111110111101000111;
    rom[54543] = 25'b1111111111110111101100011;
    rom[54544] = 25'b1111111111110111101111111;
    rom[54545] = 25'b1111111111110111110011100;
    rom[54546] = 25'b1111111111110111110111000;
    rom[54547] = 25'b1111111111110111111010101;
    rom[54548] = 25'b1111111111110111111110010;
    rom[54549] = 25'b1111111111111000000001110;
    rom[54550] = 25'b1111111111111000000101011;
    rom[54551] = 25'b1111111111111000001000111;
    rom[54552] = 25'b1111111111111000001100011;
    rom[54553] = 25'b1111111111111000010000000;
    rom[54554] = 25'b1111111111111000010011100;
    rom[54555] = 25'b1111111111111000010111000;
    rom[54556] = 25'b1111111111111000011010100;
    rom[54557] = 25'b1111111111111000011110000;
    rom[54558] = 25'b1111111111111000100001101;
    rom[54559] = 25'b1111111111111000100101001;
    rom[54560] = 25'b1111111111111000101000110;
    rom[54561] = 25'b1111111111111000101100010;
    rom[54562] = 25'b1111111111111000101111110;
    rom[54563] = 25'b1111111111111000110011010;
    rom[54564] = 25'b1111111111111000110110110;
    rom[54565] = 25'b1111111111111000111010011;
    rom[54566] = 25'b1111111111111000111101111;
    rom[54567] = 25'b1111111111111001000001011;
    rom[54568] = 25'b1111111111111001000100111;
    rom[54569] = 25'b1111111111111001001000100;
    rom[54570] = 25'b1111111111111001001011111;
    rom[54571] = 25'b1111111111111001001111100;
    rom[54572] = 25'b1111111111111001010011000;
    rom[54573] = 25'b1111111111111001010110100;
    rom[54574] = 25'b1111111111111001011010000;
    rom[54575] = 25'b1111111111111001011101100;
    rom[54576] = 25'b1111111111111001100001000;
    rom[54577] = 25'b1111111111111001100100101;
    rom[54578] = 25'b1111111111111001101000000;
    rom[54579] = 25'b1111111111111001101011101;
    rom[54580] = 25'b1111111111111001101111000;
    rom[54581] = 25'b1111111111111001110010101;
    rom[54582] = 25'b1111111111111001110110000;
    rom[54583] = 25'b1111111111111001111001100;
    rom[54584] = 25'b1111111111111001111101000;
    rom[54585] = 25'b1111111111111010000000100;
    rom[54586] = 25'b1111111111111010000100000;
    rom[54587] = 25'b1111111111111010000111100;
    rom[54588] = 25'b1111111111111010001011000;
    rom[54589] = 25'b1111111111111010001110100;
    rom[54590] = 25'b1111111111111010010010000;
    rom[54591] = 25'b1111111111111010010101011;
    rom[54592] = 25'b1111111111111010011001000;
    rom[54593] = 25'b1111111111111010011100011;
    rom[54594] = 25'b1111111111111010011111111;
    rom[54595] = 25'b1111111111111010100011011;
    rom[54596] = 25'b1111111111111010100110110;
    rom[54597] = 25'b1111111111111010101010011;
    rom[54598] = 25'b1111111111111010101101110;
    rom[54599] = 25'b1111111111111010110001010;
    rom[54600] = 25'b1111111111111010110100110;
    rom[54601] = 25'b1111111111111010111000001;
    rom[54602] = 25'b1111111111111010111011101;
    rom[54603] = 25'b1111111111111010111111000;
    rom[54604] = 25'b1111111111111011000010100;
    rom[54605] = 25'b1111111111111011000110000;
    rom[54606] = 25'b1111111111111011001001011;
    rom[54607] = 25'b1111111111111011001100111;
    rom[54608] = 25'b1111111111111011010000011;
    rom[54609] = 25'b1111111111111011010011110;
    rom[54610] = 25'b1111111111111011010111010;
    rom[54611] = 25'b1111111111111011011010110;
    rom[54612] = 25'b1111111111111011011110001;
    rom[54613] = 25'b1111111111111011100001101;
    rom[54614] = 25'b1111111111111011100101001;
    rom[54615] = 25'b1111111111111011101000011;
    rom[54616] = 25'b1111111111111011101011111;
    rom[54617] = 25'b1111111111111011101111011;
    rom[54618] = 25'b1111111111111011110010110;
    rom[54619] = 25'b1111111111111011110110010;
    rom[54620] = 25'b1111111111111011111001101;
    rom[54621] = 25'b1111111111111011111101001;
    rom[54622] = 25'b1111111111111100000000100;
    rom[54623] = 25'b1111111111111100000011111;
    rom[54624] = 25'b1111111111111100000111011;
    rom[54625] = 25'b1111111111111100001010110;
    rom[54626] = 25'b1111111111111100001110001;
    rom[54627] = 25'b1111111111111100010001101;
    rom[54628] = 25'b1111111111111100010101000;
    rom[54629] = 25'b1111111111111100011000011;
    rom[54630] = 25'b1111111111111100011011110;
    rom[54631] = 25'b1111111111111100011111010;
    rom[54632] = 25'b1111111111111100100010101;
    rom[54633] = 25'b1111111111111100100110001;
    rom[54634] = 25'b1111111111111100101001011;
    rom[54635] = 25'b1111111111111100101100111;
    rom[54636] = 25'b1111111111111100110000010;
    rom[54637] = 25'b1111111111111100110011110;
    rom[54638] = 25'b1111111111111100110111000;
    rom[54639] = 25'b1111111111111100111010011;
    rom[54640] = 25'b1111111111111100111101111;
    rom[54641] = 25'b1111111111111101000001010;
    rom[54642] = 25'b1111111111111101000100101;
    rom[54643] = 25'b1111111111111101001000000;
    rom[54644] = 25'b1111111111111101001011011;
    rom[54645] = 25'b1111111111111101001110110;
    rom[54646] = 25'b1111111111111101010010001;
    rom[54647] = 25'b1111111111111101010101100;
    rom[54648] = 25'b1111111111111101011000111;
    rom[54649] = 25'b1111111111111101011100011;
    rom[54650] = 25'b1111111111111101011111101;
    rom[54651] = 25'b1111111111111101100011000;
    rom[54652] = 25'b1111111111111101100110011;
    rom[54653] = 25'b1111111111111101101001110;
    rom[54654] = 25'b1111111111111101101101001;
    rom[54655] = 25'b1111111111111101110000100;
    rom[54656] = 25'b1111111111111101110011111;
    rom[54657] = 25'b1111111111111101110111010;
    rom[54658] = 25'b1111111111111101111010101;
    rom[54659] = 25'b1111111111111101111110000;
    rom[54660] = 25'b1111111111111110000001010;
    rom[54661] = 25'b1111111111111110000100101;
    rom[54662] = 25'b1111111111111110000111111;
    rom[54663] = 25'b1111111111111110001011010;
    rom[54664] = 25'b1111111111111110001110101;
    rom[54665] = 25'b1111111111111110010010000;
    rom[54666] = 25'b1111111111111110010101011;
    rom[54667] = 25'b1111111111111110011000101;
    rom[54668] = 25'b1111111111111110011100000;
    rom[54669] = 25'b1111111111111110011111011;
    rom[54670] = 25'b1111111111111110100010101;
    rom[54671] = 25'b1111111111111110100110000;
    rom[54672] = 25'b1111111111111110101001011;
    rom[54673] = 25'b1111111111111110101100101;
    rom[54674] = 25'b1111111111111110110000000;
    rom[54675] = 25'b1111111111111110110011011;
    rom[54676] = 25'b1111111111111110110110101;
    rom[54677] = 25'b1111111111111110111010000;
    rom[54678] = 25'b1111111111111110111101010;
    rom[54679] = 25'b1111111111111111000000101;
    rom[54680] = 25'b1111111111111111000011111;
    rom[54681] = 25'b1111111111111111000111010;
    rom[54682] = 25'b1111111111111111001010100;
    rom[54683] = 25'b1111111111111111001101110;
    rom[54684] = 25'b1111111111111111010001001;
    rom[54685] = 25'b1111111111111111010100011;
    rom[54686] = 25'b1111111111111111010111110;
    rom[54687] = 25'b1111111111111111011011000;
    rom[54688] = 25'b1111111111111111011110011;
    rom[54689] = 25'b1111111111111111100001101;
    rom[54690] = 25'b1111111111111111100100111;
    rom[54691] = 25'b1111111111111111101000010;
    rom[54692] = 25'b1111111111111111101011100;
    rom[54693] = 25'b1111111111111111101110110;
    rom[54694] = 25'b1111111111111111110010000;
    rom[54695] = 25'b1111111111111111110101010;
    rom[54696] = 25'b1111111111111111111000100;
    rom[54697] = 25'b1111111111111111111011111;
    rom[54698] = 25'b1111111111111111111111010;
    rom[54699] = 25'b0000000000000000000010011;
    rom[54700] = 25'b0000000000000000000101101;
    rom[54701] = 25'b0000000000000000001000111;
    rom[54702] = 25'b0000000000000000001100001;
    rom[54703] = 25'b0000000000000000001111100;
    rom[54704] = 25'b0000000000000000010010101;
    rom[54705] = 25'b0000000000000000010101111;
    rom[54706] = 25'b0000000000000000011001001;
    rom[54707] = 25'b0000000000000000011100011;
    rom[54708] = 25'b0000000000000000011111110;
    rom[54709] = 25'b0000000000000000100011000;
    rom[54710] = 25'b0000000000000000100110001;
    rom[54711] = 25'b0000000000000000101001011;
    rom[54712] = 25'b0000000000000000101100101;
    rom[54713] = 25'b0000000000000000110000000;
    rom[54714] = 25'b0000000000000000110011001;
    rom[54715] = 25'b0000000000000000110110011;
    rom[54716] = 25'b0000000000000000111001101;
    rom[54717] = 25'b0000000000000000111100111;
    rom[54718] = 25'b0000000000000001000000001;
    rom[54719] = 25'b0000000000000001000011010;
    rom[54720] = 25'b0000000000000001000110100;
    rom[54721] = 25'b0000000000000001001001110;
    rom[54722] = 25'b0000000000000001001101000;
    rom[54723] = 25'b0000000000000001010000001;
    rom[54724] = 25'b0000000000000001010011011;
    rom[54725] = 25'b0000000000000001010110101;
    rom[54726] = 25'b0000000000000001011001111;
    rom[54727] = 25'b0000000000000001011101000;
    rom[54728] = 25'b0000000000000001100000010;
    rom[54729] = 25'b0000000000000001100011100;
    rom[54730] = 25'b0000000000000001100110101;
    rom[54731] = 25'b0000000000000001101001111;
    rom[54732] = 25'b0000000000000001101101001;
    rom[54733] = 25'b0000000000000001110000010;
    rom[54734] = 25'b0000000000000001110011100;
    rom[54735] = 25'b0000000000000001110110101;
    rom[54736] = 25'b0000000000000001111001110;
    rom[54737] = 25'b0000000000000001111101001;
    rom[54738] = 25'b0000000000000010000000010;
    rom[54739] = 25'b0000000000000010000011011;
    rom[54740] = 25'b0000000000000010000110101;
    rom[54741] = 25'b0000000000000010001001110;
    rom[54742] = 25'b0000000000000010001101000;
    rom[54743] = 25'b0000000000000010010000001;
    rom[54744] = 25'b0000000000000010010011010;
    rom[54745] = 25'b0000000000000010010110100;
    rom[54746] = 25'b0000000000000010011001101;
    rom[54747] = 25'b0000000000000010011100111;
    rom[54748] = 25'b0000000000000010100000000;
    rom[54749] = 25'b0000000000000010100011001;
    rom[54750] = 25'b0000000000000010100110010;
    rom[54751] = 25'b0000000000000010101001011;
    rom[54752] = 25'b0000000000000010101100101;
    rom[54753] = 25'b0000000000000010101111110;
    rom[54754] = 25'b0000000000000010110010111;
    rom[54755] = 25'b0000000000000010110110000;
    rom[54756] = 25'b0000000000000010111001010;
    rom[54757] = 25'b0000000000000010111100010;
    rom[54758] = 25'b0000000000000010111111100;
    rom[54759] = 25'b0000000000000011000010100;
    rom[54760] = 25'b0000000000000011000101110;
    rom[54761] = 25'b0000000000000011001000111;
    rom[54762] = 25'b0000000000000011001100000;
    rom[54763] = 25'b0000000000000011001111001;
    rom[54764] = 25'b0000000000000011010010010;
    rom[54765] = 25'b0000000000000011010101011;
    rom[54766] = 25'b0000000000000011011000100;
    rom[54767] = 25'b0000000000000011011011101;
    rom[54768] = 25'b0000000000000011011110110;
    rom[54769] = 25'b0000000000000011100001111;
    rom[54770] = 25'b0000000000000011100100111;
    rom[54771] = 25'b0000000000000011101000001;
    rom[54772] = 25'b0000000000000011101011001;
    rom[54773] = 25'b0000000000000011101110010;
    rom[54774] = 25'b0000000000000011110001011;
    rom[54775] = 25'b0000000000000011110100100;
    rom[54776] = 25'b0000000000000011110111101;
    rom[54777] = 25'b0000000000000011111010101;
    rom[54778] = 25'b0000000000000011111101110;
    rom[54779] = 25'b0000000000000100000000111;
    rom[54780] = 25'b0000000000000100000011111;
    rom[54781] = 25'b0000000000000100000111000;
    rom[54782] = 25'b0000000000000100001010001;
    rom[54783] = 25'b0000000000000100001101001;
    rom[54784] = 25'b0000000000000100010000010;
    rom[54785] = 25'b0000000000000100010011011;
    rom[54786] = 25'b0000000000000100010110011;
    rom[54787] = 25'b0000000000000100011001100;
    rom[54788] = 25'b0000000000000100011100101;
    rom[54789] = 25'b0000000000000100011111101;
    rom[54790] = 25'b0000000000000100100010101;
    rom[54791] = 25'b0000000000000100100101110;
    rom[54792] = 25'b0000000000000100101000111;
    rom[54793] = 25'b0000000000000100101011111;
    rom[54794] = 25'b0000000000000100101110111;
    rom[54795] = 25'b0000000000000100110010000;
    rom[54796] = 25'b0000000000000100110101000;
    rom[54797] = 25'b0000000000000100111000000;
    rom[54798] = 25'b0000000000000100111011001;
    rom[54799] = 25'b0000000000000100111110001;
    rom[54800] = 25'b0000000000000101000001010;
    rom[54801] = 25'b0000000000000101000100010;
    rom[54802] = 25'b0000000000000101000111010;
    rom[54803] = 25'b0000000000000101001010011;
    rom[54804] = 25'b0000000000000101001101011;
    rom[54805] = 25'b0000000000000101010000011;
    rom[54806] = 25'b0000000000000101010011011;
    rom[54807] = 25'b0000000000000101010110011;
    rom[54808] = 25'b0000000000000101011001011;
    rom[54809] = 25'b0000000000000101011100100;
    rom[54810] = 25'b0000000000000101011111100;
    rom[54811] = 25'b0000000000000101100010011;
    rom[54812] = 25'b0000000000000101100101100;
    rom[54813] = 25'b0000000000000101101000100;
    rom[54814] = 25'b0000000000000101101011100;
    rom[54815] = 25'b0000000000000101101110100;
    rom[54816] = 25'b0000000000000101110001100;
    rom[54817] = 25'b0000000000000101110100100;
    rom[54818] = 25'b0000000000000101110111100;
    rom[54819] = 25'b0000000000000101111010011;
    rom[54820] = 25'b0000000000000101111101011;
    rom[54821] = 25'b0000000000000110000000011;
    rom[54822] = 25'b0000000000000110000011011;
    rom[54823] = 25'b0000000000000110000110011;
    rom[54824] = 25'b0000000000000110001001011;
    rom[54825] = 25'b0000000000000110001100011;
    rom[54826] = 25'b0000000000000110001111011;
    rom[54827] = 25'b0000000000000110010010011;
    rom[54828] = 25'b0000000000000110010101011;
    rom[54829] = 25'b0000000000000110011000010;
    rom[54830] = 25'b0000000000000110011011010;
    rom[54831] = 25'b0000000000000110011110010;
    rom[54832] = 25'b0000000000000110100001001;
    rom[54833] = 25'b0000000000000110100100001;
    rom[54834] = 25'b0000000000000110100111001;
    rom[54835] = 25'b0000000000000110101010000;
    rom[54836] = 25'b0000000000000110101101000;
    rom[54837] = 25'b0000000000000110110000000;
    rom[54838] = 25'b0000000000000110110010111;
    rom[54839] = 25'b0000000000000110110101111;
    rom[54840] = 25'b0000000000000110111000110;
    rom[54841] = 25'b0000000000000110111011101;
    rom[54842] = 25'b0000000000000110111110101;
    rom[54843] = 25'b0000000000000111000001100;
    rom[54844] = 25'b0000000000000111000100100;
    rom[54845] = 25'b0000000000000111000111011;
    rom[54846] = 25'b0000000000000111001010010;
    rom[54847] = 25'b0000000000000111001101010;
    rom[54848] = 25'b0000000000000111010000001;
    rom[54849] = 25'b0000000000000111010011000;
    rom[54850] = 25'b0000000000000111010110000;
    rom[54851] = 25'b0000000000000111011000111;
    rom[54852] = 25'b0000000000000111011011111;
    rom[54853] = 25'b0000000000000111011110110;
    rom[54854] = 25'b0000000000000111100001101;
    rom[54855] = 25'b0000000000000111100100100;
    rom[54856] = 25'b0000000000000111100111011;
    rom[54857] = 25'b0000000000000111101010011;
    rom[54858] = 25'b0000000000000111101101010;
    rom[54859] = 25'b0000000000000111110000001;
    rom[54860] = 25'b0000000000000111110011000;
    rom[54861] = 25'b0000000000000111110101111;
    rom[54862] = 25'b0000000000000111111000110;
    rom[54863] = 25'b0000000000000111111011101;
    rom[54864] = 25'b0000000000000111111110100;
    rom[54865] = 25'b0000000000001000000001011;
    rom[54866] = 25'b0000000000001000000100010;
    rom[54867] = 25'b0000000000001000000111001;
    rom[54868] = 25'b0000000000001000001010000;
    rom[54869] = 25'b0000000000001000001100111;
    rom[54870] = 25'b0000000000001000001111101;
    rom[54871] = 25'b0000000000001000010010101;
    rom[54872] = 25'b0000000000001000010101100;
    rom[54873] = 25'b0000000000001000011000010;
    rom[54874] = 25'b0000000000001000011011001;
    rom[54875] = 25'b0000000000001000011110000;
    rom[54876] = 25'b0000000000001000100000111;
    rom[54877] = 25'b0000000000001000100011101;
    rom[54878] = 25'b0000000000001000100110100;
    rom[54879] = 25'b0000000000001000101001011;
    rom[54880] = 25'b0000000000001000101100001;
    rom[54881] = 25'b0000000000001000101111000;
    rom[54882] = 25'b0000000000001000110001111;
    rom[54883] = 25'b0000000000001000110100101;
    rom[54884] = 25'b0000000000001000110111100;
    rom[54885] = 25'b0000000000001000111010011;
    rom[54886] = 25'b0000000000001000111101001;
    rom[54887] = 25'b0000000000001001000000000;
    rom[54888] = 25'b0000000000001001000010110;
    rom[54889] = 25'b0000000000001001000101100;
    rom[54890] = 25'b0000000000001001001000011;
    rom[54891] = 25'b0000000000001001001011001;
    rom[54892] = 25'b0000000000001001001110000;
    rom[54893] = 25'b0000000000001001010000110;
    rom[54894] = 25'b0000000000001001010011100;
    rom[54895] = 25'b0000000000001001010110011;
    rom[54896] = 25'b0000000000001001011001001;
    rom[54897] = 25'b0000000000001001011100000;
    rom[54898] = 25'b0000000000001001011110110;
    rom[54899] = 25'b0000000000001001100001101;
    rom[54900] = 25'b0000000000001001100100010;
    rom[54901] = 25'b0000000000001001100111001;
    rom[54902] = 25'b0000000000001001101001111;
    rom[54903] = 25'b0000000000001001101100101;
    rom[54904] = 25'b0000000000001001101111011;
    rom[54905] = 25'b0000000000001001110010010;
    rom[54906] = 25'b0000000000001001110100111;
    rom[54907] = 25'b0000000000001001110111110;
    rom[54908] = 25'b0000000000001001111010011;
    rom[54909] = 25'b0000000000001001111101010;
    rom[54910] = 25'b0000000000001001111111111;
    rom[54911] = 25'b0000000000001010000010110;
    rom[54912] = 25'b0000000000001010000101011;
    rom[54913] = 25'b0000000000001010001000010;
    rom[54914] = 25'b0000000000001010001011000;
    rom[54915] = 25'b0000000000001010001101110;
    rom[54916] = 25'b0000000000001010010000100;
    rom[54917] = 25'b0000000000001010010011001;
    rom[54918] = 25'b0000000000001010010101111;
    rom[54919] = 25'b0000000000001010011000101;
    rom[54920] = 25'b0000000000001010011011011;
    rom[54921] = 25'b0000000000001010011110001;
    rom[54922] = 25'b0000000000001010100000110;
    rom[54923] = 25'b0000000000001010100011100;
    rom[54924] = 25'b0000000000001010100110010;
    rom[54925] = 25'b0000000000001010101000111;
    rom[54926] = 25'b0000000000001010101011101;
    rom[54927] = 25'b0000000000001010101110011;
    rom[54928] = 25'b0000000000001010110001000;
    rom[54929] = 25'b0000000000001010110011110;
    rom[54930] = 25'b0000000000001010110110100;
    rom[54931] = 25'b0000000000001010111001001;
    rom[54932] = 25'b0000000000001010111011111;
    rom[54933] = 25'b0000000000001010111110101;
    rom[54934] = 25'b0000000000001011000001010;
    rom[54935] = 25'b0000000000001011000011111;
    rom[54936] = 25'b0000000000001011000110101;
    rom[54937] = 25'b0000000000001011001001011;
    rom[54938] = 25'b0000000000001011001011111;
    rom[54939] = 25'b0000000000001011001110101;
    rom[54940] = 25'b0000000000001011010001010;
    rom[54941] = 25'b0000000000001011010100000;
    rom[54942] = 25'b0000000000001011010110101;
    rom[54943] = 25'b0000000000001011011001010;
    rom[54944] = 25'b0000000000001011011100000;
    rom[54945] = 25'b0000000000001011011110101;
    rom[54946] = 25'b0000000000001011100001010;
    rom[54947] = 25'b0000000000001011100011111;
    rom[54948] = 25'b0000000000001011100110100;
    rom[54949] = 25'b0000000000001011101001010;
    rom[54950] = 25'b0000000000001011101011111;
    rom[54951] = 25'b0000000000001011101110100;
    rom[54952] = 25'b0000000000001011110001001;
    rom[54953] = 25'b0000000000001011110011110;
    rom[54954] = 25'b0000000000001011110110011;
    rom[54955] = 25'b0000000000001011111001000;
    rom[54956] = 25'b0000000000001011111011101;
    rom[54957] = 25'b0000000000001011111110010;
    rom[54958] = 25'b0000000000001100000000111;
    rom[54959] = 25'b0000000000001100000011100;
    rom[54960] = 25'b0000000000001100000110001;
    rom[54961] = 25'b0000000000001100001000110;
    rom[54962] = 25'b0000000000001100001011011;
    rom[54963] = 25'b0000000000001100001110000;
    rom[54964] = 25'b0000000000001100010000101;
    rom[54965] = 25'b0000000000001100010011010;
    rom[54966] = 25'b0000000000001100010101110;
    rom[54967] = 25'b0000000000001100011000011;
    rom[54968] = 25'b0000000000001100011011000;
    rom[54969] = 25'b0000000000001100011101100;
    rom[54970] = 25'b0000000000001100100000001;
    rom[54971] = 25'b0000000000001100100010110;
    rom[54972] = 25'b0000000000001100100101010;
    rom[54973] = 25'b0000000000001100100111111;
    rom[54974] = 25'b0000000000001100101010100;
    rom[54975] = 25'b0000000000001100101101000;
    rom[54976] = 25'b0000000000001100101111101;
    rom[54977] = 25'b0000000000001100110010010;
    rom[54978] = 25'b0000000000001100110100110;
    rom[54979] = 25'b0000000000001100110111010;
    rom[54980] = 25'b0000000000001100111001111;
    rom[54981] = 25'b0000000000001100111100011;
    rom[54982] = 25'b0000000000001100111111000;
    rom[54983] = 25'b0000000000001101000001100;
    rom[54984] = 25'b0000000000001101000100000;
    rom[54985] = 25'b0000000000001101000110100;
    rom[54986] = 25'b0000000000001101001001001;
    rom[54987] = 25'b0000000000001101001011110;
    rom[54988] = 25'b0000000000001101001110010;
    rom[54989] = 25'b0000000000001101010000110;
    rom[54990] = 25'b0000000000001101010011010;
    rom[54991] = 25'b0000000000001101010101110;
    rom[54992] = 25'b0000000000001101011000010;
    rom[54993] = 25'b0000000000001101011010111;
    rom[54994] = 25'b0000000000001101011101011;
    rom[54995] = 25'b0000000000001101011111111;
    rom[54996] = 25'b0000000000001101100010011;
    rom[54997] = 25'b0000000000001101100100111;
    rom[54998] = 25'b0000000000001101100111011;
    rom[54999] = 25'b0000000000001101101001111;
    rom[55000] = 25'b0000000000001101101100011;
    rom[55001] = 25'b0000000000001101101110111;
    rom[55002] = 25'b0000000000001101110001011;
    rom[55003] = 25'b0000000000001101110011111;
    rom[55004] = 25'b0000000000001101110110011;
    rom[55005] = 25'b0000000000001101111000111;
    rom[55006] = 25'b0000000000001101111011011;
    rom[55007] = 25'b0000000000001101111101111;
    rom[55008] = 25'b0000000000001110000000010;
    rom[55009] = 25'b0000000000001110000010110;
    rom[55010] = 25'b0000000000001110000101010;
    rom[55011] = 25'b0000000000001110000111110;
    rom[55012] = 25'b0000000000001110001010001;
    rom[55013] = 25'b0000000000001110001100101;
    rom[55014] = 25'b0000000000001110001111001;
    rom[55015] = 25'b0000000000001110010001100;
    rom[55016] = 25'b0000000000001110010100000;
    rom[55017] = 25'b0000000000001110010110100;
    rom[55018] = 25'b0000000000001110011000111;
    rom[55019] = 25'b0000000000001110011011011;
    rom[55020] = 25'b0000000000001110011101110;
    rom[55021] = 25'b0000000000001110100000010;
    rom[55022] = 25'b0000000000001110100010101;
    rom[55023] = 25'b0000000000001110100101000;
    rom[55024] = 25'b0000000000001110100111100;
    rom[55025] = 25'b0000000000001110101001111;
    rom[55026] = 25'b0000000000001110101100011;
    rom[55027] = 25'b0000000000001110101110110;
    rom[55028] = 25'b0000000000001110110001010;
    rom[55029] = 25'b0000000000001110110011101;
    rom[55030] = 25'b0000000000001110110110000;
    rom[55031] = 25'b0000000000001110111000100;
    rom[55032] = 25'b0000000000001110111010111;
    rom[55033] = 25'b0000000000001110111101010;
    rom[55034] = 25'b0000000000001110111111101;
    rom[55035] = 25'b0000000000001111000010000;
    rom[55036] = 25'b0000000000001111000100100;
    rom[55037] = 25'b0000000000001111000110111;
    rom[55038] = 25'b0000000000001111001001010;
    rom[55039] = 25'b0000000000001111001011101;
    rom[55040] = 25'b0000000000001111001110000;
    rom[55041] = 25'b0000000000001111010000011;
    rom[55042] = 25'b0000000000001111010010110;
    rom[55043] = 25'b0000000000001111010101001;
    rom[55044] = 25'b0000000000001111010111100;
    rom[55045] = 25'b0000000000001111011001111;
    rom[55046] = 25'b0000000000001111011100010;
    rom[55047] = 25'b0000000000001111011110101;
    rom[55048] = 25'b0000000000001111100000111;
    rom[55049] = 25'b0000000000001111100011011;
    rom[55050] = 25'b0000000000001111100101101;
    rom[55051] = 25'b0000000000001111101000000;
    rom[55052] = 25'b0000000000001111101010011;
    rom[55053] = 25'b0000000000001111101100110;
    rom[55054] = 25'b0000000000001111101111000;
    rom[55055] = 25'b0000000000001111110001011;
    rom[55056] = 25'b0000000000001111110011110;
    rom[55057] = 25'b0000000000001111110110000;
    rom[55058] = 25'b0000000000001111111000011;
    rom[55059] = 25'b0000000000001111111010110;
    rom[55060] = 25'b0000000000001111111101000;
    rom[55061] = 25'b0000000000001111111111011;
    rom[55062] = 25'b0000000000010000000001110;
    rom[55063] = 25'b0000000000010000000100000;
    rom[55064] = 25'b0000000000010000000110010;
    rom[55065] = 25'b0000000000010000001000101;
    rom[55066] = 25'b0000000000010000001011000;
    rom[55067] = 25'b0000000000010000001101001;
    rom[55068] = 25'b0000000000010000001111100;
    rom[55069] = 25'b0000000000010000010001110;
    rom[55070] = 25'b0000000000010000010100001;
    rom[55071] = 25'b0000000000010000010110011;
    rom[55072] = 25'b0000000000010000011000101;
    rom[55073] = 25'b0000000000010000011010111;
    rom[55074] = 25'b0000000000010000011101010;
    rom[55075] = 25'b0000000000010000011111100;
    rom[55076] = 25'b0000000000010000100001111;
    rom[55077] = 25'b0000000000010000100100001;
    rom[55078] = 25'b0000000000010000100110010;
    rom[55079] = 25'b0000000000010000101000100;
    rom[55080] = 25'b0000000000010000101010111;
    rom[55081] = 25'b0000000000010000101101001;
    rom[55082] = 25'b0000000000010000101111011;
    rom[55083] = 25'b0000000000010000110001101;
    rom[55084] = 25'b0000000000010000110011111;
    rom[55085] = 25'b0000000000010000110110001;
    rom[55086] = 25'b0000000000010000111000011;
    rom[55087] = 25'b0000000000010000111010101;
    rom[55088] = 25'b0000000000010000111100111;
    rom[55089] = 25'b0000000000010000111111000;
    rom[55090] = 25'b0000000000010001000001010;
    rom[55091] = 25'b0000000000010001000011100;
    rom[55092] = 25'b0000000000010001000101110;
    rom[55093] = 25'b0000000000010001001000000;
    rom[55094] = 25'b0000000000010001001010001;
    rom[55095] = 25'b0000000000010001001100011;
    rom[55096] = 25'b0000000000010001001110101;
    rom[55097] = 25'b0000000000010001010000111;
    rom[55098] = 25'b0000000000010001010011000;
    rom[55099] = 25'b0000000000010001010101010;
    rom[55100] = 25'b0000000000010001010111011;
    rom[55101] = 25'b0000000000010001011001101;
    rom[55102] = 25'b0000000000010001011011111;
    rom[55103] = 25'b0000000000010001011110000;
    rom[55104] = 25'b0000000000010001100000010;
    rom[55105] = 25'b0000000000010001100010100;
    rom[55106] = 25'b0000000000010001100100101;
    rom[55107] = 25'b0000000000010001100110111;
    rom[55108] = 25'b0000000000010001101001000;
    rom[55109] = 25'b0000000000010001101011001;
    rom[55110] = 25'b0000000000010001101101010;
    rom[55111] = 25'b0000000000010001101111100;
    rom[55112] = 25'b0000000000010001110001101;
    rom[55113] = 25'b0000000000010001110011111;
    rom[55114] = 25'b0000000000010001110110000;
    rom[55115] = 25'b0000000000010001111000001;
    rom[55116] = 25'b0000000000010001111010010;
    rom[55117] = 25'b0000000000010001111100011;
    rom[55118] = 25'b0000000000010001111110100;
    rom[55119] = 25'b0000000000010010000000110;
    rom[55120] = 25'b0000000000010010000010111;
    rom[55121] = 25'b0000000000010010000101000;
    rom[55122] = 25'b0000000000010010000111001;
    rom[55123] = 25'b0000000000010010001001010;
    rom[55124] = 25'b0000000000010010001011011;
    rom[55125] = 25'b0000000000010010001101100;
    rom[55126] = 25'b0000000000010010001111101;
    rom[55127] = 25'b0000000000010010010001110;
    rom[55128] = 25'b0000000000010010010011111;
    rom[55129] = 25'b0000000000010010010110000;
    rom[55130] = 25'b0000000000010010011000001;
    rom[55131] = 25'b0000000000010010011010010;
    rom[55132] = 25'b0000000000010010011100011;
    rom[55133] = 25'b0000000000010010011110011;
    rom[55134] = 25'b0000000000010010100000100;
    rom[55135] = 25'b0000000000010010100010101;
    rom[55136] = 25'b0000000000010010100100101;
    rom[55137] = 25'b0000000000010010100110110;
    rom[55138] = 25'b0000000000010010101000111;
    rom[55139] = 25'b0000000000010010101010111;
    rom[55140] = 25'b0000000000010010101101001;
    rom[55141] = 25'b0000000000010010101111001;
    rom[55142] = 25'b0000000000010010110001001;
    rom[55143] = 25'b0000000000010010110011010;
    rom[55144] = 25'b0000000000010010110101010;
    rom[55145] = 25'b0000000000010010110111011;
    rom[55146] = 25'b0000000000010010111001100;
    rom[55147] = 25'b0000000000010010111011100;
    rom[55148] = 25'b0000000000010010111101101;
    rom[55149] = 25'b0000000000010010111111100;
    rom[55150] = 25'b0000000000010011000001101;
    rom[55151] = 25'b0000000000010011000011101;
    rom[55152] = 25'b0000000000010011000101110;
    rom[55153] = 25'b0000000000010011000111110;
    rom[55154] = 25'b0000000000010011001001111;
    rom[55155] = 25'b0000000000010011001011111;
    rom[55156] = 25'b0000000000010011001101111;
    rom[55157] = 25'b0000000000010011001111111;
    rom[55158] = 25'b0000000000010011010010000;
    rom[55159] = 25'b0000000000010011010011111;
    rom[55160] = 25'b0000000000010011010110000;
    rom[55161] = 25'b0000000000010011010111111;
    rom[55162] = 25'b0000000000010011011010000;
    rom[55163] = 25'b0000000000010011011100000;
    rom[55164] = 25'b0000000000010011011110000;
    rom[55165] = 25'b0000000000010011100000000;
    rom[55166] = 25'b0000000000010011100010000;
    rom[55167] = 25'b0000000000010011100100000;
    rom[55168] = 25'b0000000000010011100110000;
    rom[55169] = 25'b0000000000010011101000000;
    rom[55170] = 25'b0000000000010011101010000;
    rom[55171] = 25'b0000000000010011101011111;
    rom[55172] = 25'b0000000000010011101101111;
    rom[55173] = 25'b0000000000010011101111111;
    rom[55174] = 25'b0000000000010011110001111;
    rom[55175] = 25'b0000000000010011110011111;
    rom[55176] = 25'b0000000000010011110101111;
    rom[55177] = 25'b0000000000010011110111110;
    rom[55178] = 25'b0000000000010011111001110;
    rom[55179] = 25'b0000000000010011111011110;
    rom[55180] = 25'b0000000000010011111101101;
    rom[55181] = 25'b0000000000010011111111101;
    rom[55182] = 25'b0000000000010100000001101;
    rom[55183] = 25'b0000000000010100000011100;
    rom[55184] = 25'b0000000000010100000101011;
    rom[55185] = 25'b0000000000010100000111011;
    rom[55186] = 25'b0000000000010100001001011;
    rom[55187] = 25'b0000000000010100001011010;
    rom[55188] = 25'b0000000000010100001101001;
    rom[55189] = 25'b0000000000010100001111001;
    rom[55190] = 25'b0000000000010100010001000;
    rom[55191] = 25'b0000000000010100010011000;
    rom[55192] = 25'b0000000000010100010100111;
    rom[55193] = 25'b0000000000010100010110110;
    rom[55194] = 25'b0000000000010100011000101;
    rom[55195] = 25'b0000000000010100011010101;
    rom[55196] = 25'b0000000000010100011100100;
    rom[55197] = 25'b0000000000010100011110011;
    rom[55198] = 25'b0000000000010100100000010;
    rom[55199] = 25'b0000000000010100100010001;
    rom[55200] = 25'b0000000000010100100100000;
    rom[55201] = 25'b0000000000010100100110000;
    rom[55202] = 25'b0000000000010100100111111;
    rom[55203] = 25'b0000000000010100101001110;
    rom[55204] = 25'b0000000000010100101011101;
    rom[55205] = 25'b0000000000010100101101100;
    rom[55206] = 25'b0000000000010100101111011;
    rom[55207] = 25'b0000000000010100110001010;
    rom[55208] = 25'b0000000000010100110011001;
    rom[55209] = 25'b0000000000010100110101000;
    rom[55210] = 25'b0000000000010100110110110;
    rom[55211] = 25'b0000000000010100111000101;
    rom[55212] = 25'b0000000000010100111010100;
    rom[55213] = 25'b0000000000010100111100011;
    rom[55214] = 25'b0000000000010100111110010;
    rom[55215] = 25'b0000000000010101000000000;
    rom[55216] = 25'b0000000000010101000001111;
    rom[55217] = 25'b0000000000010101000011110;
    rom[55218] = 25'b0000000000010101000101101;
    rom[55219] = 25'b0000000000010101000111011;
    rom[55220] = 25'b0000000000010101001001010;
    rom[55221] = 25'b0000000000010101001011001;
    rom[55222] = 25'b0000000000010101001100111;
    rom[55223] = 25'b0000000000010101001110110;
    rom[55224] = 25'b0000000000010101010000100;
    rom[55225] = 25'b0000000000010101010010011;
    rom[55226] = 25'b0000000000010101010100001;
    rom[55227] = 25'b0000000000010101010110000;
    rom[55228] = 25'b0000000000010101010111110;
    rom[55229] = 25'b0000000000010101011001100;
    rom[55230] = 25'b0000000000010101011011011;
    rom[55231] = 25'b0000000000010101011101010;
    rom[55232] = 25'b0000000000010101011111000;
    rom[55233] = 25'b0000000000010101100000110;
    rom[55234] = 25'b0000000000010101100010100;
    rom[55235] = 25'b0000000000010101100100010;
    rom[55236] = 25'b0000000000010101100110001;
    rom[55237] = 25'b0000000000010101100111111;
    rom[55238] = 25'b0000000000010101101001101;
    rom[55239] = 25'b0000000000010101101011011;
    rom[55240] = 25'b0000000000010101101101001;
    rom[55241] = 25'b0000000000010101101110111;
    rom[55242] = 25'b0000000000010101110000110;
    rom[55243] = 25'b0000000000010101110010011;
    rom[55244] = 25'b0000000000010101110100001;
    rom[55245] = 25'b0000000000010101110110000;
    rom[55246] = 25'b0000000000010101110111110;
    rom[55247] = 25'b0000000000010101111001011;
    rom[55248] = 25'b0000000000010101111011001;
    rom[55249] = 25'b0000000000010101111101000;
    rom[55250] = 25'b0000000000010101111110101;
    rom[55251] = 25'b0000000000010110000000011;
    rom[55252] = 25'b0000000000010110000010001;
    rom[55253] = 25'b0000000000010110000011111;
    rom[55254] = 25'b0000000000010110000101100;
    rom[55255] = 25'b0000000000010110000111010;
    rom[55256] = 25'b0000000000010110001001000;
    rom[55257] = 25'b0000000000010110001010101;
    rom[55258] = 25'b0000000000010110001100011;
    rom[55259] = 25'b0000000000010110001110001;
    rom[55260] = 25'b0000000000010110001111110;
    rom[55261] = 25'b0000000000010110010001100;
    rom[55262] = 25'b0000000000010110010011001;
    rom[55263] = 25'b0000000000010110010100111;
    rom[55264] = 25'b0000000000010110010110100;
    rom[55265] = 25'b0000000000010110011000010;
    rom[55266] = 25'b0000000000010110011010000;
    rom[55267] = 25'b0000000000010110011011101;
    rom[55268] = 25'b0000000000010110011101011;
    rom[55269] = 25'b0000000000010110011111000;
    rom[55270] = 25'b0000000000010110100000101;
    rom[55271] = 25'b0000000000010110100010010;
    rom[55272] = 25'b0000000000010110100100000;
    rom[55273] = 25'b0000000000010110100101101;
    rom[55274] = 25'b0000000000010110100111011;
    rom[55275] = 25'b0000000000010110101000111;
    rom[55276] = 25'b0000000000010110101010101;
    rom[55277] = 25'b0000000000010110101100010;
    rom[55278] = 25'b0000000000010110101101111;
    rom[55279] = 25'b0000000000010110101111100;
    rom[55280] = 25'b0000000000010110110001001;
    rom[55281] = 25'b0000000000010110110010111;
    rom[55282] = 25'b0000000000010110110100011;
    rom[55283] = 25'b0000000000010110110110001;
    rom[55284] = 25'b0000000000010110110111101;
    rom[55285] = 25'b0000000000010110111001011;
    rom[55286] = 25'b0000000000010110111011000;
    rom[55287] = 25'b0000000000010110111100100;
    rom[55288] = 25'b0000000000010110111110001;
    rom[55289] = 25'b0000000000010110111111110;
    rom[55290] = 25'b0000000000010111000001011;
    rom[55291] = 25'b0000000000010111000011000;
    rom[55292] = 25'b0000000000010111000100101;
    rom[55293] = 25'b0000000000010111000110001;
    rom[55294] = 25'b0000000000010111000111110;
    rom[55295] = 25'b0000000000010111001001011;
    rom[55296] = 25'b0000000000010111001010111;
    rom[55297] = 25'b0000000000010111001100100;
    rom[55298] = 25'b0000000000010111001110001;
    rom[55299] = 25'b0000000000010111001111101;
    rom[55300] = 25'b0000000000010111010001010;
    rom[55301] = 25'b0000000000010111010010111;
    rom[55302] = 25'b0000000000010111010100100;
    rom[55303] = 25'b0000000000010111010110000;
    rom[55304] = 25'b0000000000010111010111100;
    rom[55305] = 25'b0000000000010111011001001;
    rom[55306] = 25'b0000000000010111011010101;
    rom[55307] = 25'b0000000000010111011100010;
    rom[55308] = 25'b0000000000010111011101110;
    rom[55309] = 25'b0000000000010111011111010;
    rom[55310] = 25'b0000000000010111100000111;
    rom[55311] = 25'b0000000000010111100010011;
    rom[55312] = 25'b0000000000010111100100000;
    rom[55313] = 25'b0000000000010111100101100;
    rom[55314] = 25'b0000000000010111100111000;
    rom[55315] = 25'b0000000000010111101000100;
    rom[55316] = 25'b0000000000010111101010000;
    rom[55317] = 25'b0000000000010111101011100;
    rom[55318] = 25'b0000000000010111101101001;
    rom[55319] = 25'b0000000000010111101110101;
    rom[55320] = 25'b0000000000010111110000001;
    rom[55321] = 25'b0000000000010111110001101;
    rom[55322] = 25'b0000000000010111110011001;
    rom[55323] = 25'b0000000000010111110100101;
    rom[55324] = 25'b0000000000010111110110001;
    rom[55325] = 25'b0000000000010111110111101;
    rom[55326] = 25'b0000000000010111111001000;
    rom[55327] = 25'b0000000000010111111010100;
    rom[55328] = 25'b0000000000010111111100000;
    rom[55329] = 25'b0000000000010111111101100;
    rom[55330] = 25'b0000000000010111111111000;
    rom[55331] = 25'b0000000000011000000000100;
    rom[55332] = 25'b0000000000011000000010000;
    rom[55333] = 25'b0000000000011000000011011;
    rom[55334] = 25'b0000000000011000000100111;
    rom[55335] = 25'b0000000000011000000110011;
    rom[55336] = 25'b0000000000011000000111110;
    rom[55337] = 25'b0000000000011000001001010;
    rom[55338] = 25'b0000000000011000001010110;
    rom[55339] = 25'b0000000000011000001100010;
    rom[55340] = 25'b0000000000011000001101110;
    rom[55341] = 25'b0000000000011000001111001;
    rom[55342] = 25'b0000000000011000010000100;
    rom[55343] = 25'b0000000000011000010010000;
    rom[55344] = 25'b0000000000011000010011011;
    rom[55345] = 25'b0000000000011000010100111;
    rom[55346] = 25'b0000000000011000010110010;
    rom[55347] = 25'b0000000000011000010111101;
    rom[55348] = 25'b0000000000011000011001001;
    rom[55349] = 25'b0000000000011000011010100;
    rom[55350] = 25'b0000000000011000011100000;
    rom[55351] = 25'b0000000000011000011101011;
    rom[55352] = 25'b0000000000011000011110110;
    rom[55353] = 25'b0000000000011000100000001;
    rom[55354] = 25'b0000000000011000100001101;
    rom[55355] = 25'b0000000000011000100011000;
    rom[55356] = 25'b0000000000011000100100011;
    rom[55357] = 25'b0000000000011000100101110;
    rom[55358] = 25'b0000000000011000100111010;
    rom[55359] = 25'b0000000000011000101000101;
    rom[55360] = 25'b0000000000011000101001111;
    rom[55361] = 25'b0000000000011000101011010;
    rom[55362] = 25'b0000000000011000101100110;
    rom[55363] = 25'b0000000000011000101110001;
    rom[55364] = 25'b0000000000011000101111011;
    rom[55365] = 25'b0000000000011000110000110;
    rom[55366] = 25'b0000000000011000110010001;
    rom[55367] = 25'b0000000000011000110011100;
    rom[55368] = 25'b0000000000011000110100111;
    rom[55369] = 25'b0000000000011000110110010;
    rom[55370] = 25'b0000000000011000110111101;
    rom[55371] = 25'b0000000000011000111000111;
    rom[55372] = 25'b0000000000011000111010010;
    rom[55373] = 25'b0000000000011000111011101;
    rom[55374] = 25'b0000000000011000111101000;
    rom[55375] = 25'b0000000000011000111110010;
    rom[55376] = 25'b0000000000011000111111101;
    rom[55377] = 25'b0000000000011001000001000;
    rom[55378] = 25'b0000000000011001000010010;
    rom[55379] = 25'b0000000000011001000011101;
    rom[55380] = 25'b0000000000011001000100111;
    rom[55381] = 25'b0000000000011001000110010;
    rom[55382] = 25'b0000000000011001000111101;
    rom[55383] = 25'b0000000000011001001000111;
    rom[55384] = 25'b0000000000011001001010010;
    rom[55385] = 25'b0000000000011001001011100;
    rom[55386] = 25'b0000000000011001001100110;
    rom[55387] = 25'b0000000000011001001110000;
    rom[55388] = 25'b0000000000011001001111011;
    rom[55389] = 25'b0000000000011001010000101;
    rom[55390] = 25'b0000000000011001010010000;
    rom[55391] = 25'b0000000000011001010011010;
    rom[55392] = 25'b0000000000011001010100100;
    rom[55393] = 25'b0000000000011001010101110;
    rom[55394] = 25'b0000000000011001010111001;
    rom[55395] = 25'b0000000000011001011000010;
    rom[55396] = 25'b0000000000011001011001101;
    rom[55397] = 25'b0000000000011001011010111;
    rom[55398] = 25'b0000000000011001011100001;
    rom[55399] = 25'b0000000000011001011101011;
    rom[55400] = 25'b0000000000011001011110101;
    rom[55401] = 25'b0000000000011001011111111;
    rom[55402] = 25'b0000000000011001100001001;
    rom[55403] = 25'b0000000000011001100010011;
    rom[55404] = 25'b0000000000011001100011101;
    rom[55405] = 25'b0000000000011001100100111;
    rom[55406] = 25'b0000000000011001100110001;
    rom[55407] = 25'b0000000000011001100111011;
    rom[55408] = 25'b0000000000011001101000100;
    rom[55409] = 25'b0000000000011001101001110;
    rom[55410] = 25'b0000000000011001101011001;
    rom[55411] = 25'b0000000000011001101100010;
    rom[55412] = 25'b0000000000011001101101100;
    rom[55413] = 25'b0000000000011001101110110;
    rom[55414] = 25'b0000000000011001110000000;
    rom[55415] = 25'b0000000000011001110001001;
    rom[55416] = 25'b0000000000011001110010010;
    rom[55417] = 25'b0000000000011001110011100;
    rom[55418] = 25'b0000000000011001110100110;
    rom[55419] = 25'b0000000000011001110101111;
    rom[55420] = 25'b0000000000011001110111001;
    rom[55421] = 25'b0000000000011001111000010;
    rom[55422] = 25'b0000000000011001111001100;
    rom[55423] = 25'b0000000000011001111010101;
    rom[55424] = 25'b0000000000011001111011110;
    rom[55425] = 25'b0000000000011001111101000;
    rom[55426] = 25'b0000000000011001111110010;
    rom[55427] = 25'b0000000000011001111111011;
    rom[55428] = 25'b0000000000011010000000100;
    rom[55429] = 25'b0000000000011010000001101;
    rom[55430] = 25'b0000000000011010000010111;
    rom[55431] = 25'b0000000000011010000100000;
    rom[55432] = 25'b0000000000011010000101001;
    rom[55433] = 25'b0000000000011010000110011;
    rom[55434] = 25'b0000000000011010000111100;
    rom[55435] = 25'b0000000000011010001000101;
    rom[55436] = 25'b0000000000011010001001110;
    rom[55437] = 25'b0000000000011010001010111;
    rom[55438] = 25'b0000000000011010001100000;
    rom[55439] = 25'b0000000000011010001101001;
    rom[55440] = 25'b0000000000011010001110010;
    rom[55441] = 25'b0000000000011010001111011;
    rom[55442] = 25'b0000000000011010010000100;
    rom[55443] = 25'b0000000000011010010001101;
    rom[55444] = 25'b0000000000011010010010110;
    rom[55445] = 25'b0000000000011010010011111;
    rom[55446] = 25'b0000000000011010010101000;
    rom[55447] = 25'b0000000000011010010110001;
    rom[55448] = 25'b0000000000011010010111001;
    rom[55449] = 25'b0000000000011010011000010;
    rom[55450] = 25'b0000000000011010011001011;
    rom[55451] = 25'b0000000000011010011010100;
    rom[55452] = 25'b0000000000011010011011100;
    rom[55453] = 25'b0000000000011010011100101;
    rom[55454] = 25'b0000000000011010011101110;
    rom[55455] = 25'b0000000000011010011110111;
    rom[55456] = 25'b0000000000011010100000000;
    rom[55457] = 25'b0000000000011010100001000;
    rom[55458] = 25'b0000000000011010100010001;
    rom[55459] = 25'b0000000000011010100011001;
    rom[55460] = 25'b0000000000011010100100010;
    rom[55461] = 25'b0000000000011010100101010;
    rom[55462] = 25'b0000000000011010100110010;
    rom[55463] = 25'b0000000000011010100111011;
    rom[55464] = 25'b0000000000011010101000011;
    rom[55465] = 25'b0000000000011010101001100;
    rom[55466] = 25'b0000000000011010101010100;
    rom[55467] = 25'b0000000000011010101011101;
    rom[55468] = 25'b0000000000011010101100101;
    rom[55469] = 25'b0000000000011010101101101;
    rom[55470] = 25'b0000000000011010101110110;
    rom[55471] = 25'b0000000000011010101111110;
    rom[55472] = 25'b0000000000011010110000110;
    rom[55473] = 25'b0000000000011010110001110;
    rom[55474] = 25'b0000000000011010110010110;
    rom[55475] = 25'b0000000000011010110011111;
    rom[55476] = 25'b0000000000011010110100111;
    rom[55477] = 25'b0000000000011010110101110;
    rom[55478] = 25'b0000000000011010110110111;
    rom[55479] = 25'b0000000000011010110111111;
    rom[55480] = 25'b0000000000011010111000111;
    rom[55481] = 25'b0000000000011010111001111;
    rom[55482] = 25'b0000000000011010111010111;
    rom[55483] = 25'b0000000000011010111011111;
    rom[55484] = 25'b0000000000011010111100110;
    rom[55485] = 25'b0000000000011010111101111;
    rom[55486] = 25'b0000000000011010111110111;
    rom[55487] = 25'b0000000000011010111111110;
    rom[55488] = 25'b0000000000011011000000110;
    rom[55489] = 25'b0000000000011011000001110;
    rom[55490] = 25'b0000000000011011000010101;
    rom[55491] = 25'b0000000000011011000011110;
    rom[55492] = 25'b0000000000011011000100101;
    rom[55493] = 25'b0000000000011011000101101;
    rom[55494] = 25'b0000000000011011000110101;
    rom[55495] = 25'b0000000000011011000111100;
    rom[55496] = 25'b0000000000011011001000100;
    rom[55497] = 25'b0000000000011011001001011;
    rom[55498] = 25'b0000000000011011001010011;
    rom[55499] = 25'b0000000000011011001011010;
    rom[55500] = 25'b0000000000011011001100010;
    rom[55501] = 25'b0000000000011011001101010;
    rom[55502] = 25'b0000000000011011001110001;
    rom[55503] = 25'b0000000000011011001111000;
    rom[55504] = 25'b0000000000011011010000000;
    rom[55505] = 25'b0000000000011011010000111;
    rom[55506] = 25'b0000000000011011010001110;
    rom[55507] = 25'b0000000000011011010010110;
    rom[55508] = 25'b0000000000011011010011101;
    rom[55509] = 25'b0000000000011011010100101;
    rom[55510] = 25'b0000000000011011010101100;
    rom[55511] = 25'b0000000000011011010110011;
    rom[55512] = 25'b0000000000011011010111011;
    rom[55513] = 25'b0000000000011011011000001;
    rom[55514] = 25'b0000000000011011011001001;
    rom[55515] = 25'b0000000000011011011001111;
    rom[55516] = 25'b0000000000011011011010111;
    rom[55517] = 25'b0000000000011011011011110;
    rom[55518] = 25'b0000000000011011011100101;
    rom[55519] = 25'b0000000000011011011101100;
    rom[55520] = 25'b0000000000011011011110011;
    rom[55521] = 25'b0000000000011011011111010;
    rom[55522] = 25'b0000000000011011100000001;
    rom[55523] = 25'b0000000000011011100001000;
    rom[55524] = 25'b0000000000011011100001111;
    rom[55525] = 25'b0000000000011011100010110;
    rom[55526] = 25'b0000000000011011100011100;
    rom[55527] = 25'b0000000000011011100100100;
    rom[55528] = 25'b0000000000011011100101011;
    rom[55529] = 25'b0000000000011011100110001;
    rom[55530] = 25'b0000000000011011100111000;
    rom[55531] = 25'b0000000000011011100111111;
    rom[55532] = 25'b0000000000011011101000110;
    rom[55533] = 25'b0000000000011011101001100;
    rom[55534] = 25'b0000000000011011101010011;
    rom[55535] = 25'b0000000000011011101011010;
    rom[55536] = 25'b0000000000011011101100000;
    rom[55537] = 25'b0000000000011011101100110;
    rom[55538] = 25'b0000000000011011101101101;
    rom[55539] = 25'b0000000000011011101110100;
    rom[55540] = 25'b0000000000011011101111011;
    rom[55541] = 25'b0000000000011011110000001;
    rom[55542] = 25'b0000000000011011110000111;
    rom[55543] = 25'b0000000000011011110001110;
    rom[55544] = 25'b0000000000011011110010100;
    rom[55545] = 25'b0000000000011011110011011;
    rom[55546] = 25'b0000000000011011110100001;
    rom[55547] = 25'b0000000000011011110100111;
    rom[55548] = 25'b0000000000011011110101101;
    rom[55549] = 25'b0000000000011011110110100;
    rom[55550] = 25'b0000000000011011110111010;
    rom[55551] = 25'b0000000000011011111000001;
    rom[55552] = 25'b0000000000011011111000111;
    rom[55553] = 25'b0000000000011011111001101;
    rom[55554] = 25'b0000000000011011111010011;
    rom[55555] = 25'b0000000000011011111011001;
    rom[55556] = 25'b0000000000011011111011111;
    rom[55557] = 25'b0000000000011011111100101;
    rom[55558] = 25'b0000000000011011111101011;
    rom[55559] = 25'b0000000000011011111110001;
    rom[55560] = 25'b0000000000011011111110111;
    rom[55561] = 25'b0000000000011011111111101;
    rom[55562] = 25'b0000000000011100000000011;
    rom[55563] = 25'b0000000000011100000001001;
    rom[55564] = 25'b0000000000011100000001111;
    rom[55565] = 25'b0000000000011100000010101;
    rom[55566] = 25'b0000000000011100000011011;
    rom[55567] = 25'b0000000000011100000100001;
    rom[55568] = 25'b0000000000011100000100111;
    rom[55569] = 25'b0000000000011100000101101;
    rom[55570] = 25'b0000000000011100000110010;
    rom[55571] = 25'b0000000000011100000111000;
    rom[55572] = 25'b0000000000011100000111110;
    rom[55573] = 25'b0000000000011100001000100;
    rom[55574] = 25'b0000000000011100001001001;
    rom[55575] = 25'b0000000000011100001001111;
    rom[55576] = 25'b0000000000011100001010101;
    rom[55577] = 25'b0000000000011100001011011;
    rom[55578] = 25'b0000000000011100001100000;
    rom[55579] = 25'b0000000000011100001100101;
    rom[55580] = 25'b0000000000011100001101011;
    rom[55581] = 25'b0000000000011100001110000;
    rom[55582] = 25'b0000000000011100001110110;
    rom[55583] = 25'b0000000000011100001111100;
    rom[55584] = 25'b0000000000011100010000001;
    rom[55585] = 25'b0000000000011100010000110;
    rom[55586] = 25'b0000000000011100010001100;
    rom[55587] = 25'b0000000000011100010010001;
    rom[55588] = 25'b0000000000011100010010110;
    rom[55589] = 25'b0000000000011100010011100;
    rom[55590] = 25'b0000000000011100010100001;
    rom[55591] = 25'b0000000000011100010100110;
    rom[55592] = 25'b0000000000011100010101011;
    rom[55593] = 25'b0000000000011100010110001;
    rom[55594] = 25'b0000000000011100010110110;
    rom[55595] = 25'b0000000000011100010111011;
    rom[55596] = 25'b0000000000011100011000000;
    rom[55597] = 25'b0000000000011100011000110;
    rom[55598] = 25'b0000000000011100011001011;
    rom[55599] = 25'b0000000000011100011001111;
    rom[55600] = 25'b0000000000011100011010100;
    rom[55601] = 25'b0000000000011100011011010;
    rom[55602] = 25'b0000000000011100011011111;
    rom[55603] = 25'b0000000000011100011100011;
    rom[55604] = 25'b0000000000011100011101001;
    rom[55605] = 25'b0000000000011100011101110;
    rom[55606] = 25'b0000000000011100011110010;
    rom[55607] = 25'b0000000000011100011111000;
    rom[55608] = 25'b0000000000011100011111100;
    rom[55609] = 25'b0000000000011100100000001;
    rom[55610] = 25'b0000000000011100100000110;
    rom[55611] = 25'b0000000000011100100001010;
    rom[55612] = 25'b0000000000011100100001111;
    rom[55613] = 25'b0000000000011100100010100;
    rom[55614] = 25'b0000000000011100100011000;
    rom[55615] = 25'b0000000000011100100011110;
    rom[55616] = 25'b0000000000011100100100010;
    rom[55617] = 25'b0000000000011100100100111;
    rom[55618] = 25'b0000000000011100100101011;
    rom[55619] = 25'b0000000000011100100110000;
    rom[55620] = 25'b0000000000011100100110101;
    rom[55621] = 25'b0000000000011100100111001;
    rom[55622] = 25'b0000000000011100100111110;
    rom[55623] = 25'b0000000000011100101000010;
    rom[55624] = 25'b0000000000011100101000111;
    rom[55625] = 25'b0000000000011100101001011;
    rom[55626] = 25'b0000000000011100101010000;
    rom[55627] = 25'b0000000000011100101010011;
    rom[55628] = 25'b0000000000011100101011000;
    rom[55629] = 25'b0000000000011100101011100;
    rom[55630] = 25'b0000000000011100101100001;
    rom[55631] = 25'b0000000000011100101100101;
    rom[55632] = 25'b0000000000011100101101001;
    rom[55633] = 25'b0000000000011100101101110;
    rom[55634] = 25'b0000000000011100101110010;
    rom[55635] = 25'b0000000000011100101110110;
    rom[55636] = 25'b0000000000011100101111010;
    rom[55637] = 25'b0000000000011100101111111;
    rom[55638] = 25'b0000000000011100110000011;
    rom[55639] = 25'b0000000000011100110000111;
    rom[55640] = 25'b0000000000011100110001011;
    rom[55641] = 25'b0000000000011100110001110;
    rom[55642] = 25'b0000000000011100110010011;
    rom[55643] = 25'b0000000000011100110010111;
    rom[55644] = 25'b0000000000011100110011011;
    rom[55645] = 25'b0000000000011100110011111;
    rom[55646] = 25'b0000000000011100110100011;
    rom[55647] = 25'b0000000000011100110100110;
    rom[55648] = 25'b0000000000011100110101011;
    rom[55649] = 25'b0000000000011100110101111;
    rom[55650] = 25'b0000000000011100110110010;
    rom[55651] = 25'b0000000000011100110110110;
    rom[55652] = 25'b0000000000011100110111010;
    rom[55653] = 25'b0000000000011100110111110;
    rom[55654] = 25'b0000000000011100111000001;
    rom[55655] = 25'b0000000000011100111000101;
    rom[55656] = 25'b0000000000011100111001001;
    rom[55657] = 25'b0000000000011100111001100;
    rom[55658] = 25'b0000000000011100111010000;
    rom[55659] = 25'b0000000000011100111010100;
    rom[55660] = 25'b0000000000011100111011000;
    rom[55661] = 25'b0000000000011100111011011;
    rom[55662] = 25'b0000000000011100111011110;
    rom[55663] = 25'b0000000000011100111100010;
    rom[55664] = 25'b0000000000011100111100110;
    rom[55665] = 25'b0000000000011100111101001;
    rom[55666] = 25'b0000000000011100111101101;
    rom[55667] = 25'b0000000000011100111110000;
    rom[55668] = 25'b0000000000011100111110011;
    rom[55669] = 25'b0000000000011100111110111;
    rom[55670] = 25'b0000000000011100111111010;
    rom[55671] = 25'b0000000000011100111111110;
    rom[55672] = 25'b0000000000011101000000001;
    rom[55673] = 25'b0000000000011101000000101;
    rom[55674] = 25'b0000000000011101000001000;
    rom[55675] = 25'b0000000000011101000001010;
    rom[55676] = 25'b0000000000011101000001110;
    rom[55677] = 25'b0000000000011101000010001;
    rom[55678] = 25'b0000000000011101000010100;
    rom[55679] = 25'b0000000000011101000010111;
    rom[55680] = 25'b0000000000011101000011011;
    rom[55681] = 25'b0000000000011101000011110;
    rom[55682] = 25'b0000000000011101000100001;
    rom[55683] = 25'b0000000000011101000100100;
    rom[55684] = 25'b0000000000011101000100111;
    rom[55685] = 25'b0000000000011101000101010;
    rom[55686] = 25'b0000000000011101000101101;
    rom[55687] = 25'b0000000000011101000110000;
    rom[55688] = 25'b0000000000011101000110011;
    rom[55689] = 25'b0000000000011101000110110;
    rom[55690] = 25'b0000000000011101000111001;
    rom[55691] = 25'b0000000000011101000111100;
    rom[55692] = 25'b0000000000011101000111111;
    rom[55693] = 25'b0000000000011101001000001;
    rom[55694] = 25'b0000000000011101001000100;
    rom[55695] = 25'b0000000000011101001000111;
    rom[55696] = 25'b0000000000011101001001001;
    rom[55697] = 25'b0000000000011101001001100;
    rom[55698] = 25'b0000000000011101001001111;
    rom[55699] = 25'b0000000000011101001010001;
    rom[55700] = 25'b0000000000011101001010100;
    rom[55701] = 25'b0000000000011101001010111;
    rom[55702] = 25'b0000000000011101001011010;
    rom[55703] = 25'b0000000000011101001011100;
    rom[55704] = 25'b0000000000011101001011111;
    rom[55705] = 25'b0000000000011101001100001;
    rom[55706] = 25'b0000000000011101001100100;
    rom[55707] = 25'b0000000000011101001100110;
    rom[55708] = 25'b0000000000011101001101001;
    rom[55709] = 25'b0000000000011101001101100;
    rom[55710] = 25'b0000000000011101001101110;
    rom[55711] = 25'b0000000000011101001110000;
    rom[55712] = 25'b0000000000011101001110010;
    rom[55713] = 25'b0000000000011101001110101;
    rom[55714] = 25'b0000000000011101001111000;
    rom[55715] = 25'b0000000000011101001111010;
    rom[55716] = 25'b0000000000011101001111100;
    rom[55717] = 25'b0000000000011101001111110;
    rom[55718] = 25'b0000000000011101010000001;
    rom[55719] = 25'b0000000000011101010000011;
    rom[55720] = 25'b0000000000011101010000101;
    rom[55721] = 25'b0000000000011101010000111;
    rom[55722] = 25'b0000000000011101010001010;
    rom[55723] = 25'b0000000000011101010001100;
    rom[55724] = 25'b0000000000011101010001101;
    rom[55725] = 25'b0000000000011101010001111;
    rom[55726] = 25'b0000000000011101010010010;
    rom[55727] = 25'b0000000000011101010010100;
    rom[55728] = 25'b0000000000011101010010101;
    rom[55729] = 25'b0000000000011101010011000;
    rom[55730] = 25'b0000000000011101010011010;
    rom[55731] = 25'b0000000000011101010011011;
    rom[55732] = 25'b0000000000011101010011110;
    rom[55733] = 25'b0000000000011101010011111;
    rom[55734] = 25'b0000000000011101010100001;
    rom[55735] = 25'b0000000000011101010100011;
    rom[55736] = 25'b0000000000011101010100101;
    rom[55737] = 25'b0000000000011101010100111;
    rom[55738] = 25'b0000000000011101010101001;
    rom[55739] = 25'b0000000000011101010101010;
    rom[55740] = 25'b0000000000011101010101100;
    rom[55741] = 25'b0000000000011101010101110;
    rom[55742] = 25'b0000000000011101010110000;
    rom[55743] = 25'b0000000000011101010110001;
    rom[55744] = 25'b0000000000011101010110011;
    rom[55745] = 25'b0000000000011101010110101;
    rom[55746] = 25'b0000000000011101010110110;
    rom[55747] = 25'b0000000000011101010111000;
    rom[55748] = 25'b0000000000011101010111001;
    rom[55749] = 25'b0000000000011101010111011;
    rom[55750] = 25'b0000000000011101010111100;
    rom[55751] = 25'b0000000000011101010111110;
    rom[55752] = 25'b0000000000011101010111111;
    rom[55753] = 25'b0000000000011101011000001;
    rom[55754] = 25'b0000000000011101011000010;
    rom[55755] = 25'b0000000000011101011000100;
    rom[55756] = 25'b0000000000011101011000101;
    rom[55757] = 25'b0000000000011101011000110;
    rom[55758] = 25'b0000000000011101011001000;
    rom[55759] = 25'b0000000000011101011001001;
    rom[55760] = 25'b0000000000011101011001010;
    rom[55761] = 25'b0000000000011101011001011;
    rom[55762] = 25'b0000000000011101011001101;
    rom[55763] = 25'b0000000000011101011001110;
    rom[55764] = 25'b0000000000011101011001111;
    rom[55765] = 25'b0000000000011101011010000;
    rom[55766] = 25'b0000000000011101011010010;
    rom[55767] = 25'b0000000000011101011010011;
    rom[55768] = 25'b0000000000011101011010100;
    rom[55769] = 25'b0000000000011101011010101;
    rom[55770] = 25'b0000000000011101011010110;
    rom[55771] = 25'b0000000000011101011010111;
    rom[55772] = 25'b0000000000011101011011000;
    rom[55773] = 25'b0000000000011101011011001;
    rom[55774] = 25'b0000000000011101011011010;
    rom[55775] = 25'b0000000000011101011011011;
    rom[55776] = 25'b0000000000011101011011100;
    rom[55777] = 25'b0000000000011101011011101;
    rom[55778] = 25'b0000000000011101011011110;
    rom[55779] = 25'b0000000000011101011011111;
    rom[55780] = 25'b0000000000011101011011111;
    rom[55781] = 25'b0000000000011101011100000;
    rom[55782] = 25'b0000000000011101011100001;
    rom[55783] = 25'b0000000000011101011100010;
    rom[55784] = 25'b0000000000011101011100010;
    rom[55785] = 25'b0000000000011101011100011;
    rom[55786] = 25'b0000000000011101011100100;
    rom[55787] = 25'b0000000000011101011100101;
    rom[55788] = 25'b0000000000011101011100101;
    rom[55789] = 25'b0000000000011101011100110;
    rom[55790] = 25'b0000000000011101011100111;
    rom[55791] = 25'b0000000000011101011101000;
    rom[55792] = 25'b0000000000011101011101000;
    rom[55793] = 25'b0000000000011101011101000;
    rom[55794] = 25'b0000000000011101011101001;
    rom[55795] = 25'b0000000000011101011101001;
    rom[55796] = 25'b0000000000011101011101010;
    rom[55797] = 25'b0000000000011101011101011;
    rom[55798] = 25'b0000000000011101011101011;
    rom[55799] = 25'b0000000000011101011101011;
    rom[55800] = 25'b0000000000011101011101011;
    rom[55801] = 25'b0000000000011101011101100;
    rom[55802] = 25'b0000000000011101011101100;
    rom[55803] = 25'b0000000000011101011101101;
    rom[55804] = 25'b0000000000011101011101101;
    rom[55805] = 25'b0000000000011101011101110;
    rom[55806] = 25'b0000000000011101011101110;
    rom[55807] = 25'b0000000000011101011101110;
    rom[55808] = 25'b0000000000011101011101110;
    rom[55809] = 25'b0000000000011101011101110;
    rom[55810] = 25'b0000000000011101011101110;
    rom[55811] = 25'b0000000000011101011101110;
    rom[55812] = 25'b0000000000011101011101111;
    rom[55813] = 25'b0000000000011101011101111;
    rom[55814] = 25'b0000000000011101011101111;
    rom[55815] = 25'b0000000000011101011101111;
    rom[55816] = 25'b0000000000011101011101111;
    rom[55817] = 25'b0000000000011101011101111;
    rom[55818] = 25'b0000000000011101011101111;
    rom[55819] = 25'b0000000000011101011101111;
    rom[55820] = 25'b0000000000011101011101111;
    rom[55821] = 25'b0000000000011101011101111;
    rom[55822] = 25'b0000000000011101011101111;
    rom[55823] = 25'b0000000000011101011101111;
    rom[55824] = 25'b0000000000011101011101111;
    rom[55825] = 25'b0000000000011101011101110;
    rom[55826] = 25'b0000000000011101011101110;
    rom[55827] = 25'b0000000000011101011101110;
    rom[55828] = 25'b0000000000011101011101110;
    rom[55829] = 25'b0000000000011101011101110;
    rom[55830] = 25'b0000000000011101011101110;
    rom[55831] = 25'b0000000000011101011101110;
    rom[55832] = 25'b0000000000011101011101101;
    rom[55833] = 25'b0000000000011101011101101;
    rom[55834] = 25'b0000000000011101011101100;
    rom[55835] = 25'b0000000000011101011101100;
    rom[55836] = 25'b0000000000011101011101011;
    rom[55837] = 25'b0000000000011101011101011;
    rom[55838] = 25'b0000000000011101011101011;
    rom[55839] = 25'b0000000000011101011101011;
    rom[55840] = 25'b0000000000011101011101010;
    rom[55841] = 25'b0000000000011101011101001;
    rom[55842] = 25'b0000000000011101011101001;
    rom[55843] = 25'b0000000000011101011101000;
    rom[55844] = 25'b0000000000011101011101000;
    rom[55845] = 25'b0000000000011101011101000;
    rom[55846] = 25'b0000000000011101011100111;
    rom[55847] = 25'b0000000000011101011100110;
    rom[55848] = 25'b0000000000011101011100101;
    rom[55849] = 25'b0000000000011101011100101;
    rom[55850] = 25'b0000000000011101011100100;
    rom[55851] = 25'b0000000000011101011100011;
    rom[55852] = 25'b0000000000011101011100010;
    rom[55853] = 25'b0000000000011101011100010;
    rom[55854] = 25'b0000000000011101011100001;
    rom[55855] = 25'b0000000000011101011100000;
    rom[55856] = 25'b0000000000011101011011111;
    rom[55857] = 25'b0000000000011101011011111;
    rom[55858] = 25'b0000000000011101011011110;
    rom[55859] = 25'b0000000000011101011011101;
    rom[55860] = 25'b0000000000011101011011100;
    rom[55861] = 25'b0000000000011101011011011;
    rom[55862] = 25'b0000000000011101011011010;
    rom[55863] = 25'b0000000000011101011011001;
    rom[55864] = 25'b0000000000011101011011001;
    rom[55865] = 25'b0000000000011101011010111;
    rom[55866] = 25'b0000000000011101011010110;
    rom[55867] = 25'b0000000000011101011010101;
    rom[55868] = 25'b0000000000011101011010100;
    rom[55869] = 25'b0000000000011101011010011;
    rom[55870] = 25'b0000000000011101011010010;
    rom[55871] = 25'b0000000000011101011010001;
    rom[55872] = 25'b0000000000011101011010000;
    rom[55873] = 25'b0000000000011101011001111;
    rom[55874] = 25'b0000000000011101011001101;
    rom[55875] = 25'b0000000000011101011001100;
    rom[55876] = 25'b0000000000011101011001011;
    rom[55877] = 25'b0000000000011101011001010;
    rom[55878] = 25'b0000000000011101011001000;
    rom[55879] = 25'b0000000000011101011001000;
    rom[55880] = 25'b0000000000011101011000110;
    rom[55881] = 25'b0000000000011101011000101;
    rom[55882] = 25'b0000000000011101011000011;
    rom[55883] = 25'b0000000000011101011000010;
    rom[55884] = 25'b0000000000011101011000001;
    rom[55885] = 25'b0000000000011101010111111;
    rom[55886] = 25'b0000000000011101010111110;
    rom[55887] = 25'b0000000000011101010111100;
    rom[55888] = 25'b0000000000011101010111011;
    rom[55889] = 25'b0000000000011101010111001;
    rom[55890] = 25'b0000000000011101010111000;
    rom[55891] = 25'b0000000000011101010110110;
    rom[55892] = 25'b0000000000011101010110101;
    rom[55893] = 25'b0000000000011101010110011;
    rom[55894] = 25'b0000000000011101010110001;
    rom[55895] = 25'b0000000000011101010110000;
    rom[55896] = 25'b0000000000011101010101110;
    rom[55897] = 25'b0000000000011101010101101;
    rom[55898] = 25'b0000000000011101010101011;
    rom[55899] = 25'b0000000000011101010101001;
    rom[55900] = 25'b0000000000011101010100111;
    rom[55901] = 25'b0000000000011101010100110;
    rom[55902] = 25'b0000000000011101010100100;
    rom[55903] = 25'b0000000000011101010100010;
    rom[55904] = 25'b0000000000011101010100001;
    rom[55905] = 25'b0000000000011101010011110;
    rom[55906] = 25'b0000000000011101010011101;
    rom[55907] = 25'b0000000000011101010011011;
    rom[55908] = 25'b0000000000011101010011001;
    rom[55909] = 25'b0000000000011101010010111;
    rom[55910] = 25'b0000000000011101010010101;
    rom[55911] = 25'b0000000000011101010010011;
    rom[55912] = 25'b0000000000011101010010001;
    rom[55913] = 25'b0000000000011101010001111;
    rom[55914] = 25'b0000000000011101010001101;
    rom[55915] = 25'b0000000000011101010001011;
    rom[55916] = 25'b0000000000011101010001001;
    rom[55917] = 25'b0000000000011101010000111;
    rom[55918] = 25'b0000000000011101010000101;
    rom[55919] = 25'b0000000000011101010000011;
    rom[55920] = 25'b0000000000011101010000001;
    rom[55921] = 25'b0000000000011101001111110;
    rom[55922] = 25'b0000000000011101001111100;
    rom[55923] = 25'b0000000000011101001111011;
    rom[55924] = 25'b0000000000011101001111000;
    rom[55925] = 25'b0000000000011101001110110;
    rom[55926] = 25'b0000000000011101001110100;
    rom[55927] = 25'b0000000000011101001110010;
    rom[55928] = 25'b0000000000011101001101111;
    rom[55929] = 25'b0000000000011101001101100;
    rom[55930] = 25'b0000000000011101001101010;
    rom[55931] = 25'b0000000000011101001101000;
    rom[55932] = 25'b0000000000011101001100110;
    rom[55933] = 25'b0000000000011101001100011;
    rom[55934] = 25'b0000000000011101001100001;
    rom[55935] = 25'b0000000000011101001011110;
    rom[55936] = 25'b0000000000011101001011100;
    rom[55937] = 25'b0000000000011101001011010;
    rom[55938] = 25'b0000000000011101001010111;
    rom[55939] = 25'b0000000000011101001010100;
    rom[55940] = 25'b0000000000011101001010010;
    rom[55941] = 25'b0000000000011101001001111;
    rom[55942] = 25'b0000000000011101001001101;
    rom[55943] = 25'b0000000000011101001001010;
    rom[55944] = 25'b0000000000011101001001000;
    rom[55945] = 25'b0000000000011101001000101;
    rom[55946] = 25'b0000000000011101001000011;
    rom[55947] = 25'b0000000000011101001000000;
    rom[55948] = 25'b0000000000011101000111101;
    rom[55949] = 25'b0000000000011101000111010;
    rom[55950] = 25'b0000000000011101000110111;
    rom[55951] = 25'b0000000000011101000110101;
    rom[55952] = 25'b0000000000011101000110010;
    rom[55953] = 25'b0000000000011101000101111;
    rom[55954] = 25'b0000000000011101000101101;
    rom[55955] = 25'b0000000000011101000101010;
    rom[55956] = 25'b0000000000011101000100111;
    rom[55957] = 25'b0000000000011101000100100;
    rom[55958] = 25'b0000000000011101000100001;
    rom[55959] = 25'b0000000000011101000011110;
    rom[55960] = 25'b0000000000011101000011011;
    rom[55961] = 25'b0000000000011101000011001;
    rom[55962] = 25'b0000000000011101000010110;
    rom[55963] = 25'b0000000000011101000010011;
    rom[55964] = 25'b0000000000011101000010000;
    rom[55965] = 25'b0000000000011101000001101;
    rom[55966] = 25'b0000000000011101000001010;
    rom[55967] = 25'b0000000000011101000000110;
    rom[55968] = 25'b0000000000011101000000011;
    rom[55969] = 25'b0000000000011101000000000;
    rom[55970] = 25'b0000000000011100111111101;
    rom[55971] = 25'b0000000000011100111111010;
    rom[55972] = 25'b0000000000011100111110111;
    rom[55973] = 25'b0000000000011100111110011;
    rom[55974] = 25'b0000000000011100111110000;
    rom[55975] = 25'b0000000000011100111101101;
    rom[55976] = 25'b0000000000011100111101010;
    rom[55977] = 25'b0000000000011100111100111;
    rom[55978] = 25'b0000000000011100111100100;
    rom[55979] = 25'b0000000000011100111100000;
    rom[55980] = 25'b0000000000011100111011101;
    rom[55981] = 25'b0000000000011100111011001;
    rom[55982] = 25'b0000000000011100111010110;
    rom[55983] = 25'b0000000000011100111010011;
    rom[55984] = 25'b0000000000011100111001111;
    rom[55985] = 25'b0000000000011100111001100;
    rom[55986] = 25'b0000000000011100111001001;
    rom[55987] = 25'b0000000000011100111000101;
    rom[55988] = 25'b0000000000011100111000010;
    rom[55989] = 25'b0000000000011100110111110;
    rom[55990] = 25'b0000000000011100110111011;
    rom[55991] = 25'b0000000000011100110111000;
    rom[55992] = 25'b0000000000011100110110100;
    rom[55993] = 25'b0000000000011100110110000;
    rom[55994] = 25'b0000000000011100110101100;
    rom[55995] = 25'b0000000000011100110101001;
    rom[55996] = 25'b0000000000011100110100110;
    rom[55997] = 25'b0000000000011100110100010;
    rom[55998] = 25'b0000000000011100110011110;
    rom[55999] = 25'b0000000000011100110011010;
    rom[56000] = 25'b0000000000011100110010111;
    rom[56001] = 25'b0000000000011100110010011;
    rom[56002] = 25'b0000000000011100110001111;
    rom[56003] = 25'b0000000000011100110001011;
    rom[56004] = 25'b0000000000011100110001000;
    rom[56005] = 25'b0000000000011100110000100;
    rom[56006] = 25'b0000000000011100110000000;
    rom[56007] = 25'b0000000000011100101111101;
    rom[56008] = 25'b0000000000011100101111001;
    rom[56009] = 25'b0000000000011100101110101;
    rom[56010] = 25'b0000000000011100101110001;
    rom[56011] = 25'b0000000000011100101101101;
    rom[56012] = 25'b0000000000011100101101001;
    rom[56013] = 25'b0000000000011100101100101;
    rom[56014] = 25'b0000000000011100101100010;
    rom[56015] = 25'b0000000000011100101011101;
    rom[56016] = 25'b0000000000011100101011001;
    rom[56017] = 25'b0000000000011100101010110;
    rom[56018] = 25'b0000000000011100101010001;
    rom[56019] = 25'b0000000000011100101001101;
    rom[56020] = 25'b0000000000011100101001001;
    rom[56021] = 25'b0000000000011100101000101;
    rom[56022] = 25'b0000000000011100101000001;
    rom[56023] = 25'b0000000000011100100111101;
    rom[56024] = 25'b0000000000011100100111001;
    rom[56025] = 25'b0000000000011100100110101;
    rom[56026] = 25'b0000000000011100100110000;
    rom[56027] = 25'b0000000000011100100101101;
    rom[56028] = 25'b0000000000011100100101000;
    rom[56029] = 25'b0000000000011100100100100;
    rom[56030] = 25'b0000000000011100100100000;
    rom[56031] = 25'b0000000000011100100011011;
    rom[56032] = 25'b0000000000011100100010111;
    rom[56033] = 25'b0000000000011100100010011;
    rom[56034] = 25'b0000000000011100100001111;
    rom[56035] = 25'b0000000000011100100001010;
    rom[56036] = 25'b0000000000011100100000110;
    rom[56037] = 25'b0000000000011100100000001;
    rom[56038] = 25'b0000000000011100011111110;
    rom[56039] = 25'b0000000000011100011111001;
    rom[56040] = 25'b0000000000011100011110101;
    rom[56041] = 25'b0000000000011100011110000;
    rom[56042] = 25'b0000000000011100011101100;
    rom[56043] = 25'b0000000000011100011100111;
    rom[56044] = 25'b0000000000011100011100011;
    rom[56045] = 25'b0000000000011100011011110;
    rom[56046] = 25'b0000000000011100011011010;
    rom[56047] = 25'b0000000000011100011010101;
    rom[56048] = 25'b0000000000011100011010001;
    rom[56049] = 25'b0000000000011100011001011;
    rom[56050] = 25'b0000000000011100011000111;
    rom[56051] = 25'b0000000000011100011000011;
    rom[56052] = 25'b0000000000011100010111110;
    rom[56053] = 25'b0000000000011100010111010;
    rom[56054] = 25'b0000000000011100010110100;
    rom[56055] = 25'b0000000000011100010110000;
    rom[56056] = 25'b0000000000011100010101011;
    rom[56057] = 25'b0000000000011100010100111;
    rom[56058] = 25'b0000000000011100010100010;
    rom[56059] = 25'b0000000000011100010011101;
    rom[56060] = 25'b0000000000011100010011000;
    rom[56061] = 25'b0000000000011100010010011;
    rom[56062] = 25'b0000000000011100010001111;
    rom[56063] = 25'b0000000000011100010001010;
    rom[56064] = 25'b0000000000011100010000101;
    rom[56065] = 25'b0000000000011100010000000;
    rom[56066] = 25'b0000000000011100001111100;
    rom[56067] = 25'b0000000000011100001110110;
    rom[56068] = 25'b0000000000011100001110010;
    rom[56069] = 25'b0000000000011100001101101;
    rom[56070] = 25'b0000000000011100001100111;
    rom[56071] = 25'b0000000000011100001100011;
    rom[56072] = 25'b0000000000011100001011110;
    rom[56073] = 25'b0000000000011100001011000;
    rom[56074] = 25'b0000000000011100001010100;
    rom[56075] = 25'b0000000000011100001001111;
    rom[56076] = 25'b0000000000011100001001001;
    rom[56077] = 25'b0000000000011100001000100;
    rom[56078] = 25'b0000000000011100000111111;
    rom[56079] = 25'b0000000000011100000111011;
    rom[56080] = 25'b0000000000011100000110101;
    rom[56081] = 25'b0000000000011100000110000;
    rom[56082] = 25'b0000000000011100000101011;
    rom[56083] = 25'b0000000000011100000100110;
    rom[56084] = 25'b0000000000011100000100000;
    rom[56085] = 25'b0000000000011100000011011;
    rom[56086] = 25'b0000000000011100000010110;
    rom[56087] = 25'b0000000000011100000010001;
    rom[56088] = 25'b0000000000011100000001011;
    rom[56089] = 25'b0000000000011100000000110;
    rom[56090] = 25'b0000000000011100000000001;
    rom[56091] = 25'b0000000000011011111111100;
    rom[56092] = 25'b0000000000011011111110111;
    rom[56093] = 25'b0000000000011011111110001;
    rom[56094] = 25'b0000000000011011111101011;
    rom[56095] = 25'b0000000000011011111100110;
    rom[56096] = 25'b0000000000011011111100001;
    rom[56097] = 25'b0000000000011011111011100;
    rom[56098] = 25'b0000000000011011111010110;
    rom[56099] = 25'b0000000000011011111010000;
    rom[56100] = 25'b0000000000011011111001011;
    rom[56101] = 25'b0000000000011011111000110;
    rom[56102] = 25'b0000000000011011111000000;
    rom[56103] = 25'b0000000000011011110111011;
    rom[56104] = 25'b0000000000011011110110101;
    rom[56105] = 25'b0000000000011011110110000;
    rom[56106] = 25'b0000000000011011110101010;
    rom[56107] = 25'b0000000000011011110100100;
    rom[56108] = 25'b0000000000011011110011111;
    rom[56109] = 25'b0000000000011011110011001;
    rom[56110] = 25'b0000000000011011110010011;
    rom[56111] = 25'b0000000000011011110001110;
    rom[56112] = 25'b0000000000011011110001000;
    rom[56113] = 25'b0000000000011011110000011;
    rom[56114] = 25'b0000000000011011101111101;
    rom[56115] = 25'b0000000000011011101110111;
    rom[56116] = 25'b0000000000011011101110010;
    rom[56117] = 25'b0000000000011011101101100;
    rom[56118] = 25'b0000000000011011101100110;
    rom[56119] = 25'b0000000000011011101100000;
    rom[56120] = 25'b0000000000011011101011010;
    rom[56121] = 25'b0000000000011011101010100;
    rom[56122] = 25'b0000000000011011101001110;
    rom[56123] = 25'b0000000000011011101001001;
    rom[56124] = 25'b0000000000011011101000011;
    rom[56125] = 25'b0000000000011011100111101;
    rom[56126] = 25'b0000000000011011100110111;
    rom[56127] = 25'b0000000000011011100110001;
    rom[56128] = 25'b0000000000011011100101011;
    rom[56129] = 25'b0000000000011011100100101;
    rom[56130] = 25'b0000000000011011100011111;
    rom[56131] = 25'b0000000000011011100011001;
    rom[56132] = 25'b0000000000011011100010011;
    rom[56133] = 25'b0000000000011011100001101;
    rom[56134] = 25'b0000000000011011100000111;
    rom[56135] = 25'b0000000000011011100000010;
    rom[56136] = 25'b0000000000011011011111100;
    rom[56137] = 25'b0000000000011011011110110;
    rom[56138] = 25'b0000000000011011011110000;
    rom[56139] = 25'b0000000000011011011101001;
    rom[56140] = 25'b0000000000011011011100011;
    rom[56141] = 25'b0000000000011011011011101;
    rom[56142] = 25'b0000000000011011011010111;
    rom[56143] = 25'b0000000000011011011010000;
    rom[56144] = 25'b0000000000011011011001010;
    rom[56145] = 25'b0000000000011011011000100;
    rom[56146] = 25'b0000000000011011010111110;
    rom[56147] = 25'b0000000000011011010111000;
    rom[56148] = 25'b0000000000011011010110010;
    rom[56149] = 25'b0000000000011011010101011;
    rom[56150] = 25'b0000000000011011010100101;
    rom[56151] = 25'b0000000000011011010011111;
    rom[56152] = 25'b0000000000011011010011000;
    rom[56153] = 25'b0000000000011011010010010;
    rom[56154] = 25'b0000000000011011010001011;
    rom[56155] = 25'b0000000000011011010000101;
    rom[56156] = 25'b0000000000011011001111111;
    rom[56157] = 25'b0000000000011011001111001;
    rom[56158] = 25'b0000000000011011001110010;
    rom[56159] = 25'b0000000000011011001101011;
    rom[56160] = 25'b0000000000011011001100101;
    rom[56161] = 25'b0000000000011011001011111;
    rom[56162] = 25'b0000000000011011001011001;
    rom[56163] = 25'b0000000000011011001010010;
    rom[56164] = 25'b0000000000011011001001011;
    rom[56165] = 25'b0000000000011011001000101;
    rom[56166] = 25'b0000000000011011000111111;
    rom[56167] = 25'b0000000000011011000111000;
    rom[56168] = 25'b0000000000011011000110001;
    rom[56169] = 25'b0000000000011011000101010;
    rom[56170] = 25'b0000000000011011000100100;
    rom[56171] = 25'b0000000000011011000011110;
    rom[56172] = 25'b0000000000011011000010111;
    rom[56173] = 25'b0000000000011011000010000;
    rom[56174] = 25'b0000000000011011000001001;
    rom[56175] = 25'b0000000000011011000000011;
    rom[56176] = 25'b0000000000011010111111100;
    rom[56177] = 25'b0000000000011010111110101;
    rom[56178] = 25'b0000000000011010111101111;
    rom[56179] = 25'b0000000000011010111101000;
    rom[56180] = 25'b0000000000011010111100001;
    rom[56181] = 25'b0000000000011010111011010;
    rom[56182] = 25'b0000000000011010111010100;
    rom[56183] = 25'b0000000000011010111001101;
    rom[56184] = 25'b0000000000011010111000110;
    rom[56185] = 25'b0000000000011010111000000;
    rom[56186] = 25'b0000000000011010110111000;
    rom[56187] = 25'b0000000000011010110110001;
    rom[56188] = 25'b0000000000011010110101011;
    rom[56189] = 25'b0000000000011010110100100;
    rom[56190] = 25'b0000000000011010110011101;
    rom[56191] = 25'b0000000000011010110010110;
    rom[56192] = 25'b0000000000011010110001111;
    rom[56193] = 25'b0000000000011010110001000;
    rom[56194] = 25'b0000000000011010110000010;
    rom[56195] = 25'b0000000000011010101111010;
    rom[56196] = 25'b0000000000011010101110011;
    rom[56197] = 25'b0000000000011010101101100;
    rom[56198] = 25'b0000000000011010101100101;
    rom[56199] = 25'b0000000000011010101011110;
    rom[56200] = 25'b0000000000011010101010111;
    rom[56201] = 25'b0000000000011010101010000;
    rom[56202] = 25'b0000000000011010101001001;
    rom[56203] = 25'b0000000000011010101000010;
    rom[56204] = 25'b0000000000011010100111011;
    rom[56205] = 25'b0000000000011010100110100;
    rom[56206] = 25'b0000000000011010100101100;
    rom[56207] = 25'b0000000000011010100100110;
    rom[56208] = 25'b0000000000011010100011110;
    rom[56209] = 25'b0000000000011010100010111;
    rom[56210] = 25'b0000000000011010100010000;
    rom[56211] = 25'b0000000000011010100001000;
    rom[56212] = 25'b0000000000011010100000001;
    rom[56213] = 25'b0000000000011010011111010;
    rom[56214] = 25'b0000000000011010011110011;
    rom[56215] = 25'b0000000000011010011101011;
    rom[56216] = 25'b0000000000011010011100101;
    rom[56217] = 25'b0000000000011010011011101;
    rom[56218] = 25'b0000000000011010011010110;
    rom[56219] = 25'b0000000000011010011001110;
    rom[56220] = 25'b0000000000011010011000111;
    rom[56221] = 25'b0000000000011010010111111;
    rom[56222] = 25'b0000000000011010010111001;
    rom[56223] = 25'b0000000000011010010110001;
    rom[56224] = 25'b0000000000011010010101010;
    rom[56225] = 25'b0000000000011010010100010;
    rom[56226] = 25'b0000000000011010010011011;
    rom[56227] = 25'b0000000000011010010010011;
    rom[56228] = 25'b0000000000011010010001100;
    rom[56229] = 25'b0000000000011010010000100;
    rom[56230] = 25'b0000000000011010001111101;
    rom[56231] = 25'b0000000000011010001110101;
    rom[56232] = 25'b0000000000011010001101110;
    rom[56233] = 25'b0000000000011010001100110;
    rom[56234] = 25'b0000000000011010001011111;
    rom[56235] = 25'b0000000000011010001010111;
    rom[56236] = 25'b0000000000011010001001111;
    rom[56237] = 25'b0000000000011010001001000;
    rom[56238] = 25'b0000000000011010001000000;
    rom[56239] = 25'b0000000000011010000111001;
    rom[56240] = 25'b0000000000011010000110001;
    rom[56241] = 25'b0000000000011010000101010;
    rom[56242] = 25'b0000000000011010000100010;
    rom[56243] = 25'b0000000000011010000011010;
    rom[56244] = 25'b0000000000011010000010011;
    rom[56245] = 25'b0000000000011010000001010;
    rom[56246] = 25'b0000000000011010000000011;
    rom[56247] = 25'b0000000000011001111111100;
    rom[56248] = 25'b0000000000011001111110011;
    rom[56249] = 25'b0000000000011001111101100;
    rom[56250] = 25'b0000000000011001111100100;
    rom[56251] = 25'b0000000000011001111011100;
    rom[56252] = 25'b0000000000011001111010101;
    rom[56253] = 25'b0000000000011001111001100;
    rom[56254] = 25'b0000000000011001111000101;
    rom[56255] = 25'b0000000000011001110111101;
    rom[56256] = 25'b0000000000011001110110101;
    rom[56257] = 25'b0000000000011001110101101;
    rom[56258] = 25'b0000000000011001110100110;
    rom[56259] = 25'b0000000000011001110011101;
    rom[56260] = 25'b0000000000011001110010110;
    rom[56261] = 25'b0000000000011001110001110;
    rom[56262] = 25'b0000000000011001110000101;
    rom[56263] = 25'b0000000000011001101111110;
    rom[56264] = 25'b0000000000011001101110110;
    rom[56265] = 25'b0000000000011001101101110;
    rom[56266] = 25'b0000000000011001101100110;
    rom[56267] = 25'b0000000000011001101011110;
    rom[56268] = 25'b0000000000011001101010110;
    rom[56269] = 25'b0000000000011001101001110;
    rom[56270] = 25'b0000000000011001101000110;
    rom[56271] = 25'b0000000000011001100111110;
    rom[56272] = 25'b0000000000011001100110110;
    rom[56273] = 25'b0000000000011001100101101;
    rom[56274] = 25'b0000000000011001100100110;
    rom[56275] = 25'b0000000000011001100011110;
    rom[56276] = 25'b0000000000011001100010101;
    rom[56277] = 25'b0000000000011001100001101;
    rom[56278] = 25'b0000000000011001100000101;
    rom[56279] = 25'b0000000000011001011111101;
    rom[56280] = 25'b0000000000011001011110101;
    rom[56281] = 25'b0000000000011001011101100;
    rom[56282] = 25'b0000000000011001011100100;
    rom[56283] = 25'b0000000000011001011011100;
    rom[56284] = 25'b0000000000011001011010100;
    rom[56285] = 25'b0000000000011001011001011;
    rom[56286] = 25'b0000000000011001011000011;
    rom[56287] = 25'b0000000000011001010111011;
    rom[56288] = 25'b0000000000011001010110011;
    rom[56289] = 25'b0000000000011001010101011;
    rom[56290] = 25'b0000000000011001010100010;
    rom[56291] = 25'b0000000000011001010011010;
    rom[56292] = 25'b0000000000011001010010010;
    rom[56293] = 25'b0000000000011001010001001;
    rom[56294] = 25'b0000000000011001010000001;
    rom[56295] = 25'b0000000000011001001111001;
    rom[56296] = 25'b0000000000011001001110000;
    rom[56297] = 25'b0000000000011001001101000;
    rom[56298] = 25'b0000000000011001001011111;
    rom[56299] = 25'b0000000000011001001010111;
    rom[56300] = 25'b0000000000011001001001111;
    rom[56301] = 25'b0000000000011001001000110;
    rom[56302] = 25'b0000000000011001000111110;
    rom[56303] = 25'b0000000000011001000110101;
    rom[56304] = 25'b0000000000011001000101101;
    rom[56305] = 25'b0000000000011001000100100;
    rom[56306] = 25'b0000000000011001000011100;
    rom[56307] = 25'b0000000000011001000010011;
    rom[56308] = 25'b0000000000011001000001011;
    rom[56309] = 25'b0000000000011001000000010;
    rom[56310] = 25'b0000000000011000111111010;
    rom[56311] = 25'b0000000000011000111110001;
    rom[56312] = 25'b0000000000011000111101000;
    rom[56313] = 25'b0000000000011000111100000;
    rom[56314] = 25'b0000000000011000111010111;
    rom[56315] = 25'b0000000000011000111001111;
    rom[56316] = 25'b0000000000011000111000110;
    rom[56317] = 25'b0000000000011000110111101;
    rom[56318] = 25'b0000000000011000110110101;
    rom[56319] = 25'b0000000000011000110101100;
    rom[56320] = 25'b0000000000011000110100100;
    rom[56321] = 25'b0000000000011000110011011;
    rom[56322] = 25'b0000000000011000110010010;
    rom[56323] = 25'b0000000000011000110001001;
    rom[56324] = 25'b0000000000011000110000000;
    rom[56325] = 25'b0000000000011000101111000;
    rom[56326] = 25'b0000000000011000101101111;
    rom[56327] = 25'b0000000000011000101100110;
    rom[56328] = 25'b0000000000011000101011101;
    rom[56329] = 25'b0000000000011000101010100;
    rom[56330] = 25'b0000000000011000101001011;
    rom[56331] = 25'b0000000000011000101000011;
    rom[56332] = 25'b0000000000011000100111010;
    rom[56333] = 25'b0000000000011000100110001;
    rom[56334] = 25'b0000000000011000100101000;
    rom[56335] = 25'b0000000000011000100011111;
    rom[56336] = 25'b0000000000011000100010110;
    rom[56337] = 25'b0000000000011000100001101;
    rom[56338] = 25'b0000000000011000100000101;
    rom[56339] = 25'b0000000000011000011111100;
    rom[56340] = 25'b0000000000011000011110011;
    rom[56341] = 25'b0000000000011000011101010;
    rom[56342] = 25'b0000000000011000011100001;
    rom[56343] = 25'b0000000000011000011011000;
    rom[56344] = 25'b0000000000011000011001111;
    rom[56345] = 25'b0000000000011000011000110;
    rom[56346] = 25'b0000000000011000010111101;
    rom[56347] = 25'b0000000000011000010110101;
    rom[56348] = 25'b0000000000011000010101100;
    rom[56349] = 25'b0000000000011000010100010;
    rom[56350] = 25'b0000000000011000010011001;
    rom[56351] = 25'b0000000000011000010010000;
    rom[56352] = 25'b0000000000011000010000111;
    rom[56353] = 25'b0000000000011000001111110;
    rom[56354] = 25'b0000000000011000001110101;
    rom[56355] = 25'b0000000000011000001101100;
    rom[56356] = 25'b0000000000011000001100010;
    rom[56357] = 25'b0000000000011000001011001;
    rom[56358] = 25'b0000000000011000001010000;
    rom[56359] = 25'b0000000000011000001000111;
    rom[56360] = 25'b0000000000011000000111110;
    rom[56361] = 25'b0000000000011000000110101;
    rom[56362] = 25'b0000000000011000000101100;
    rom[56363] = 25'b0000000000011000000100011;
    rom[56364] = 25'b0000000000011000000011001;
    rom[56365] = 25'b0000000000011000000010000;
    rom[56366] = 25'b0000000000011000000000110;
    rom[56367] = 25'b0000000000010111111111101;
    rom[56368] = 25'b0000000000010111111110101;
    rom[56369] = 25'b0000000000010111111101011;
    rom[56370] = 25'b0000000000010111111100010;
    rom[56371] = 25'b0000000000010111111011000;
    rom[56372] = 25'b0000000000010111111001111;
    rom[56373] = 25'b0000000000010111111000110;
    rom[56374] = 25'b0000000000010111110111100;
    rom[56375] = 25'b0000000000010111110110100;
    rom[56376] = 25'b0000000000010111110101010;
    rom[56377] = 25'b0000000000010111110100001;
    rom[56378] = 25'b0000000000010111110010111;
    rom[56379] = 25'b0000000000010111110001110;
    rom[56380] = 25'b0000000000010111110000100;
    rom[56381] = 25'b0000000000010111101111011;
    rom[56382] = 25'b0000000000010111101110010;
    rom[56383] = 25'b0000000000010111101101000;
    rom[56384] = 25'b0000000000010111101011111;
    rom[56385] = 25'b0000000000010111101010101;
    rom[56386] = 25'b0000000000010111101001100;
    rom[56387] = 25'b0000000000010111101000011;
    rom[56388] = 25'b0000000000010111100111001;
    rom[56389] = 25'b0000000000010111100101111;
    rom[56390] = 25'b0000000000010111100100110;
    rom[56391] = 25'b0000000000010111100011101;
    rom[56392] = 25'b0000000000010111100010011;
    rom[56393] = 25'b0000000000010111100001001;
    rom[56394] = 25'b0000000000010111100000000;
    rom[56395] = 25'b0000000000010111011110111;
    rom[56396] = 25'b0000000000010111011101101;
    rom[56397] = 25'b0000000000010111011100011;
    rom[56398] = 25'b0000000000010111011011001;
    rom[56399] = 25'b0000000000010111011010000;
    rom[56400] = 25'b0000000000010111011000111;
    rom[56401] = 25'b0000000000010111010111101;
    rom[56402] = 25'b0000000000010111010110011;
    rom[56403] = 25'b0000000000010111010101010;
    rom[56404] = 25'b0000000000010111010100000;
    rom[56405] = 25'b0000000000010111010010110;
    rom[56406] = 25'b0000000000010111010001100;
    rom[56407] = 25'b0000000000010111010000011;
    rom[56408] = 25'b0000000000010111001111001;
    rom[56409] = 25'b0000000000010111001101111;
    rom[56410] = 25'b0000000000010111001100110;
    rom[56411] = 25'b0000000000010111001011100;
    rom[56412] = 25'b0000000000010111001010010;
    rom[56413] = 25'b0000000000010111001001000;
    rom[56414] = 25'b0000000000010111000111111;
    rom[56415] = 25'b0000000000010111000110101;
    rom[56416] = 25'b0000000000010111000101011;
    rom[56417] = 25'b0000000000010111000100010;
    rom[56418] = 25'b0000000000010111000011000;
    rom[56419] = 25'b0000000000010111000001110;
    rom[56420] = 25'b0000000000010111000000100;
    rom[56421] = 25'b0000000000010110111111010;
    rom[56422] = 25'b0000000000010110111110000;
    rom[56423] = 25'b0000000000010110111100111;
    rom[56424] = 25'b0000000000010110111011101;
    rom[56425] = 25'b0000000000010110111010011;
    rom[56426] = 25'b0000000000010110111001001;
    rom[56427] = 25'b0000000000010110110111111;
    rom[56428] = 25'b0000000000010110110110101;
    rom[56429] = 25'b0000000000010110110101100;
    rom[56430] = 25'b0000000000010110110100001;
    rom[56431] = 25'b0000000000010110110010111;
    rom[56432] = 25'b0000000000010110110001110;
    rom[56433] = 25'b0000000000010110110000100;
    rom[56434] = 25'b0000000000010110101111001;
    rom[56435] = 25'b0000000000010110101110000;
    rom[56436] = 25'b0000000000010110101100110;
    rom[56437] = 25'b0000000000010110101011100;
    rom[56438] = 25'b0000000000010110101010010;
    rom[56439] = 25'b0000000000010110101000111;
    rom[56440] = 25'b0000000000010110100111110;
    rom[56441] = 25'b0000000000010110100110100;
    rom[56442] = 25'b0000000000010110100101010;
    rom[56443] = 25'b0000000000010110100100000;
    rom[56444] = 25'b0000000000010110100010101;
    rom[56445] = 25'b0000000000010110100001100;
    rom[56446] = 25'b0000000000010110100000001;
    rom[56447] = 25'b0000000000010110011111000;
    rom[56448] = 25'b0000000000010110011101101;
    rom[56449] = 25'b0000000000010110011100011;
    rom[56450] = 25'b0000000000010110011011001;
    rom[56451] = 25'b0000000000010110011001111;
    rom[56452] = 25'b0000000000010110011000101;
    rom[56453] = 25'b0000000000010110010111011;
    rom[56454] = 25'b0000000000010110010110001;
    rom[56455] = 25'b0000000000010110010100110;
    rom[56456] = 25'b0000000000010110010011100;
    rom[56457] = 25'b0000000000010110010010010;
    rom[56458] = 25'b0000000000010110010000111;
    rom[56459] = 25'b0000000000010110001111110;
    rom[56460] = 25'b0000000000010110001110011;
    rom[56461] = 25'b0000000000010110001101010;
    rom[56462] = 25'b0000000000010110001011111;
    rom[56463] = 25'b0000000000010110001010101;
    rom[56464] = 25'b0000000000010110001001010;
    rom[56465] = 25'b0000000000010110001000000;
    rom[56466] = 25'b0000000000010110000110110;
    rom[56467] = 25'b0000000000010110000101100;
    rom[56468] = 25'b0000000000010110000100001;
    rom[56469] = 25'b0000000000010110000010111;
    rom[56470] = 25'b0000000000010110000001101;
    rom[56471] = 25'b0000000000010110000000010;
    rom[56472] = 25'b0000000000010101111111000;
    rom[56473] = 25'b0000000000010101111101110;
    rom[56474] = 25'b0000000000010101111100100;
    rom[56475] = 25'b0000000000010101111011001;
    rom[56476] = 25'b0000000000010101111001111;
    rom[56477] = 25'b0000000000010101111000100;
    rom[56478] = 25'b0000000000010101110111010;
    rom[56479] = 25'b0000000000010101110110000;
    rom[56480] = 25'b0000000000010101110100101;
    rom[56481] = 25'b0000000000010101110011011;
    rom[56482] = 25'b0000000000010101110010001;
    rom[56483] = 25'b0000000000010101110000110;
    rom[56484] = 25'b0000000000010101101111100;
    rom[56485] = 25'b0000000000010101101110010;
    rom[56486] = 25'b0000000000010101101100111;
    rom[56487] = 25'b0000000000010101101011101;
    rom[56488] = 25'b0000000000010101101010010;
    rom[56489] = 25'b0000000000010101101001000;
    rom[56490] = 25'b0000000000010101100111101;
    rom[56491] = 25'b0000000000010101100110011;
    rom[56492] = 25'b0000000000010101100101000;
    rom[56493] = 25'b0000000000010101100011110;
    rom[56494] = 25'b0000000000010101100010011;
    rom[56495] = 25'b0000000000010101100001000;
    rom[56496] = 25'b0000000000010101011111110;
    rom[56497] = 25'b0000000000010101011110011;
    rom[56498] = 25'b0000000000010101011101001;
    rom[56499] = 25'b0000000000010101011011110;
    rom[56500] = 25'b0000000000010101011010100;
    rom[56501] = 25'b0000000000010101011001001;
    rom[56502] = 25'b0000000000010101010111110;
    rom[56503] = 25'b0000000000010101010110100;
    rom[56504] = 25'b0000000000010101010101001;
    rom[56505] = 25'b0000000000010101010011111;
    rom[56506] = 25'b0000000000010101010010100;
    rom[56507] = 25'b0000000000010101010001010;
    rom[56508] = 25'b0000000000010101001111111;
    rom[56509] = 25'b0000000000010101001110100;
    rom[56510] = 25'b0000000000010101001101010;
    rom[56511] = 25'b0000000000010101001011111;
    rom[56512] = 25'b0000000000010101001010100;
    rom[56513] = 25'b0000000000010101001001010;
    rom[56514] = 25'b0000000000010101000111111;
    rom[56515] = 25'b0000000000010101000110100;
    rom[56516] = 25'b0000000000010101000101010;
    rom[56517] = 25'b0000000000010101000011111;
    rom[56518] = 25'b0000000000010101000010100;
    rom[56519] = 25'b0000000000010101000001001;
    rom[56520] = 25'b0000000000010100111111111;
    rom[56521] = 25'b0000000000010100111110100;
    rom[56522] = 25'b0000000000010100111101001;
    rom[56523] = 25'b0000000000010100111011111;
    rom[56524] = 25'b0000000000010100111010100;
    rom[56525] = 25'b0000000000010100111001001;
    rom[56526] = 25'b0000000000010100110111110;
    rom[56527] = 25'b0000000000010100110110100;
    rom[56528] = 25'b0000000000010100110101000;
    rom[56529] = 25'b0000000000010100110011110;
    rom[56530] = 25'b0000000000010100110010011;
    rom[56531] = 25'b0000000000010100110001000;
    rom[56532] = 25'b0000000000010100101111101;
    rom[56533] = 25'b0000000000010100101110011;
    rom[56534] = 25'b0000000000010100101100111;
    rom[56535] = 25'b0000000000010100101011101;
    rom[56536] = 25'b0000000000010100101010010;
    rom[56537] = 25'b0000000000010100101000111;
    rom[56538] = 25'b0000000000010100100111100;
    rom[56539] = 25'b0000000000010100100110010;
    rom[56540] = 25'b0000000000010100100100110;
    rom[56541] = 25'b0000000000010100100011100;
    rom[56542] = 25'b0000000000010100100010001;
    rom[56543] = 25'b0000000000010100100000101;
    rom[56544] = 25'b0000000000010100011111011;
    rom[56545] = 25'b0000000000010100011110000;
    rom[56546] = 25'b0000000000010100011100101;
    rom[56547] = 25'b0000000000010100011011010;
    rom[56548] = 25'b0000000000010100011001111;
    rom[56549] = 25'b0000000000010100011000100;
    rom[56550] = 25'b0000000000010100010111001;
    rom[56551] = 25'b0000000000010100010101110;
    rom[56552] = 25'b0000000000010100010100100;
    rom[56553] = 25'b0000000000010100010011000;
    rom[56554] = 25'b0000000000010100010001101;
    rom[56555] = 25'b0000000000010100010000010;
    rom[56556] = 25'b0000000000010100001110111;
    rom[56557] = 25'b0000000000010100001101100;
    rom[56558] = 25'b0000000000010100001100001;
    rom[56559] = 25'b0000000000010100001010110;
    rom[56560] = 25'b0000000000010100001001011;
    rom[56561] = 25'b0000000000010100001000000;
    rom[56562] = 25'b0000000000010100000110101;
    rom[56563] = 25'b0000000000010100000101010;
    rom[56564] = 25'b0000000000010100000011111;
    rom[56565] = 25'b0000000000010100000010100;
    rom[56566] = 25'b0000000000010100000001001;
    rom[56567] = 25'b0000000000010011111111110;
    rom[56568] = 25'b0000000000010011111110010;
    rom[56569] = 25'b0000000000010011111100111;
    rom[56570] = 25'b0000000000010011111011100;
    rom[56571] = 25'b0000000000010011111010001;
    rom[56572] = 25'b0000000000010011111000110;
    rom[56573] = 25'b0000000000010011110111011;
    rom[56574] = 25'b0000000000010011110110000;
    rom[56575] = 25'b0000000000010011110100101;
    rom[56576] = 25'b0000000000010011110011010;
    rom[56577] = 25'b0000000000010011110001110;
    rom[56578] = 25'b0000000000010011110000011;
    rom[56579] = 25'b0000000000010011101111000;
    rom[56580] = 25'b0000000000010011101101101;
    rom[56581] = 25'b0000000000010011101100010;
    rom[56582] = 25'b0000000000010011101010110;
    rom[56583] = 25'b0000000000010011101001011;
    rom[56584] = 25'b0000000000010011101000000;
    rom[56585] = 25'b0000000000010011100110101;
    rom[56586] = 25'b0000000000010011100101010;
    rom[56587] = 25'b0000000000010011100011110;
    rom[56588] = 25'b0000000000010011100010011;
    rom[56589] = 25'b0000000000010011100001000;
    rom[56590] = 25'b0000000000010011011111101;
    rom[56591] = 25'b0000000000010011011110001;
    rom[56592] = 25'b0000000000010011011100110;
    rom[56593] = 25'b0000000000010011011011011;
    rom[56594] = 25'b0000000000010011011010000;
    rom[56595] = 25'b0000000000010011011000101;
    rom[56596] = 25'b0000000000010011010111001;
    rom[56597] = 25'b0000000000010011010101110;
    rom[56598] = 25'b0000000000010011010100010;
    rom[56599] = 25'b0000000000010011010010111;
    rom[56600] = 25'b0000000000010011010001100;
    rom[56601] = 25'b0000000000010011010000001;
    rom[56602] = 25'b0000000000010011001110101;
    rom[56603] = 25'b0000000000010011001101010;
    rom[56604] = 25'b0000000000010011001011110;
    rom[56605] = 25'b0000000000010011001010011;
    rom[56606] = 25'b0000000000010011001001000;
    rom[56607] = 25'b0000000000010011000111101;
    rom[56608] = 25'b0000000000010011000110001;
    rom[56609] = 25'b0000000000010011000100110;
    rom[56610] = 25'b0000000000010011000011010;
    rom[56611] = 25'b0000000000010011000001111;
    rom[56612] = 25'b0000000000010011000000100;
    rom[56613] = 25'b0000000000010010111111000;
    rom[56614] = 25'b0000000000010010111101101;
    rom[56615] = 25'b0000000000010010111100010;
    rom[56616] = 25'b0000000000010010111010110;
    rom[56617] = 25'b0000000000010010111001010;
    rom[56618] = 25'b0000000000010010110111111;
    rom[56619] = 25'b0000000000010010110110100;
    rom[56620] = 25'b0000000000010010110101001;
    rom[56621] = 25'b0000000000010010110011101;
    rom[56622] = 25'b0000000000010010110010010;
    rom[56623] = 25'b0000000000010010110000110;
    rom[56624] = 25'b0000000000010010101111010;
    rom[56625] = 25'b0000000000010010101101111;
    rom[56626] = 25'b0000000000010010101100100;
    rom[56627] = 25'b0000000000010010101011000;
    rom[56628] = 25'b0000000000010010101001101;
    rom[56629] = 25'b0000000000010010101000001;
    rom[56630] = 25'b0000000000010010100110110;
    rom[56631] = 25'b0000000000010010100101011;
    rom[56632] = 25'b0000000000010010100011111;
    rom[56633] = 25'b0000000000010010100010011;
    rom[56634] = 25'b0000000000010010100000111;
    rom[56635] = 25'b0000000000010010011111100;
    rom[56636] = 25'b0000000000010010011110001;
    rom[56637] = 25'b0000000000010010011100101;
    rom[56638] = 25'b0000000000010010011011010;
    rom[56639] = 25'b0000000000010010011001110;
    rom[56640] = 25'b0000000000010010011000011;
    rom[56641] = 25'b0000000000010010010110111;
    rom[56642] = 25'b0000000000010010010101100;
    rom[56643] = 25'b0000000000010010010100000;
    rom[56644] = 25'b0000000000010010010010100;
    rom[56645] = 25'b0000000000010010010001000;
    rom[56646] = 25'b0000000000010010001111101;
    rom[56647] = 25'b0000000000010010001110001;
    rom[56648] = 25'b0000000000010010001100110;
    rom[56649] = 25'b0000000000010010001011010;
    rom[56650] = 25'b0000000000010010001001111;
    rom[56651] = 25'b0000000000010010001000011;
    rom[56652] = 25'b0000000000010010000111000;
    rom[56653] = 25'b0000000000010010000101100;
    rom[56654] = 25'b0000000000010010000100001;
    rom[56655] = 25'b0000000000010010000010101;
    rom[56656] = 25'b0000000000010010000001001;
    rom[56657] = 25'b0000000000010001111111101;
    rom[56658] = 25'b0000000000010001111110001;
    rom[56659] = 25'b0000000000010001111100110;
    rom[56660] = 25'b0000000000010001111011010;
    rom[56661] = 25'b0000000000010001111001110;
    rom[56662] = 25'b0000000000010001111000011;
    rom[56663] = 25'b0000000000010001110110111;
    rom[56664] = 25'b0000000000010001110101100;
    rom[56665] = 25'b0000000000010001110100000;
    rom[56666] = 25'b0000000000010001110010100;
    rom[56667] = 25'b0000000000010001110001001;
    rom[56668] = 25'b0000000000010001101111101;
    rom[56669] = 25'b0000000000010001101110001;
    rom[56670] = 25'b0000000000010001101100110;
    rom[56671] = 25'b0000000000010001101011010;
    rom[56672] = 25'b0000000000010001101001110;
    rom[56673] = 25'b0000000000010001101000011;
    rom[56674] = 25'b0000000000010001100110111;
    rom[56675] = 25'b0000000000010001100101011;
    rom[56676] = 25'b0000000000010001100100000;
    rom[56677] = 25'b0000000000010001100010100;
    rom[56678] = 25'b0000000000010001100001000;
    rom[56679] = 25'b0000000000010001011111100;
    rom[56680] = 25'b0000000000010001011110000;
    rom[56681] = 25'b0000000000010001011100101;
    rom[56682] = 25'b0000000000010001011011001;
    rom[56683] = 25'b0000000000010001011001101;
    rom[56684] = 25'b0000000000010001011000001;
    rom[56685] = 25'b0000000000010001010110101;
    rom[56686] = 25'b0000000000010001010101010;
    rom[56687] = 25'b0000000000010001010011110;
    rom[56688] = 25'b0000000000010001010010010;
    rom[56689] = 25'b0000000000010001010000110;
    rom[56690] = 25'b0000000000010001001111010;
    rom[56691] = 25'b0000000000010001001101110;
    rom[56692] = 25'b0000000000010001001100011;
    rom[56693] = 25'b0000000000010001001010111;
    rom[56694] = 25'b0000000000010001001001011;
    rom[56695] = 25'b0000000000010001000111111;
    rom[56696] = 25'b0000000000010001000110011;
    rom[56697] = 25'b0000000000010001000101000;
    rom[56698] = 25'b0000000000010001000011100;
    rom[56699] = 25'b0000000000010001000010000;
    rom[56700] = 25'b0000000000010001000000100;
    rom[56701] = 25'b0000000000010000111111000;
    rom[56702] = 25'b0000000000010000111101100;
    rom[56703] = 25'b0000000000010000111100001;
    rom[56704] = 25'b0000000000010000111010101;
    rom[56705] = 25'b0000000000010000111001001;
    rom[56706] = 25'b0000000000010000110111101;
    rom[56707] = 25'b0000000000010000110110001;
    rom[56708] = 25'b0000000000010000110100110;
    rom[56709] = 25'b0000000000010000110011010;
    rom[56710] = 25'b0000000000010000110001110;
    rom[56711] = 25'b0000000000010000110000010;
    rom[56712] = 25'b0000000000010000101110110;
    rom[56713] = 25'b0000000000010000101101010;
    rom[56714] = 25'b0000000000010000101011110;
    rom[56715] = 25'b0000000000010000101010010;
    rom[56716] = 25'b0000000000010000101000110;
    rom[56717] = 25'b0000000000010000100111010;
    rom[56718] = 25'b0000000000010000100101110;
    rom[56719] = 25'b0000000000010000100100010;
    rom[56720] = 25'b0000000000010000100010110;
    rom[56721] = 25'b0000000000010000100001010;
    rom[56722] = 25'b0000000000010000011111110;
    rom[56723] = 25'b0000000000010000011110010;
    rom[56724] = 25'b0000000000010000011100110;
    rom[56725] = 25'b0000000000010000011011010;
    rom[56726] = 25'b0000000000010000011001110;
    rom[56727] = 25'b0000000000010000011000010;
    rom[56728] = 25'b0000000000010000010110110;
    rom[56729] = 25'b0000000000010000010101010;
    rom[56730] = 25'b0000000000010000010011111;
    rom[56731] = 25'b0000000000010000010010011;
    rom[56732] = 25'b0000000000010000010000111;
    rom[56733] = 25'b0000000000010000001111011;
    rom[56734] = 25'b0000000000010000001101111;
    rom[56735] = 25'b0000000000010000001100011;
    rom[56736] = 25'b0000000000010000001010111;
    rom[56737] = 25'b0000000000010000001001011;
    rom[56738] = 25'b0000000000010000000111111;
    rom[56739] = 25'b0000000000010000000110011;
    rom[56740] = 25'b0000000000010000000100111;
    rom[56741] = 25'b0000000000010000000011011;
    rom[56742] = 25'b0000000000010000000001111;
    rom[56743] = 25'b0000000000010000000000011;
    rom[56744] = 25'b0000000000001111111110111;
    rom[56745] = 25'b0000000000001111111101011;
    rom[56746] = 25'b0000000000001111111011111;
    rom[56747] = 25'b0000000000001111111010011;
    rom[56748] = 25'b0000000000001111111000111;
    rom[56749] = 25'b0000000000001111110111011;
    rom[56750] = 25'b0000000000001111110101111;
    rom[56751] = 25'b0000000000001111110100011;
    rom[56752] = 25'b0000000000001111110010111;
    rom[56753] = 25'b0000000000001111110001011;
    rom[56754] = 25'b0000000000001111101111111;
    rom[56755] = 25'b0000000000001111101110010;
    rom[56756] = 25'b0000000000001111101100110;
    rom[56757] = 25'b0000000000001111101011010;
    rom[56758] = 25'b0000000000001111101001110;
    rom[56759] = 25'b0000000000001111101000010;
    rom[56760] = 25'b0000000000001111100110110;
    rom[56761] = 25'b0000000000001111100101010;
    rom[56762] = 25'b0000000000001111100011110;
    rom[56763] = 25'b0000000000001111100010010;
    rom[56764] = 25'b0000000000001111100000110;
    rom[56765] = 25'b0000000000001111011111010;
    rom[56766] = 25'b0000000000001111011101110;
    rom[56767] = 25'b0000000000001111011100001;
    rom[56768] = 25'b0000000000001111011010101;
    rom[56769] = 25'b0000000000001111011001001;
    rom[56770] = 25'b0000000000001111010111101;
    rom[56771] = 25'b0000000000001111010110001;
    rom[56772] = 25'b0000000000001111010100101;
    rom[56773] = 25'b0000000000001111010011001;
    rom[56774] = 25'b0000000000001111010001101;
    rom[56775] = 25'b0000000000001111010000001;
    rom[56776] = 25'b0000000000001111001110101;
    rom[56777] = 25'b0000000000001111001101000;
    rom[56778] = 25'b0000000000001111001011100;
    rom[56779] = 25'b0000000000001111001010000;
    rom[56780] = 25'b0000000000001111001000100;
    rom[56781] = 25'b0000000000001111000111000;
    rom[56782] = 25'b0000000000001111000101100;
    rom[56783] = 25'b0000000000001111000100000;
    rom[56784] = 25'b0000000000001111000010100;
    rom[56785] = 25'b0000000000001111000000111;
    rom[56786] = 25'b0000000000001110111111011;
    rom[56787] = 25'b0000000000001110111101111;
    rom[56788] = 25'b0000000000001110111100011;
    rom[56789] = 25'b0000000000001110111010111;
    rom[56790] = 25'b0000000000001110111001011;
    rom[56791] = 25'b0000000000001110110111111;
    rom[56792] = 25'b0000000000001110110110011;
    rom[56793] = 25'b0000000000001110110100110;
    rom[56794] = 25'b0000000000001110110011010;
    rom[56795] = 25'b0000000000001110110001110;
    rom[56796] = 25'b0000000000001110110000001;
    rom[56797] = 25'b0000000000001110101110101;
    rom[56798] = 25'b0000000000001110101101001;
    rom[56799] = 25'b0000000000001110101011110;
    rom[56800] = 25'b0000000000001110101010001;
    rom[56801] = 25'b0000000000001110101000101;
    rom[56802] = 25'b0000000000001110100111001;
    rom[56803] = 25'b0000000000001110100101100;
    rom[56804] = 25'b0000000000001110100100000;
    rom[56805] = 25'b0000000000001110100010100;
    rom[56806] = 25'b0000000000001110100001000;
    rom[56807] = 25'b0000000000001110011111100;
    rom[56808] = 25'b0000000000001110011110000;
    rom[56809] = 25'b0000000000001110011100011;
    rom[56810] = 25'b0000000000001110011010111;
    rom[56811] = 25'b0000000000001110011001011;
    rom[56812] = 25'b0000000000001110010111110;
    rom[56813] = 25'b0000000000001110010110010;
    rom[56814] = 25'b0000000000001110010100110;
    rom[56815] = 25'b0000000000001110010011010;
    rom[56816] = 25'b0000000000001110010001110;
    rom[56817] = 25'b0000000000001110010000010;
    rom[56818] = 25'b0000000000001110001110101;
    rom[56819] = 25'b0000000000001110001101001;
    rom[56820] = 25'b0000000000001110001011101;
    rom[56821] = 25'b0000000000001110001010001;
    rom[56822] = 25'b0000000000001110001000101;
    rom[56823] = 25'b0000000000001110000111001;
    rom[56824] = 25'b0000000000001110000101100;
    rom[56825] = 25'b0000000000001110000100000;
    rom[56826] = 25'b0000000000001110000010011;
    rom[56827] = 25'b0000000000001110000000111;
    rom[56828] = 25'b0000000000001101111111011;
    rom[56829] = 25'b0000000000001101111101111;
    rom[56830] = 25'b0000000000001101111100011;
    rom[56831] = 25'b0000000000001101111010110;
    rom[56832] = 25'b0000000000001101111001010;
    rom[56833] = 25'b0000000000001101110111110;
    rom[56834] = 25'b0000000000001101110110001;
    rom[56835] = 25'b0000000000001101110100101;
    rom[56836] = 25'b0000000000001101110011010;
    rom[56837] = 25'b0000000000001101110001101;
    rom[56838] = 25'b0000000000001101110000001;
    rom[56839] = 25'b0000000000001101101110100;
    rom[56840] = 25'b0000000000001101101101000;
    rom[56841] = 25'b0000000000001101101011100;
    rom[56842] = 25'b0000000000001101101010000;
    rom[56843] = 25'b0000000000001101101000100;
    rom[56844] = 25'b0000000000001101100110111;
    rom[56845] = 25'b0000000000001101100101011;
    rom[56846] = 25'b0000000000001101100011110;
    rom[56847] = 25'b0000000000001101100010010;
    rom[56848] = 25'b0000000000001101100000110;
    rom[56849] = 25'b0000000000001101011111010;
    rom[56850] = 25'b0000000000001101011101110;
    rom[56851] = 25'b0000000000001101011100001;
    rom[56852] = 25'b0000000000001101011010101;
    rom[56853] = 25'b0000000000001101011001000;
    rom[56854] = 25'b0000000000001101010111100;
    rom[56855] = 25'b0000000000001101010110000;
    rom[56856] = 25'b0000000000001101010100100;
    rom[56857] = 25'b0000000000001101010011000;
    rom[56858] = 25'b0000000000001101010001011;
    rom[56859] = 25'b0000000000001101001111111;
    rom[56860] = 25'b0000000000001101001110010;
    rom[56861] = 25'b0000000000001101001100110;
    rom[56862] = 25'b0000000000001101001011010;
    rom[56863] = 25'b0000000000001101001001110;
    rom[56864] = 25'b0000000000001101001000010;
    rom[56865] = 25'b0000000000001101000110101;
    rom[56866] = 25'b0000000000001101000101001;
    rom[56867] = 25'b0000000000001101000011101;
    rom[56868] = 25'b0000000000001101000010001;
    rom[56869] = 25'b0000000000001101000000100;
    rom[56870] = 25'b0000000000001100111111000;
    rom[56871] = 25'b0000000000001100111101011;
    rom[56872] = 25'b0000000000001100111011111;
    rom[56873] = 25'b0000000000001100111010011;
    rom[56874] = 25'b0000000000001100111000111;
    rom[56875] = 25'b0000000000001100110111011;
    rom[56876] = 25'b0000000000001100110101110;
    rom[56877] = 25'b0000000000001100110100010;
    rom[56878] = 25'b0000000000001100110010101;
    rom[56879] = 25'b0000000000001100110001001;
    rom[56880] = 25'b0000000000001100101111101;
    rom[56881] = 25'b0000000000001100101110001;
    rom[56882] = 25'b0000000000001100101100100;
    rom[56883] = 25'b0000000000001100101011000;
    rom[56884] = 25'b0000000000001100101001011;
    rom[56885] = 25'b0000000000001100100111111;
    rom[56886] = 25'b0000000000001100100110011;
    rom[56887] = 25'b0000000000001100100100111;
    rom[56888] = 25'b0000000000001100100011010;
    rom[56889] = 25'b0000000000001100100001110;
    rom[56890] = 25'b0000000000001100100000001;
    rom[56891] = 25'b0000000000001100011110101;
    rom[56892] = 25'b0000000000001100011101001;
    rom[56893] = 25'b0000000000001100011011101;
    rom[56894] = 25'b0000000000001100011010000;
    rom[56895] = 25'b0000000000001100011000100;
    rom[56896] = 25'b0000000000001100010110111;
    rom[56897] = 25'b0000000000001100010101011;
    rom[56898] = 25'b0000000000001100010011111;
    rom[56899] = 25'b0000000000001100010010011;
    rom[56900] = 25'b0000000000001100010000111;
    rom[56901] = 25'b0000000000001100001111010;
    rom[56902] = 25'b0000000000001100001101110;
    rom[56903] = 25'b0000000000001100001100001;
    rom[56904] = 25'b0000000000001100001010110;
    rom[56905] = 25'b0000000000001100001001001;
    rom[56906] = 25'b0000000000001100000111101;
    rom[56907] = 25'b0000000000001100000110000;
    rom[56908] = 25'b0000000000001100000100100;
    rom[56909] = 25'b0000000000001100000011000;
    rom[56910] = 25'b0000000000001100000001100;
    rom[56911] = 25'b0000000000001011111111111;
    rom[56912] = 25'b0000000000001011111110011;
    rom[56913] = 25'b0000000000001011111100110;
    rom[56914] = 25'b0000000000001011111011010;
    rom[56915] = 25'b0000000000001011111001110;
    rom[56916] = 25'b0000000000001011111000010;
    rom[56917] = 25'b0000000000001011110110101;
    rom[56918] = 25'b0000000000001011110101001;
    rom[56919] = 25'b0000000000001011110011100;
    rom[56920] = 25'b0000000000001011110010000;
    rom[56921] = 25'b0000000000001011110000100;
    rom[56922] = 25'b0000000000001011101111000;
    rom[56923] = 25'b0000000000001011101101011;
    rom[56924] = 25'b0000000000001011101011111;
    rom[56925] = 25'b0000000000001011101010010;
    rom[56926] = 25'b0000000000001011101000110;
    rom[56927] = 25'b0000000000001011100111010;
    rom[56928] = 25'b0000000000001011100101110;
    rom[56929] = 25'b0000000000001011100100001;
    rom[56930] = 25'b0000000000001011100010101;
    rom[56931] = 25'b0000000000001011100001000;
    rom[56932] = 25'b0000000000001011011111100;
    rom[56933] = 25'b0000000000001011011110000;
    rom[56934] = 25'b0000000000001011011100100;
    rom[56935] = 25'b0000000000001011011010111;
    rom[56936] = 25'b0000000000001011011001011;
    rom[56937] = 25'b0000000000001011010111110;
    rom[56938] = 25'b0000000000001011010110010;
    rom[56939] = 25'b0000000000001011010100110;
    rom[56940] = 25'b0000000000001011010011010;
    rom[56941] = 25'b0000000000001011010001101;
    rom[56942] = 25'b0000000000001011010000001;
    rom[56943] = 25'b0000000000001011001110100;
    rom[56944] = 25'b0000000000001011001101000;
    rom[56945] = 25'b0000000000001011001011100;
    rom[56946] = 25'b0000000000001011001010000;
    rom[56947] = 25'b0000000000001011001000011;
    rom[56948] = 25'b0000000000001011000110111;
    rom[56949] = 25'b0000000000001011000101010;
    rom[56950] = 25'b0000000000001011000011110;
    rom[56951] = 25'b0000000000001011000010010;
    rom[56952] = 25'b0000000000001011000000110;
    rom[56953] = 25'b0000000000001010111111001;
    rom[56954] = 25'b0000000000001010111101101;
    rom[56955] = 25'b0000000000001010111100000;
    rom[56956] = 25'b0000000000001010111010101;
    rom[56957] = 25'b0000000000001010111001001;
    rom[56958] = 25'b0000000000001010110111100;
    rom[56959] = 25'b0000000000001010110110000;
    rom[56960] = 25'b0000000000001010110100011;
    rom[56961] = 25'b0000000000001010110010111;
    rom[56962] = 25'b0000000000001010110001011;
    rom[56963] = 25'b0000000000001010101111111;
    rom[56964] = 25'b0000000000001010101110010;
    rom[56965] = 25'b0000000000001010101100110;
    rom[56966] = 25'b0000000000001010101011001;
    rom[56967] = 25'b0000000000001010101001101;
    rom[56968] = 25'b0000000000001010101000001;
    rom[56969] = 25'b0000000000001010100110101;
    rom[56970] = 25'b0000000000001010100101000;
    rom[56971] = 25'b0000000000001010100011100;
    rom[56972] = 25'b0000000000001010100001111;
    rom[56973] = 25'b0000000000001010100000011;
    rom[56974] = 25'b0000000000001010011110111;
    rom[56975] = 25'b0000000000001010011101011;
    rom[56976] = 25'b0000000000001010011011111;
    rom[56977] = 25'b0000000000001010011010010;
    rom[56978] = 25'b0000000000001010011000110;
    rom[56979] = 25'b0000000000001010010111001;
    rom[56980] = 25'b0000000000001010010101101;
    rom[56981] = 25'b0000000000001010010100001;
    rom[56982] = 25'b0000000000001010010010101;
    rom[56983] = 25'b0000000000001010010001000;
    rom[56984] = 25'b0000000000001010001111100;
    rom[56985] = 25'b0000000000001010001101111;
    rom[56986] = 25'b0000000000001010001100011;
    rom[56987] = 25'b0000000000001010001011000;
    rom[56988] = 25'b0000000000001010001001011;
    rom[56989] = 25'b0000000000001010000111111;
    rom[56990] = 25'b0000000000001010000110010;
    rom[56991] = 25'b0000000000001010000100110;
    rom[56992] = 25'b0000000000001010000011001;
    rom[56993] = 25'b0000000000001010000001110;
    rom[56994] = 25'b0000000000001010000000001;
    rom[56995] = 25'b0000000000001001111110101;
    rom[56996] = 25'b0000000000001001111101001;
    rom[56997] = 25'b0000000000001001111011100;
    rom[56998] = 25'b0000000000001001111010000;
    rom[56999] = 25'b0000000000001001111000100;
    rom[57000] = 25'b0000000000001001110111000;
    rom[57001] = 25'b0000000000001001110101011;
    rom[57002] = 25'b0000000000001001110011111;
    rom[57003] = 25'b0000000000001001110010011;
    rom[57004] = 25'b0000000000001001110000110;
    rom[57005] = 25'b0000000000001001101111010;
    rom[57006] = 25'b0000000000001001101101110;
    rom[57007] = 25'b0000000000001001101100010;
    rom[57008] = 25'b0000000000001001101010101;
    rom[57009] = 25'b0000000000001001101001001;
    rom[57010] = 25'b0000000000001001100111101;
    rom[57011] = 25'b0000000000001001100110000;
    rom[57012] = 25'b0000000000001001100100100;
    rom[57013] = 25'b0000000000001001100011000;
    rom[57014] = 25'b0000000000001001100001100;
    rom[57015] = 25'b0000000000001001100000000;
    rom[57016] = 25'b0000000000001001011110011;
    rom[57017] = 25'b0000000000001001011100111;
    rom[57018] = 25'b0000000000001001011011010;
    rom[57019] = 25'b0000000000001001011001111;
    rom[57020] = 25'b0000000000001001011000011;
    rom[57021] = 25'b0000000000001001010110110;
    rom[57022] = 25'b0000000000001001010101010;
    rom[57023] = 25'b0000000000001001010011110;
    rom[57024] = 25'b0000000000001001010010001;
    rom[57025] = 25'b0000000000001001010000101;
    rom[57026] = 25'b0000000000001001001111001;
    rom[57027] = 25'b0000000000001001001101101;
    rom[57028] = 25'b0000000000001001001100001;
    rom[57029] = 25'b0000000000001001001010100;
    rom[57030] = 25'b0000000000001001001001000;
    rom[57031] = 25'b0000000000001001000111100;
    rom[57032] = 25'b0000000000001001000101111;
    rom[57033] = 25'b0000000000001001000100011;
    rom[57034] = 25'b0000000000001001000010111;
    rom[57035] = 25'b0000000000001001000001011;
    rom[57036] = 25'b0000000000001000111111111;
    rom[57037] = 25'b0000000000001000111110010;
    rom[57038] = 25'b0000000000001000111100110;
    rom[57039] = 25'b0000000000001000111011010;
    rom[57040] = 25'b0000000000001000111001110;
    rom[57041] = 25'b0000000000001000111000010;
    rom[57042] = 25'b0000000000001000110110110;
    rom[57043] = 25'b0000000000001000110101001;
    rom[57044] = 25'b0000000000001000110011101;
    rom[57045] = 25'b0000000000001000110010001;
    rom[57046] = 25'b0000000000001000110000100;
    rom[57047] = 25'b0000000000001000101111000;
    rom[57048] = 25'b0000000000001000101101100;
    rom[57049] = 25'b0000000000001000101100000;
    rom[57050] = 25'b0000000000001000101010100;
    rom[57051] = 25'b0000000000001000101001000;
    rom[57052] = 25'b0000000000001000100111100;
    rom[57053] = 25'b0000000000001000100101111;
    rom[57054] = 25'b0000000000001000100100011;
    rom[57055] = 25'b0000000000001000100010111;
    rom[57056] = 25'b0000000000001000100001011;
    rom[57057] = 25'b0000000000001000011111111;
    rom[57058] = 25'b0000000000001000011110011;
    rom[57059] = 25'b0000000000001000011100111;
    rom[57060] = 25'b0000000000001000011011010;
    rom[57061] = 25'b0000000000001000011001110;
    rom[57062] = 25'b0000000000001000011000010;
    rom[57063] = 25'b0000000000001000010110101;
    rom[57064] = 25'b0000000000001000010101001;
    rom[57065] = 25'b0000000000001000010011101;
    rom[57066] = 25'b0000000000001000010010010;
    rom[57067] = 25'b0000000000001000010000101;
    rom[57068] = 25'b0000000000001000001111001;
    rom[57069] = 25'b0000000000001000001101101;
    rom[57070] = 25'b0000000000001000001100001;
    rom[57071] = 25'b0000000000001000001010100;
    rom[57072] = 25'b0000000000001000001001000;
    rom[57073] = 25'b0000000000001000000111100;
    rom[57074] = 25'b0000000000001000000110000;
    rom[57075] = 25'b0000000000001000000100100;
    rom[57076] = 25'b0000000000001000000011000;
    rom[57077] = 25'b0000000000001000000001100;
    rom[57078] = 25'b0000000000001000000000000;
    rom[57079] = 25'b0000000000000111111110100;
    rom[57080] = 25'b0000000000000111111100111;
    rom[57081] = 25'b0000000000000111111011011;
    rom[57082] = 25'b0000000000000111111001111;
    rom[57083] = 25'b0000000000000111111000011;
    rom[57084] = 25'b0000000000000111110110111;
    rom[57085] = 25'b0000000000000111110101011;
    rom[57086] = 25'b0000000000000111110011111;
    rom[57087] = 25'b0000000000000111110010011;
    rom[57088] = 25'b0000000000000111110000111;
    rom[57089] = 25'b0000000000000111101111011;
    rom[57090] = 25'b0000000000000111101101110;
    rom[57091] = 25'b0000000000000111101100010;
    rom[57092] = 25'b0000000000000111101010110;
    rom[57093] = 25'b0000000000000111101001010;
    rom[57094] = 25'b0000000000000111100111110;
    rom[57095] = 25'b0000000000000111100110010;
    rom[57096] = 25'b0000000000000111100100110;
    rom[57097] = 25'b0000000000000111100011010;
    rom[57098] = 25'b0000000000000111100001110;
    rom[57099] = 25'b0000000000000111100000010;
    rom[57100] = 25'b0000000000000111011110110;
    rom[57101] = 25'b0000000000000111011101010;
    rom[57102] = 25'b0000000000000111011011110;
    rom[57103] = 25'b0000000000000111011010001;
    rom[57104] = 25'b0000000000000111011000101;
    rom[57105] = 25'b0000000000000111010111001;
    rom[57106] = 25'b0000000000000111010101101;
    rom[57107] = 25'b0000000000000111010100001;
    rom[57108] = 25'b0000000000000111010010101;
    rom[57109] = 25'b0000000000000111010001010;
    rom[57110] = 25'b0000000000000111001111110;
    rom[57111] = 25'b0000000000000111001110010;
    rom[57112] = 25'b0000000000000111001100101;
    rom[57113] = 25'b0000000000000111001011001;
    rom[57114] = 25'b0000000000000111001001101;
    rom[57115] = 25'b0000000000000111001000001;
    rom[57116] = 25'b0000000000000111000110101;
    rom[57117] = 25'b0000000000000111000101001;
    rom[57118] = 25'b0000000000000111000011101;
    rom[57119] = 25'b0000000000000111000010001;
    rom[57120] = 25'b0000000000000111000000101;
    rom[57121] = 25'b0000000000000110111111001;
    rom[57122] = 25'b0000000000000110111101101;
    rom[57123] = 25'b0000000000000110111100001;
    rom[57124] = 25'b0000000000000110111010101;
    rom[57125] = 25'b0000000000000110111001010;
    rom[57126] = 25'b0000000000000110110111110;
    rom[57127] = 25'b0000000000000110110110010;
    rom[57128] = 25'b0000000000000110110100110;
    rom[57129] = 25'b0000000000000110110011010;
    rom[57130] = 25'b0000000000000110110001110;
    rom[57131] = 25'b0000000000000110110000010;
    rom[57132] = 25'b0000000000000110101110110;
    rom[57133] = 25'b0000000000000110101101010;
    rom[57134] = 25'b0000000000000110101011110;
    rom[57135] = 25'b0000000000000110101010010;
    rom[57136] = 25'b0000000000000110101000110;
    rom[57137] = 25'b0000000000000110100111010;
    rom[57138] = 25'b0000000000000110100101110;
    rom[57139] = 25'b0000000000000110100100010;
    rom[57140] = 25'b0000000000000110100010110;
    rom[57141] = 25'b0000000000000110100001010;
    rom[57142] = 25'b0000000000000110011111110;
    rom[57143] = 25'b0000000000000110011110010;
    rom[57144] = 25'b0000000000000110011100110;
    rom[57145] = 25'b0000000000000110011011010;
    rom[57146] = 25'b0000000000000110011001111;
    rom[57147] = 25'b0000000000000110011000011;
    rom[57148] = 25'b0000000000000110010110111;
    rom[57149] = 25'b0000000000000110010101011;
    rom[57150] = 25'b0000000000000110010011111;
    rom[57151] = 25'b0000000000000110010010011;
    rom[57152] = 25'b0000000000000110010001000;
    rom[57153] = 25'b0000000000000110001111100;
    rom[57154] = 25'b0000000000000110001110000;
    rom[57155] = 25'b0000000000000110001100100;
    rom[57156] = 25'b0000000000000110001011000;
    rom[57157] = 25'b0000000000000110001001100;
    rom[57158] = 25'b0000000000000110001000000;
    rom[57159] = 25'b0000000000000110000110100;
    rom[57160] = 25'b0000000000000110000101001;
    rom[57161] = 25'b0000000000000110000011101;
    rom[57162] = 25'b0000000000000110000010001;
    rom[57163] = 25'b0000000000000110000000101;
    rom[57164] = 25'b0000000000000101111111001;
    rom[57165] = 25'b0000000000000101111101101;
    rom[57166] = 25'b0000000000000101111100001;
    rom[57167] = 25'b0000000000000101111010110;
    rom[57168] = 25'b0000000000000101111001010;
    rom[57169] = 25'b0000000000000101110111110;
    rom[57170] = 25'b0000000000000101110110010;
    rom[57171] = 25'b0000000000000101110100110;
    rom[57172] = 25'b0000000000000101110011011;
    rom[57173] = 25'b0000000000000101110001111;
    rom[57174] = 25'b0000000000000101110000011;
    rom[57175] = 25'b0000000000000101101110111;
    rom[57176] = 25'b0000000000000101101101011;
    rom[57177] = 25'b0000000000000101101100000;
    rom[57178] = 25'b0000000000000101101010100;
    rom[57179] = 25'b0000000000000101101001000;
    rom[57180] = 25'b0000000000000101100111100;
    rom[57181] = 25'b0000000000000101100110001;
    rom[57182] = 25'b0000000000000101100100101;
    rom[57183] = 25'b0000000000000101100011001;
    rom[57184] = 25'b0000000000000101100001101;
    rom[57185] = 25'b0000000000000101100000010;
    rom[57186] = 25'b0000000000000101011110110;
    rom[57187] = 25'b0000000000000101011101010;
    rom[57188] = 25'b0000000000000101011011110;
    rom[57189] = 25'b0000000000000101011010010;
    rom[57190] = 25'b0000000000000101011000111;
    rom[57191] = 25'b0000000000000101010111011;
    rom[57192] = 25'b0000000000000101010101111;
    rom[57193] = 25'b0000000000000101010100011;
    rom[57194] = 25'b0000000000000101010010111;
    rom[57195] = 25'b0000000000000101010001100;
    rom[57196] = 25'b0000000000000101010000000;
    rom[57197] = 25'b0000000000000101001110100;
    rom[57198] = 25'b0000000000000101001101001;
    rom[57199] = 25'b0000000000000101001011101;
    rom[57200] = 25'b0000000000000101001010001;
    rom[57201] = 25'b0000000000000101001000110;
    rom[57202] = 25'b0000000000000101000111010;
    rom[57203] = 25'b0000000000000101000101111;
    rom[57204] = 25'b0000000000000101000100011;
    rom[57205] = 25'b0000000000000101000010111;
    rom[57206] = 25'b0000000000000101000001100;
    rom[57207] = 25'b0000000000000101000000000;
    rom[57208] = 25'b0000000000000100111110101;
    rom[57209] = 25'b0000000000000100111101001;
    rom[57210] = 25'b0000000000000100111011101;
    rom[57211] = 25'b0000000000000100111010001;
    rom[57212] = 25'b0000000000000100111000110;
    rom[57213] = 25'b0000000000000100110111010;
    rom[57214] = 25'b0000000000000100110101110;
    rom[57215] = 25'b0000000000000100110100011;
    rom[57216] = 25'b0000000000000100110010111;
    rom[57217] = 25'b0000000000000100110001011;
    rom[57218] = 25'b0000000000000100110000000;
    rom[57219] = 25'b0000000000000100101110100;
    rom[57220] = 25'b0000000000000100101101001;
    rom[57221] = 25'b0000000000000100101011101;
    rom[57222] = 25'b0000000000000100101010010;
    rom[57223] = 25'b0000000000000100101000110;
    rom[57224] = 25'b0000000000000100100111011;
    rom[57225] = 25'b0000000000000100100101111;
    rom[57226] = 25'b0000000000000100100100011;
    rom[57227] = 25'b0000000000000100100010111;
    rom[57228] = 25'b0000000000000100100001100;
    rom[57229] = 25'b0000000000000100100000001;
    rom[57230] = 25'b0000000000000100011110101;
    rom[57231] = 25'b0000000000000100011101010;
    rom[57232] = 25'b0000000000000100011011110;
    rom[57233] = 25'b0000000000000100011010011;
    rom[57234] = 25'b0000000000000100011000111;
    rom[57235] = 25'b0000000000000100010111100;
    rom[57236] = 25'b0000000000000100010110000;
    rom[57237] = 25'b0000000000000100010100100;
    rom[57238] = 25'b0000000000000100010011001;
    rom[57239] = 25'b0000000000000100010001101;
    rom[57240] = 25'b0000000000000100010000010;
    rom[57241] = 25'b0000000000000100001110111;
    rom[57242] = 25'b0000000000000100001101011;
    rom[57243] = 25'b0000000000000100001100000;
    rom[57244] = 25'b0000000000000100001010100;
    rom[57245] = 25'b0000000000000100001001001;
    rom[57246] = 25'b0000000000000100000111101;
    rom[57247] = 25'b0000000000000100000110001;
    rom[57248] = 25'b0000000000000100000100110;
    rom[57249] = 25'b0000000000000100000011011;
    rom[57250] = 25'b0000000000000100000001111;
    rom[57251] = 25'b0000000000000100000000100;
    rom[57252] = 25'b0000000000000011111111001;
    rom[57253] = 25'b0000000000000011111101101;
    rom[57254] = 25'b0000000000000011111100001;
    rom[57255] = 25'b0000000000000011111010110;
    rom[57256] = 25'b0000000000000011111001011;
    rom[57257] = 25'b0000000000000011110111111;
    rom[57258] = 25'b0000000000000011110110100;
    rom[57259] = 25'b0000000000000011110101001;
    rom[57260] = 25'b0000000000000011110011101;
    rom[57261] = 25'b0000000000000011110010001;
    rom[57262] = 25'b0000000000000011110000110;
    rom[57263] = 25'b0000000000000011101111011;
    rom[57264] = 25'b0000000000000011101110000;
    rom[57265] = 25'b0000000000000011101100100;
    rom[57266] = 25'b0000000000000011101011001;
    rom[57267] = 25'b0000000000000011101001101;
    rom[57268] = 25'b0000000000000011101000010;
    rom[57269] = 25'b0000000000000011100110111;
    rom[57270] = 25'b0000000000000011100101011;
    rom[57271] = 25'b0000000000000011100100000;
    rom[57272] = 25'b0000000000000011100010101;
    rom[57273] = 25'b0000000000000011100001001;
    rom[57274] = 25'b0000000000000011011111110;
    rom[57275] = 25'b0000000000000011011110011;
    rom[57276] = 25'b0000000000000011011101000;
    rom[57277] = 25'b0000000000000011011011100;
    rom[57278] = 25'b0000000000000011011010001;
    rom[57279] = 25'b0000000000000011011000110;
    rom[57280] = 25'b0000000000000011010111010;
    rom[57281] = 25'b0000000000000011010101111;
    rom[57282] = 25'b0000000000000011010100100;
    rom[57283] = 25'b0000000000000011010011001;
    rom[57284] = 25'b0000000000000011010001101;
    rom[57285] = 25'b0000000000000011010000010;
    rom[57286] = 25'b0000000000000011001110111;
    rom[57287] = 25'b0000000000000011001101100;
    rom[57288] = 25'b0000000000000011001100000;
    rom[57289] = 25'b0000000000000011001010101;
    rom[57290] = 25'b0000000000000011001001001;
    rom[57291] = 25'b0000000000000011000111110;
    rom[57292] = 25'b0000000000000011000110011;
    rom[57293] = 25'b0000000000000011000101000;
    rom[57294] = 25'b0000000000000011000011101;
    rom[57295] = 25'b0000000000000011000010001;
    rom[57296] = 25'b0000000000000011000000110;
    rom[57297] = 25'b0000000000000010111111011;
    rom[57298] = 25'b0000000000000010111110000;
    rom[57299] = 25'b0000000000000010111100101;
    rom[57300] = 25'b0000000000000010111011010;
    rom[57301] = 25'b0000000000000010111001111;
    rom[57302] = 25'b0000000000000010111000100;
    rom[57303] = 25'b0000000000000010110111001;
    rom[57304] = 25'b0000000000000010110101101;
    rom[57305] = 25'b0000000000000010110100010;
    rom[57306] = 25'b0000000000000010110010111;
    rom[57307] = 25'b0000000000000010110001100;
    rom[57308] = 25'b0000000000000010110000001;
    rom[57309] = 25'b0000000000000010101110101;
    rom[57310] = 25'b0000000000000010101101010;
    rom[57311] = 25'b0000000000000010101100000;
    rom[57312] = 25'b0000000000000010101010100;
    rom[57313] = 25'b0000000000000010101001001;
    rom[57314] = 25'b0000000000000010100111110;
    rom[57315] = 25'b0000000000000010100110011;
    rom[57316] = 25'b0000000000000010100101000;
    rom[57317] = 25'b0000000000000010100011100;
    rom[57318] = 25'b0000000000000010100010010;
    rom[57319] = 25'b0000000000000010100000111;
    rom[57320] = 25'b0000000000000010011111100;
    rom[57321] = 25'b0000000000000010011110000;
    rom[57322] = 25'b0000000000000010011100101;
    rom[57323] = 25'b0000000000000010011011011;
    rom[57324] = 25'b0000000000000010011001111;
    rom[57325] = 25'b0000000000000010011000100;
    rom[57326] = 25'b0000000000000010010111001;
    rom[57327] = 25'b0000000000000010010101111;
    rom[57328] = 25'b0000000000000010010100011;
    rom[57329] = 25'b0000000000000010010011000;
    rom[57330] = 25'b0000000000000010010001110;
    rom[57331] = 25'b0000000000000010010000011;
    rom[57332] = 25'b0000000000000010001110111;
    rom[57333] = 25'b0000000000000010001101100;
    rom[57334] = 25'b0000000000000010001100010;
    rom[57335] = 25'b0000000000000010001010110;
    rom[57336] = 25'b0000000000000010001001011;
    rom[57337] = 25'b0000000000000010001000001;
    rom[57338] = 25'b0000000000000010000110110;
    rom[57339] = 25'b0000000000000010000101010;
    rom[57340] = 25'b0000000000000010000100000;
    rom[57341] = 25'b0000000000000010000010101;
    rom[57342] = 25'b0000000000000010000001010;
    rom[57343] = 25'b0000000000000001111111111;
    rom[57344] = 25'b0000000000000001111110100;
    rom[57345] = 25'b0000000000000001111101001;
    rom[57346] = 25'b0000000000000001111011110;
    rom[57347] = 25'b0000000000000001111010100;
    rom[57348] = 25'b0000000000000001111001000;
    rom[57349] = 25'b0000000000000001110111110;
    rom[57350] = 25'b0000000000000001110110011;
    rom[57351] = 25'b0000000000000001110101000;
    rom[57352] = 25'b0000000000000001110011101;
    rom[57353] = 25'b0000000000000001110010010;
    rom[57354] = 25'b0000000000000001110000111;
    rom[57355] = 25'b0000000000000001101111100;
    rom[57356] = 25'b0000000000000001101110010;
    rom[57357] = 25'b0000000000000001101100111;
    rom[57358] = 25'b0000000000000001101011100;
    rom[57359] = 25'b0000000000000001101010001;
    rom[57360] = 25'b0000000000000001101000110;
    rom[57361] = 25'b0000000000000001100111011;
    rom[57362] = 25'b0000000000000001100110001;
    rom[57363] = 25'b0000000000000001100100110;
    rom[57364] = 25'b0000000000000001100011011;
    rom[57365] = 25'b0000000000000001100010001;
    rom[57366] = 25'b0000000000000001100000101;
    rom[57367] = 25'b0000000000000001011111011;
    rom[57368] = 25'b0000000000000001011110001;
    rom[57369] = 25'b0000000000000001011100101;
    rom[57370] = 25'b0000000000000001011011011;
    rom[57371] = 25'b0000000000000001011010000;
    rom[57372] = 25'b0000000000000001011000101;
    rom[57373] = 25'b0000000000000001010111011;
    rom[57374] = 25'b0000000000000001010110000;
    rom[57375] = 25'b0000000000000001010100101;
    rom[57376] = 25'b0000000000000001010011011;
    rom[57377] = 25'b0000000000000001010001111;
    rom[57378] = 25'b0000000000000001010000101;
    rom[57379] = 25'b0000000000000001001111011;
    rom[57380] = 25'b0000000000000001001110000;
    rom[57381] = 25'b0000000000000001001100101;
    rom[57382] = 25'b0000000000000001001011010;
    rom[57383] = 25'b0000000000000001001010000;
    rom[57384] = 25'b0000000000000001001000101;
    rom[57385] = 25'b0000000000000001000111010;
    rom[57386] = 25'b0000000000000001000110000;
    rom[57387] = 25'b0000000000000001000100101;
    rom[57388] = 25'b0000000000000001000011011;
    rom[57389] = 25'b0000000000000001000010000;
    rom[57390] = 25'b0000000000000001000000101;
    rom[57391] = 25'b0000000000000000111111011;
    rom[57392] = 25'b0000000000000000111110000;
    rom[57393] = 25'b0000000000000000111100110;
    rom[57394] = 25'b0000000000000000111011011;
    rom[57395] = 25'b0000000000000000111010000;
    rom[57396] = 25'b0000000000000000111000110;
    rom[57397] = 25'b0000000000000000110111011;
    rom[57398] = 25'b0000000000000000110110001;
    rom[57399] = 25'b0000000000000000110100110;
    rom[57400] = 25'b0000000000000000110011100;
    rom[57401] = 25'b0000000000000000110010001;
    rom[57402] = 25'b0000000000000000110000111;
    rom[57403] = 25'b0000000000000000101111100;
    rom[57404] = 25'b0000000000000000101110001;
    rom[57405] = 25'b0000000000000000101100111;
    rom[57406] = 25'b0000000000000000101011100;
    rom[57407] = 25'b0000000000000000101010010;
    rom[57408] = 25'b0000000000000000101000111;
    rom[57409] = 25'b0000000000000000100111101;
    rom[57410] = 25'b0000000000000000100110011;
    rom[57411] = 25'b0000000000000000100101000;
    rom[57412] = 25'b0000000000000000100011110;
    rom[57413] = 25'b0000000000000000100010011;
    rom[57414] = 25'b0000000000000000100001001;
    rom[57415] = 25'b0000000000000000011111110;
    rom[57416] = 25'b0000000000000000011110100;
    rom[57417] = 25'b0000000000000000011101001;
    rom[57418] = 25'b0000000000000000011011111;
    rom[57419] = 25'b0000000000000000011010101;
    rom[57420] = 25'b0000000000000000011001011;
    rom[57421] = 25'b0000000000000000011000000;
    rom[57422] = 25'b0000000000000000010110110;
    rom[57423] = 25'b0000000000000000010101011;
    rom[57424] = 25'b0000000000000000010100001;
    rom[57425] = 25'b0000000000000000010010110;
    rom[57426] = 25'b0000000000000000010001100;
    rom[57427] = 25'b0000000000000000010000001;
    rom[57428] = 25'b0000000000000000001111000;
    rom[57429] = 25'b0000000000000000001101101;
    rom[57430] = 25'b0000000000000000001100011;
    rom[57431] = 25'b0000000000000000001011000;
    rom[57432] = 25'b0000000000000000001001110;
    rom[57433] = 25'b0000000000000000001000100;
    rom[57434] = 25'b0000000000000000000111010;
    rom[57435] = 25'b0000000000000000000101111;
    rom[57436] = 25'b0000000000000000000100101;
    rom[57437] = 25'b0000000000000000000011010;
    rom[57438] = 25'b0000000000000000000010001;
    rom[57439] = 25'b0000000000000000000000110;
    rom[57440] = 25'b1111111111111111111111101;
    rom[57441] = 25'b1111111111111111111110011;
    rom[57442] = 25'b1111111111111111111101000;
    rom[57443] = 25'b1111111111111111111011110;
    rom[57444] = 25'b1111111111111111111010011;
    rom[57445] = 25'b1111111111111111111001010;
    rom[57446] = 25'b1111111111111111110111111;
    rom[57447] = 25'b1111111111111111110110110;
    rom[57448] = 25'b1111111111111111110101011;
    rom[57449] = 25'b1111111111111111110100001;
    rom[57450] = 25'b1111111111111111110010111;
    rom[57451] = 25'b1111111111111111110001100;
    rom[57452] = 25'b1111111111111111110000010;
    rom[57453] = 25'b1111111111111111101111000;
    rom[57454] = 25'b1111111111111111101101110;
    rom[57455] = 25'b1111111111111111101100100;
    rom[57456] = 25'b1111111111111111101011010;
    rom[57457] = 25'b1111111111111111101010000;
    rom[57458] = 25'b1111111111111111101000101;
    rom[57459] = 25'b1111111111111111100111011;
    rom[57460] = 25'b1111111111111111100110001;
    rom[57461] = 25'b1111111111111111100100111;
    rom[57462] = 25'b1111111111111111100011101;
    rom[57463] = 25'b1111111111111111100010011;
    rom[57464] = 25'b1111111111111111100001001;
    rom[57465] = 25'b1111111111111111011111110;
    rom[57466] = 25'b1111111111111111011110101;
    rom[57467] = 25'b1111111111111111011101011;
    rom[57468] = 25'b1111111111111111011100001;
    rom[57469] = 25'b1111111111111111011010111;
    rom[57470] = 25'b1111111111111111011001100;
    rom[57471] = 25'b1111111111111111011000011;
    rom[57472] = 25'b1111111111111111010111000;
    rom[57473] = 25'b1111111111111111010101111;
    rom[57474] = 25'b1111111111111111010100101;
    rom[57475] = 25'b1111111111111111010011010;
    rom[57476] = 25'b1111111111111111010010001;
    rom[57477] = 25'b1111111111111111010000111;
    rom[57478] = 25'b1111111111111111001111101;
    rom[57479] = 25'b1111111111111111001110011;
    rom[57480] = 25'b1111111111111111001101001;
    rom[57481] = 25'b1111111111111111001011111;
    rom[57482] = 25'b1111111111111111001010101;
    rom[57483] = 25'b1111111111111111001001011;
    rom[57484] = 25'b1111111111111111001000001;
    rom[57485] = 25'b1111111111111111000110111;
    rom[57486] = 25'b1111111111111111000101101;
    rom[57487] = 25'b1111111111111111000100100;
    rom[57488] = 25'b1111111111111111000011001;
    rom[57489] = 25'b1111111111111111000001111;
    rom[57490] = 25'b1111111111111111000000110;
    rom[57491] = 25'b1111111111111110111111100;
    rom[57492] = 25'b1111111111111110111110010;
    rom[57493] = 25'b1111111111111110111101000;
    rom[57494] = 25'b1111111111111110111011110;
    rom[57495] = 25'b1111111111111110111010100;
    rom[57496] = 25'b1111111111111110111001011;
    rom[57497] = 25'b1111111111111110111000001;
    rom[57498] = 25'b1111111111111110110110111;
    rom[57499] = 25'b1111111111111110110101101;
    rom[57500] = 25'b1111111111111110110100011;
    rom[57501] = 25'b1111111111111110110011001;
    rom[57502] = 25'b1111111111111110110010000;
    rom[57503] = 25'b1111111111111110110000110;
    rom[57504] = 25'b1111111111111110101111100;
    rom[57505] = 25'b1111111111111110101110011;
    rom[57506] = 25'b1111111111111110101101001;
    rom[57507] = 25'b1111111111111110101011111;
    rom[57508] = 25'b1111111111111110101010101;
    rom[57509] = 25'b1111111111111110101001100;
    rom[57510] = 25'b1111111111111110101000010;
    rom[57511] = 25'b1111111111111110100111000;
    rom[57512] = 25'b1111111111111110100101111;
    rom[57513] = 25'b1111111111111110100100101;
    rom[57514] = 25'b1111111111111110100011011;
    rom[57515] = 25'b1111111111111110100010001;
    rom[57516] = 25'b1111111111111110100001000;
    rom[57517] = 25'b1111111111111110011111110;
    rom[57518] = 25'b1111111111111110011110100;
    rom[57519] = 25'b1111111111111110011101011;
    rom[57520] = 25'b1111111111111110011100001;
    rom[57521] = 25'b1111111111111110011010111;
    rom[57522] = 25'b1111111111111110011001110;
    rom[57523] = 25'b1111111111111110011000100;
    rom[57524] = 25'b1111111111111110010111011;
    rom[57525] = 25'b1111111111111110010110001;
    rom[57526] = 25'b1111111111111110010100111;
    rom[57527] = 25'b1111111111111110010011110;
    rom[57528] = 25'b1111111111111110010010101;
    rom[57529] = 25'b1111111111111110010001011;
    rom[57530] = 25'b1111111111111110010000001;
    rom[57531] = 25'b1111111111111110001111000;
    rom[57532] = 25'b1111111111111110001101110;
    rom[57533] = 25'b1111111111111110001100101;
    rom[57534] = 25'b1111111111111110001011011;
    rom[57535] = 25'b1111111111111110001010001;
    rom[57536] = 25'b1111111111111110001001000;
    rom[57537] = 25'b1111111111111110000111111;
    rom[57538] = 25'b1111111111111110000110101;
    rom[57539] = 25'b1111111111111110000101011;
    rom[57540] = 25'b1111111111111110000100010;
    rom[57541] = 25'b1111111111111110000011001;
    rom[57542] = 25'b1111111111111110000001111;
    rom[57543] = 25'b1111111111111110000000110;
    rom[57544] = 25'b1111111111111101111111100;
    rom[57545] = 25'b1111111111111101111110011;
    rom[57546] = 25'b1111111111111101111101010;
    rom[57547] = 25'b1111111111111101111100000;
    rom[57548] = 25'b1111111111111101111010111;
    rom[57549] = 25'b1111111111111101111001101;
    rom[57550] = 25'b1111111111111101111000100;
    rom[57551] = 25'b1111111111111101110111010;
    rom[57552] = 25'b1111111111111101110110001;
    rom[57553] = 25'b1111111111111101110101000;
    rom[57554] = 25'b1111111111111101110011110;
    rom[57555] = 25'b1111111111111101110010101;
    rom[57556] = 25'b1111111111111101110001011;
    rom[57557] = 25'b1111111111111101110000010;
    rom[57558] = 25'b1111111111111101101111001;
    rom[57559] = 25'b1111111111111101101110000;
    rom[57560] = 25'b1111111111111101101100110;
    rom[57561] = 25'b1111111111111101101011101;
    rom[57562] = 25'b1111111111111101101010100;
    rom[57563] = 25'b1111111111111101101001010;
    rom[57564] = 25'b1111111111111101101000001;
    rom[57565] = 25'b1111111111111101100111000;
    rom[57566] = 25'b1111111111111101100101111;
    rom[57567] = 25'b1111111111111101100100110;
    rom[57568] = 25'b1111111111111101100011100;
    rom[57569] = 25'b1111111111111101100010011;
    rom[57570] = 25'b1111111111111101100001001;
    rom[57571] = 25'b1111111111111101100000000;
    rom[57572] = 25'b1111111111111101011111000;
    rom[57573] = 25'b1111111111111101011101111;
    rom[57574] = 25'b1111111111111101011100101;
    rom[57575] = 25'b1111111111111101011011100;
    rom[57576] = 25'b1111111111111101011010011;
    rom[57577] = 25'b1111111111111101011001001;
    rom[57578] = 25'b1111111111111101011000000;
    rom[57579] = 25'b1111111111111101010110111;
    rom[57580] = 25'b1111111111111101010101110;
    rom[57581] = 25'b1111111111111101010100101;
    rom[57582] = 25'b1111111111111101010011100;
    rom[57583] = 25'b1111111111111101010010011;
    rom[57584] = 25'b1111111111111101010001010;
    rom[57585] = 25'b1111111111111101010000001;
    rom[57586] = 25'b1111111111111101001111000;
    rom[57587] = 25'b1111111111111101001101110;
    rom[57588] = 25'b1111111111111101001100101;
    rom[57589] = 25'b1111111111111101001011100;
    rom[57590] = 25'b1111111111111101001010011;
    rom[57591] = 25'b1111111111111101001001010;
    rom[57592] = 25'b1111111111111101001000001;
    rom[57593] = 25'b1111111111111101000111000;
    rom[57594] = 25'b1111111111111101000101111;
    rom[57595] = 25'b1111111111111101000100110;
    rom[57596] = 25'b1111111111111101000011101;
    rom[57597] = 25'b1111111111111101000010100;
    rom[57598] = 25'b1111111111111101000001011;
    rom[57599] = 25'b1111111111111101000000010;
    rom[57600] = 25'b1111111111111100111111001;
    rom[57601] = 25'b1111111111111100111110000;
    rom[57602] = 25'b1111111111111100111101000;
    rom[57603] = 25'b1111111111111100111011111;
    rom[57604] = 25'b1111111111111100111010110;
    rom[57605] = 25'b1111111111111100111001101;
    rom[57606] = 25'b1111111111111100111000100;
    rom[57607] = 25'b1111111111111100110111011;
    rom[57608] = 25'b1111111111111100110110010;
    rom[57609] = 25'b1111111111111100110101001;
    rom[57610] = 25'b1111111111111100110100000;
    rom[57611] = 25'b1111111111111100110010111;
    rom[57612] = 25'b1111111111111100110001110;
    rom[57613] = 25'b1111111111111100110000110;
    rom[57614] = 25'b1111111111111100101111101;
    rom[57615] = 25'b1111111111111100101110100;
    rom[57616] = 25'b1111111111111100101101011;
    rom[57617] = 25'b1111111111111100101100010;
    rom[57618] = 25'b1111111111111100101011001;
    rom[57619] = 25'b1111111111111100101010001;
    rom[57620] = 25'b1111111111111100101001000;
    rom[57621] = 25'b1111111111111100100111111;
    rom[57622] = 25'b1111111111111100100110110;
    rom[57623] = 25'b1111111111111100100101110;
    rom[57624] = 25'b1111111111111100100100101;
    rom[57625] = 25'b1111111111111100100011100;
    rom[57626] = 25'b1111111111111100100010011;
    rom[57627] = 25'b1111111111111100100001010;
    rom[57628] = 25'b1111111111111100100000001;
    rom[57629] = 25'b1111111111111100011111001;
    rom[57630] = 25'b1111111111111100011110000;
    rom[57631] = 25'b1111111111111100011100111;
    rom[57632] = 25'b1111111111111100011011111;
    rom[57633] = 25'b1111111111111100011010110;
    rom[57634] = 25'b1111111111111100011001101;
    rom[57635] = 25'b1111111111111100011000101;
    rom[57636] = 25'b1111111111111100010111100;
    rom[57637] = 25'b1111111111111100010110100;
    rom[57638] = 25'b1111111111111100010101011;
    rom[57639] = 25'b1111111111111100010100011;
    rom[57640] = 25'b1111111111111100010011010;
    rom[57641] = 25'b1111111111111100010010001;
    rom[57642] = 25'b1111111111111100010001000;
    rom[57643] = 25'b1111111111111100010000000;
    rom[57644] = 25'b1111111111111100001110111;
    rom[57645] = 25'b1111111111111100001101111;
    rom[57646] = 25'b1111111111111100001100110;
    rom[57647] = 25'b1111111111111100001011110;
    rom[57648] = 25'b1111111111111100001010101;
    rom[57649] = 25'b1111111111111100001001101;
    rom[57650] = 25'b1111111111111100001000100;
    rom[57651] = 25'b1111111111111100000111011;
    rom[57652] = 25'b1111111111111100000110011;
    rom[57653] = 25'b1111111111111100000101010;
    rom[57654] = 25'b1111111111111100000100010;
    rom[57655] = 25'b1111111111111100000011010;
    rom[57656] = 25'b1111111111111100000010001;
    rom[57657] = 25'b1111111111111100000001001;
    rom[57658] = 25'b1111111111111100000000000;
    rom[57659] = 25'b1111111111111011111110111;
    rom[57660] = 25'b1111111111111011111101111;
    rom[57661] = 25'b1111111111111011111100111;
    rom[57662] = 25'b1111111111111011111011111;
    rom[57663] = 25'b1111111111111011111010110;
    rom[57664] = 25'b1111111111111011111001110;
    rom[57665] = 25'b1111111111111011111000101;
    rom[57666] = 25'b1111111111111011110111101;
    rom[57667] = 25'b1111111111111011110110100;
    rom[57668] = 25'b1111111111111011110101100;
    rom[57669] = 25'b1111111111111011110100100;
    rom[57670] = 25'b1111111111111011110011100;
    rom[57671] = 25'b1111111111111011110010011;
    rom[57672] = 25'b1111111111111011110001011;
    rom[57673] = 25'b1111111111111011110000010;
    rom[57674] = 25'b1111111111111011101111010;
    rom[57675] = 25'b1111111111111011101110010;
    rom[57676] = 25'b1111111111111011101101010;
    rom[57677] = 25'b1111111111111011101100001;
    rom[57678] = 25'b1111111111111011101011001;
    rom[57679] = 25'b1111111111111011101010001;
    rom[57680] = 25'b1111111111111011101001001;
    rom[57681] = 25'b1111111111111011101000000;
    rom[57682] = 25'b1111111111111011100111000;
    rom[57683] = 25'b1111111111111011100110000;
    rom[57684] = 25'b1111111111111011100101000;
    rom[57685] = 25'b1111111111111011100100000;
    rom[57686] = 25'b1111111111111011100010111;
    rom[57687] = 25'b1111111111111011100001111;
    rom[57688] = 25'b1111111111111011100000111;
    rom[57689] = 25'b1111111111111011011111111;
    rom[57690] = 25'b1111111111111011011110110;
    rom[57691] = 25'b1111111111111011011101110;
    rom[57692] = 25'b1111111111111011011100110;
    rom[57693] = 25'b1111111111111011011011110;
    rom[57694] = 25'b1111111111111011011010110;
    rom[57695] = 25'b1111111111111011011001110;
    rom[57696] = 25'b1111111111111011011000110;
    rom[57697] = 25'b1111111111111011010111110;
    rom[57698] = 25'b1111111111111011010110101;
    rom[57699] = 25'b1111111111111011010101101;
    rom[57700] = 25'b1111111111111011010100110;
    rom[57701] = 25'b1111111111111011010011110;
    rom[57702] = 25'b1111111111111011010010101;
    rom[57703] = 25'b1111111111111011010001101;
    rom[57704] = 25'b1111111111111011010000110;
    rom[57705] = 25'b1111111111111011001111101;
    rom[57706] = 25'b1111111111111011001110101;
    rom[57707] = 25'b1111111111111011001101101;
    rom[57708] = 25'b1111111111111011001100110;
    rom[57709] = 25'b1111111111111011001011101;
    rom[57710] = 25'b1111111111111011001010101;
    rom[57711] = 25'b1111111111111011001001110;
    rom[57712] = 25'b1111111111111011001000101;
    rom[57713] = 25'b1111111111111011000111101;
    rom[57714] = 25'b1111111111111011000110110;
    rom[57715] = 25'b1111111111111011000101110;
    rom[57716] = 25'b1111111111111011000100110;
    rom[57717] = 25'b1111111111111011000011110;
    rom[57718] = 25'b1111111111111011000010110;
    rom[57719] = 25'b1111111111111011000001110;
    rom[57720] = 25'b1111111111111011000000110;
    rom[57721] = 25'b1111111111111010111111110;
    rom[57722] = 25'b1111111111111010111110110;
    rom[57723] = 25'b1111111111111010111101111;
    rom[57724] = 25'b1111111111111010111100111;
    rom[57725] = 25'b1111111111111010111011111;
    rom[57726] = 25'b1111111111111010111010111;
    rom[57727] = 25'b1111111111111010111001111;
    rom[57728] = 25'b1111111111111010111000111;
    rom[57729] = 25'b1111111111111010111000000;
    rom[57730] = 25'b1111111111111010110111000;
    rom[57731] = 25'b1111111111111010110110000;
    rom[57732] = 25'b1111111111111010110101001;
    rom[57733] = 25'b1111111111111010110100000;
    rom[57734] = 25'b1111111111111010110011001;
    rom[57735] = 25'b1111111111111010110010001;
    rom[57736] = 25'b1111111111111010110001001;
    rom[57737] = 25'b1111111111111010110000010;
    rom[57738] = 25'b1111111111111010101111010;
    rom[57739] = 25'b1111111111111010101110010;
    rom[57740] = 25'b1111111111111010101101011;
    rom[57741] = 25'b1111111111111010101100011;
    rom[57742] = 25'b1111111111111010101011100;
    rom[57743] = 25'b1111111111111010101010011;
    rom[57744] = 25'b1111111111111010101001100;
    rom[57745] = 25'b1111111111111010101000100;
    rom[57746] = 25'b1111111111111010100111101;
    rom[57747] = 25'b1111111111111010100110101;
    rom[57748] = 25'b1111111111111010100101101;
    rom[57749] = 25'b1111111111111010100100110;
    rom[57750] = 25'b1111111111111010100011110;
    rom[57751] = 25'b1111111111111010100010111;
    rom[57752] = 25'b1111111111111010100001111;
    rom[57753] = 25'b1111111111111010100000111;
    rom[57754] = 25'b1111111111111010100000000;
    rom[57755] = 25'b1111111111111010011111000;
    rom[57756] = 25'b1111111111111010011110001;
    rom[57757] = 25'b1111111111111010011101001;
    rom[57758] = 25'b1111111111111010011100010;
    rom[57759] = 25'b1111111111111010011011010;
    rom[57760] = 25'b1111111111111010011010011;
    rom[57761] = 25'b1111111111111010011001011;
    rom[57762] = 25'b1111111111111010011000100;
    rom[57763] = 25'b1111111111111010010111100;
    rom[57764] = 25'b1111111111111010010110101;
    rom[57765] = 25'b1111111111111010010101110;
    rom[57766] = 25'b1111111111111010010100110;
    rom[57767] = 25'b1111111111111010010011111;
    rom[57768] = 25'b1111111111111010010010111;
    rom[57769] = 25'b1111111111111010010010000;
    rom[57770] = 25'b1111111111111010010001000;
    rom[57771] = 25'b1111111111111010010000001;
    rom[57772] = 25'b1111111111111010001111010;
    rom[57773] = 25'b1111111111111010001110010;
    rom[57774] = 25'b1111111111111010001101011;
    rom[57775] = 25'b1111111111111010001100100;
    rom[57776] = 25'b1111111111111010001011100;
    rom[57777] = 25'b1111111111111010001010101;
    rom[57778] = 25'b1111111111111010001001101;
    rom[57779] = 25'b1111111111111010001000110;
    rom[57780] = 25'b1111111111111010000111111;
    rom[57781] = 25'b1111111111111010000110111;
    rom[57782] = 25'b1111111111111010000110000;
    rom[57783] = 25'b1111111111111010000101001;
    rom[57784] = 25'b1111111111111010000100010;
    rom[57785] = 25'b1111111111111010000011010;
    rom[57786] = 25'b1111111111111010000010100;
    rom[57787] = 25'b1111111111111010000001100;
    rom[57788] = 25'b1111111111111010000000101;
    rom[57789] = 25'b1111111111111001111111101;
    rom[57790] = 25'b1111111111111001111110110;
    rom[57791] = 25'b1111111111111001111101111;
    rom[57792] = 25'b1111111111111001111101000;
    rom[57793] = 25'b1111111111111001111100001;
    rom[57794] = 25'b1111111111111001111011001;
    rom[57795] = 25'b1111111111111001111010011;
    rom[57796] = 25'b1111111111111001111001011;
    rom[57797] = 25'b1111111111111001111000100;
    rom[57798] = 25'b1111111111111001110111101;
    rom[57799] = 25'b1111111111111001110110110;
    rom[57800] = 25'b1111111111111001110101111;
    rom[57801] = 25'b1111111111111001110101000;
    rom[57802] = 25'b1111111111111001110100001;
    rom[57803] = 25'b1111111111111001110011010;
    rom[57804] = 25'b1111111111111001110010010;
    rom[57805] = 25'b1111111111111001110001100;
    rom[57806] = 25'b1111111111111001110000100;
    rom[57807] = 25'b1111111111111001101111101;
    rom[57808] = 25'b1111111111111001101110110;
    rom[57809] = 25'b1111111111111001101101111;
    rom[57810] = 25'b1111111111111001101101001;
    rom[57811] = 25'b1111111111111001101100001;
    rom[57812] = 25'b1111111111111001101011010;
    rom[57813] = 25'b1111111111111001101010011;
    rom[57814] = 25'b1111111111111001101001100;
    rom[57815] = 25'b1111111111111001101000101;
    rom[57816] = 25'b1111111111111001100111110;
    rom[57817] = 25'b1111111111111001100110111;
    rom[57818] = 25'b1111111111111001100110000;
    rom[57819] = 25'b1111111111111001100101010;
    rom[57820] = 25'b1111111111111001100100010;
    rom[57821] = 25'b1111111111111001100011100;
    rom[57822] = 25'b1111111111111001100010101;
    rom[57823] = 25'b1111111111111001100001110;
    rom[57824] = 25'b1111111111111001100000111;
    rom[57825] = 25'b1111111111111001100000000;
    rom[57826] = 25'b1111111111111001011111001;
    rom[57827] = 25'b1111111111111001011110010;
    rom[57828] = 25'b1111111111111001011101100;
    rom[57829] = 25'b1111111111111001011100101;
    rom[57830] = 25'b1111111111111001011011110;
    rom[57831] = 25'b1111111111111001011010111;
    rom[57832] = 25'b1111111111111001011010000;
    rom[57833] = 25'b1111111111111001011001001;
    rom[57834] = 25'b1111111111111001011000011;
    rom[57835] = 25'b1111111111111001010111100;
    rom[57836] = 25'b1111111111111001010110101;
    rom[57837] = 25'b1111111111111001010101111;
    rom[57838] = 25'b1111111111111001010101000;
    rom[57839] = 25'b1111111111111001010100001;
    rom[57840] = 25'b1111111111111001010011010;
    rom[57841] = 25'b1111111111111001010010100;
    rom[57842] = 25'b1111111111111001010001101;
    rom[57843] = 25'b1111111111111001010000110;
    rom[57844] = 25'b1111111111111001001111111;
    rom[57845] = 25'b1111111111111001001111001;
    rom[57846] = 25'b1111111111111001001110010;
    rom[57847] = 25'b1111111111111001001101011;
    rom[57848] = 25'b1111111111111001001100101;
    rom[57849] = 25'b1111111111111001001011111;
    rom[57850] = 25'b1111111111111001001011000;
    rom[57851] = 25'b1111111111111001001010001;
    rom[57852] = 25'b1111111111111001001001010;
    rom[57853] = 25'b1111111111111001001000100;
    rom[57854] = 25'b1111111111111001000111101;
    rom[57855] = 25'b1111111111111001000110111;
    rom[57856] = 25'b1111111111111001000110000;
    rom[57857] = 25'b1111111111111001000101010;
    rom[57858] = 25'b1111111111111001000100011;
    rom[57859] = 25'b1111111111111001000011101;
    rom[57860] = 25'b1111111111111001000010110;
    rom[57861] = 25'b1111111111111001000001111;
    rom[57862] = 25'b1111111111111001000001001;
    rom[57863] = 25'b1111111111111001000000011;
    rom[57864] = 25'b1111111111111000111111100;
    rom[57865] = 25'b1111111111111000111110101;
    rom[57866] = 25'b1111111111111000111101111;
    rom[57867] = 25'b1111111111111000111101001;
    rom[57868] = 25'b1111111111111000111100010;
    rom[57869] = 25'b1111111111111000111011100;
    rom[57870] = 25'b1111111111111000111010101;
    rom[57871] = 25'b1111111111111000111001111;
    rom[57872] = 25'b1111111111111000111001000;
    rom[57873] = 25'b1111111111111000111000010;
    rom[57874] = 25'b1111111111111000110111100;
    rom[57875] = 25'b1111111111111000110110101;
    rom[57876] = 25'b1111111111111000110101111;
    rom[57877] = 25'b1111111111111000110101000;
    rom[57878] = 25'b1111111111111000110100010;
    rom[57879] = 25'b1111111111111000110011100;
    rom[57880] = 25'b1111111111111000110010110;
    rom[57881] = 25'b1111111111111000110010000;
    rom[57882] = 25'b1111111111111000110001001;
    rom[57883] = 25'b1111111111111000110000011;
    rom[57884] = 25'b1111111111111000101111100;
    rom[57885] = 25'b1111111111111000101110110;
    rom[57886] = 25'b1111111111111000101110000;
    rom[57887] = 25'b1111111111111000101101010;
    rom[57888] = 25'b1111111111111000101100100;
    rom[57889] = 25'b1111111111111000101011101;
    rom[57890] = 25'b1111111111111000101010111;
    rom[57891] = 25'b1111111111111000101010001;
    rom[57892] = 25'b1111111111111000101001010;
    rom[57893] = 25'b1111111111111000101000100;
    rom[57894] = 25'b1111111111111000100111110;
    rom[57895] = 25'b1111111111111000100111000;
    rom[57896] = 25'b1111111111111000100110001;
    rom[57897] = 25'b1111111111111000100101100;
    rom[57898] = 25'b1111111111111000100100110;
    rom[57899] = 25'b1111111111111000100100000;
    rom[57900] = 25'b1111111111111000100011010;
    rom[57901] = 25'b1111111111111000100010011;
    rom[57902] = 25'b1111111111111000100001101;
    rom[57903] = 25'b1111111111111000100000111;
    rom[57904] = 25'b1111111111111000100000001;
    rom[57905] = 25'b1111111111111000011111011;
    rom[57906] = 25'b1111111111111000011110101;
    rom[57907] = 25'b1111111111111000011101111;
    rom[57908] = 25'b1111111111111000011101000;
    rom[57909] = 25'b1111111111111000011100010;
    rom[57910] = 25'b1111111111111000011011100;
    rom[57911] = 25'b1111111111111000011010110;
    rom[57912] = 25'b1111111111111000011010000;
    rom[57913] = 25'b1111111111111000011001010;
    rom[57914] = 25'b1111111111111000011000100;
    rom[57915] = 25'b1111111111111000010111110;
    rom[57916] = 25'b1111111111111000010111000;
    rom[57917] = 25'b1111111111111000010110010;
    rom[57918] = 25'b1111111111111000010101100;
    rom[57919] = 25'b1111111111111000010100111;
    rom[57920] = 25'b1111111111111000010100001;
    rom[57921] = 25'b1111111111111000010011011;
    rom[57922] = 25'b1111111111111000010010101;
    rom[57923] = 25'b1111111111111000010001111;
    rom[57924] = 25'b1111111111111000010001001;
    rom[57925] = 25'b1111111111111000010000011;
    rom[57926] = 25'b1111111111111000001111101;
    rom[57927] = 25'b1111111111111000001110111;
    rom[57928] = 25'b1111111111111000001110001;
    rom[57929] = 25'b1111111111111000001101100;
    rom[57930] = 25'b1111111111111000001100110;
    rom[57931] = 25'b1111111111111000001100000;
    rom[57932] = 25'b1111111111111000001011010;
    rom[57933] = 25'b1111111111111000001010101;
    rom[57934] = 25'b1111111111111000001001111;
    rom[57935] = 25'b1111111111111000001001001;
    rom[57936] = 25'b1111111111111000001000011;
    rom[57937] = 25'b1111111111111000000111110;
    rom[57938] = 25'b1111111111111000000111000;
    rom[57939] = 25'b1111111111111000000110010;
    rom[57940] = 25'b1111111111111000000101101;
    rom[57941] = 25'b1111111111111000000100111;
    rom[57942] = 25'b1111111111111000000100001;
    rom[57943] = 25'b1111111111111000000011100;
    rom[57944] = 25'b1111111111111000000010110;
    rom[57945] = 25'b1111111111111000000010000;
    rom[57946] = 25'b1111111111111000000001010;
    rom[57947] = 25'b1111111111111000000000100;
    rom[57948] = 25'b1111111111110111111111111;
    rom[57949] = 25'b1111111111110111111111001;
    rom[57950] = 25'b1111111111110111111110100;
    rom[57951] = 25'b1111111111110111111101110;
    rom[57952] = 25'b1111111111110111111101001;
    rom[57953] = 25'b1111111111110111111100011;
    rom[57954] = 25'b1111111111110111111011110;
    rom[57955] = 25'b1111111111110111111011000;
    rom[57956] = 25'b1111111111110111111010010;
    rom[57957] = 25'b1111111111110111111001100;
    rom[57958] = 25'b1111111111110111111000111;
    rom[57959] = 25'b1111111111110111111000010;
    rom[57960] = 25'b1111111111110111110111100;
    rom[57961] = 25'b1111111111110111110110111;
    rom[57962] = 25'b1111111111110111110110001;
    rom[57963] = 25'b1111111111110111110101011;
    rom[57964] = 25'b1111111111110111110100110;
    rom[57965] = 25'b1111111111110111110100000;
    rom[57966] = 25'b1111111111110111110011011;
    rom[57967] = 25'b1111111111110111110010110;
    rom[57968] = 25'b1111111111110111110010001;
    rom[57969] = 25'b1111111111110111110001011;
    rom[57970] = 25'b1111111111110111110000101;
    rom[57971] = 25'b1111111111110111110000000;
    rom[57972] = 25'b1111111111110111101111011;
    rom[57973] = 25'b1111111111110111101110101;
    rom[57974] = 25'b1111111111110111101110000;
    rom[57975] = 25'b1111111111110111101101010;
    rom[57976] = 25'b1111111111110111101100101;
    rom[57977] = 25'b1111111111110111101100000;
    rom[57978] = 25'b1111111111110111101011011;
    rom[57979] = 25'b1111111111110111101010101;
    rom[57980] = 25'b1111111111110111101010000;
    rom[57981] = 25'b1111111111110111101001010;
    rom[57982] = 25'b1111111111110111101000101;
    rom[57983] = 25'b1111111111110111101000000;
    rom[57984] = 25'b1111111111110111100111011;
    rom[57985] = 25'b1111111111110111100110101;
    rom[57986] = 25'b1111111111110111100110000;
    rom[57987] = 25'b1111111111110111100101011;
    rom[57988] = 25'b1111111111110111100100110;
    rom[57989] = 25'b1111111111110111100100001;
    rom[57990] = 25'b1111111111110111100011011;
    rom[57991] = 25'b1111111111110111100010110;
    rom[57992] = 25'b1111111111110111100010001;
    rom[57993] = 25'b1111111111110111100001100;
    rom[57994] = 25'b1111111111110111100000110;
    rom[57995] = 25'b1111111111110111100000001;
    rom[57996] = 25'b1111111111110111011111100;
    rom[57997] = 25'b1111111111110111011110111;
    rom[57998] = 25'b1111111111110111011110001;
    rom[57999] = 25'b1111111111110111011101101;
    rom[58000] = 25'b1111111111110111011101000;
    rom[58001] = 25'b1111111111110111011100011;
    rom[58002] = 25'b1111111111110111011011101;
    rom[58003] = 25'b1111111111110111011011000;
    rom[58004] = 25'b1111111111110111011010011;
    rom[58005] = 25'b1111111111110111011001110;
    rom[58006] = 25'b1111111111110111011001001;
    rom[58007] = 25'b1111111111110111011000100;
    rom[58008] = 25'b1111111111110111010111111;
    rom[58009] = 25'b1111111111110111010111010;
    rom[58010] = 25'b1111111111110111010110101;
    rom[58011] = 25'b1111111111110111010110000;
    rom[58012] = 25'b1111111111110111010101011;
    rom[58013] = 25'b1111111111110111010100110;
    rom[58014] = 25'b1111111111110111010100001;
    rom[58015] = 25'b1111111111110111010011100;
    rom[58016] = 25'b1111111111110111010010111;
    rom[58017] = 25'b1111111111110111010010010;
    rom[58018] = 25'b1111111111110111010001101;
    rom[58019] = 25'b1111111111110111010001000;
    rom[58020] = 25'b1111111111110111010000100;
    rom[58021] = 25'b1111111111110111001111110;
    rom[58022] = 25'b1111111111110111001111001;
    rom[58023] = 25'b1111111111110111001110101;
    rom[58024] = 25'b1111111111110111001101111;
    rom[58025] = 25'b1111111111110111001101011;
    rom[58026] = 25'b1111111111110111001100110;
    rom[58027] = 25'b1111111111110111001100001;
    rom[58028] = 25'b1111111111110111001011100;
    rom[58029] = 25'b1111111111110111001011000;
    rom[58030] = 25'b1111111111110111001010010;
    rom[58031] = 25'b1111111111110111001001110;
    rom[58032] = 25'b1111111111110111001001001;
    rom[58033] = 25'b1111111111110111001000100;
    rom[58034] = 25'b1111111111110111001000000;
    rom[58035] = 25'b1111111111110111000111010;
    rom[58036] = 25'b1111111111110111000110110;
    rom[58037] = 25'b1111111111110111000110001;
    rom[58038] = 25'b1111111111110111000101100;
    rom[58039] = 25'b1111111111110111000101000;
    rom[58040] = 25'b1111111111110111000100011;
    rom[58041] = 25'b1111111111110111000011110;
    rom[58042] = 25'b1111111111110111000011010;
    rom[58043] = 25'b1111111111110111000010101;
    rom[58044] = 25'b1111111111110111000010001;
    rom[58045] = 25'b1111111111110111000001011;
    rom[58046] = 25'b1111111111110111000000111;
    rom[58047] = 25'b1111111111110111000000010;
    rom[58048] = 25'b1111111111110110111111110;
    rom[58049] = 25'b1111111111110110111111001;
    rom[58050] = 25'b1111111111110110111110100;
    rom[58051] = 25'b1111111111110110111110000;
    rom[58052] = 25'b1111111111110110111101011;
    rom[58053] = 25'b1111111111110110111100111;
    rom[58054] = 25'b1111111111110110111100010;
    rom[58055] = 25'b1111111111110110111011110;
    rom[58056] = 25'b1111111111110110111011001;
    rom[58057] = 25'b1111111111110110111010101;
    rom[58058] = 25'b1111111111110110111010000;
    rom[58059] = 25'b1111111111110110111001011;
    rom[58060] = 25'b1111111111110110111000111;
    rom[58061] = 25'b1111111111110110111000010;
    rom[58062] = 25'b1111111111110110110111110;
    rom[58063] = 25'b1111111111110110110111001;
    rom[58064] = 25'b1111111111110110110110101;
    rom[58065] = 25'b1111111111110110110110000;
    rom[58066] = 25'b1111111111110110110101100;
    rom[58067] = 25'b1111111111110110110101000;
    rom[58068] = 25'b1111111111110110110100100;
    rom[58069] = 25'b1111111111110110110011111;
    rom[58070] = 25'b1111111111110110110011011;
    rom[58071] = 25'b1111111111110110110010110;
    rom[58072] = 25'b1111111111110110110010010;
    rom[58073] = 25'b1111111111110110110001101;
    rom[58074] = 25'b1111111111110110110001001;
    rom[58075] = 25'b1111111111110110110000100;
    rom[58076] = 25'b1111111111110110110000000;
    rom[58077] = 25'b1111111111110110101111100;
    rom[58078] = 25'b1111111111110110101110111;
    rom[58079] = 25'b1111111111110110101110011;
    rom[58080] = 25'b1111111111110110101101110;
    rom[58081] = 25'b1111111111110110101101011;
    rom[58082] = 25'b1111111111110110101100110;
    rom[58083] = 25'b1111111111110110101100010;
    rom[58084] = 25'b1111111111110110101011110;
    rom[58085] = 25'b1111111111110110101011010;
    rom[58086] = 25'b1111111111110110101010101;
    rom[58087] = 25'b1111111111110110101010001;
    rom[58088] = 25'b1111111111110110101001101;
    rom[58089] = 25'b1111111111110110101001000;
    rom[58090] = 25'b1111111111110110101000101;
    rom[58091] = 25'b1111111111110110101000000;
    rom[58092] = 25'b1111111111110110100111100;
    rom[58093] = 25'b1111111111110110100111000;
    rom[58094] = 25'b1111111111110110100110011;
    rom[58095] = 25'b1111111111110110100110000;
    rom[58096] = 25'b1111111111110110100101011;
    rom[58097] = 25'b1111111111110110100100111;
    rom[58098] = 25'b1111111111110110100100011;
    rom[58099] = 25'b1111111111110110100011111;
    rom[58100] = 25'b1111111111110110100011011;
    rom[58101] = 25'b1111111111110110100010110;
    rom[58102] = 25'b1111111111110110100010011;
    rom[58103] = 25'b1111111111110110100001110;
    rom[58104] = 25'b1111111111110110100001010;
    rom[58105] = 25'b1111111111110110100000111;
    rom[58106] = 25'b1111111111110110100000010;
    rom[58107] = 25'b1111111111110110011111110;
    rom[58108] = 25'b1111111111110110011111010;
    rom[58109] = 25'b1111111111110110011110110;
    rom[58110] = 25'b1111111111110110011110010;
    rom[58111] = 25'b1111111111110110011101110;
    rom[58112] = 25'b1111111111110110011101010;
    rom[58113] = 25'b1111111111110110011100111;
    rom[58114] = 25'b1111111111110110011100010;
    rom[58115] = 25'b1111111111110110011011110;
    rom[58116] = 25'b1111111111110110011011011;
    rom[58117] = 25'b1111111111110110011010110;
    rom[58118] = 25'b1111111111110110011010010;
    rom[58119] = 25'b1111111111110110011001111;
    rom[58120] = 25'b1111111111110110011001011;
    rom[58121] = 25'b1111111111110110011000111;
    rom[58122] = 25'b1111111111110110011000011;
    rom[58123] = 25'b1111111111110110010111111;
    rom[58124] = 25'b1111111111110110010111011;
    rom[58125] = 25'b1111111111110110010110111;
    rom[58126] = 25'b1111111111110110010110100;
    rom[58127] = 25'b1111111111110110010101111;
    rom[58128] = 25'b1111111111110110010101011;
    rom[58129] = 25'b1111111111110110010101000;
    rom[58130] = 25'b1111111111110110010100100;
    rom[58131] = 25'b1111111111110110010100000;
    rom[58132] = 25'b1111111111110110010011101;
    rom[58133] = 25'b1111111111110110010011001;
    rom[58134] = 25'b1111111111110110010010101;
    rom[58135] = 25'b1111111111110110010010001;
    rom[58136] = 25'b1111111111110110010001110;
    rom[58137] = 25'b1111111111110110010001010;
    rom[58138] = 25'b1111111111110110010000110;
    rom[58139] = 25'b1111111111110110010000010;
    rom[58140] = 25'b1111111111110110001111111;
    rom[58141] = 25'b1111111111110110001111011;
    rom[58142] = 25'b1111111111110110001110111;
    rom[58143] = 25'b1111111111110110001110011;
    rom[58144] = 25'b1111111111110110001110000;
    rom[58145] = 25'b1111111111110110001101100;
    rom[58146] = 25'b1111111111110110001101000;
    rom[58147] = 25'b1111111111110110001100101;
    rom[58148] = 25'b1111111111110110001100010;
    rom[58149] = 25'b1111111111110110001011110;
    rom[58150] = 25'b1111111111110110001011010;
    rom[58151] = 25'b1111111111110110001010110;
    rom[58152] = 25'b1111111111110110001010011;
    rom[58153] = 25'b1111111111110110001010000;
    rom[58154] = 25'b1111111111110110001001100;
    rom[58155] = 25'b1111111111110110001001000;
    rom[58156] = 25'b1111111111110110001000100;
    rom[58157] = 25'b1111111111110110001000001;
    rom[58158] = 25'b1111111111110110000111110;
    rom[58159] = 25'b1111111111110110000111010;
    rom[58160] = 25'b1111111111110110000110110;
    rom[58161] = 25'b1111111111110110000110011;
    rom[58162] = 25'b1111111111110110000101111;
    rom[58163] = 25'b1111111111110110000101100;
    rom[58164] = 25'b1111111111110110000101001;
    rom[58165] = 25'b1111111111110110000100101;
    rom[58166] = 25'b1111111111110110000100010;
    rom[58167] = 25'b1111111111110110000011110;
    rom[58168] = 25'b1111111111110110000011011;
    rom[58169] = 25'b1111111111110110000011000;
    rom[58170] = 25'b1111111111110110000010100;
    rom[58171] = 25'b1111111111110110000010001;
    rom[58172] = 25'b1111111111110110000001101;
    rom[58173] = 25'b1111111111110110000001010;
    rom[58174] = 25'b1111111111110110000000110;
    rom[58175] = 25'b1111111111110110000000011;
    rom[58176] = 25'b1111111111110110000000000;
    rom[58177] = 25'b1111111111110101111111101;
    rom[58178] = 25'b1111111111110101111111001;
    rom[58179] = 25'b1111111111110101111110110;
    rom[58180] = 25'b1111111111110101111110010;
    rom[58181] = 25'b1111111111110101111101111;
    rom[58182] = 25'b1111111111110101111101100;
    rom[58183] = 25'b1111111111110101111101000;
    rom[58184] = 25'b1111111111110101111100110;
    rom[58185] = 25'b1111111111110101111100010;
    rom[58186] = 25'b1111111111110101111011111;
    rom[58187] = 25'b1111111111110101111011100;
    rom[58188] = 25'b1111111111110101111011000;
    rom[58189] = 25'b1111111111110101111010101;
    rom[58190] = 25'b1111111111110101111010010;
    rom[58191] = 25'b1111111111110101111001110;
    rom[58192] = 25'b1111111111110101111001011;
    rom[58193] = 25'b1111111111110101111001000;
    rom[58194] = 25'b1111111111110101111000101;
    rom[58195] = 25'b1111111111110101111000010;
    rom[58196] = 25'b1111111111110101110111111;
    rom[58197] = 25'b1111111111110101110111100;
    rom[58198] = 25'b1111111111110101110111001;
    rom[58199] = 25'b1111111111110101110110110;
    rom[58200] = 25'b1111111111110101110110011;
    rom[58201] = 25'b1111111111110101110101111;
    rom[58202] = 25'b1111111111110101110101100;
    rom[58203] = 25'b1111111111110101110101001;
    rom[58204] = 25'b1111111111110101110100110;
    rom[58205] = 25'b1111111111110101110100011;
    rom[58206] = 25'b1111111111110101110100000;
    rom[58207] = 25'b1111111111110101110011101;
    rom[58208] = 25'b1111111111110101110011010;
    rom[58209] = 25'b1111111111110101110010111;
    rom[58210] = 25'b1111111111110101110010100;
    rom[58211] = 25'b1111111111110101110010001;
    rom[58212] = 25'b1111111111110101110001110;
    rom[58213] = 25'b1111111111110101110001011;
    rom[58214] = 25'b1111111111110101110001000;
    rom[58215] = 25'b1111111111110101110000101;
    rom[58216] = 25'b1111111111110101110000010;
    rom[58217] = 25'b1111111111110101101111111;
    rom[58218] = 25'b1111111111110101101111100;
    rom[58219] = 25'b1111111111110101101111001;
    rom[58220] = 25'b1111111111110101101110110;
    rom[58221] = 25'b1111111111110101101110011;
    rom[58222] = 25'b1111111111110101101110000;
    rom[58223] = 25'b1111111111110101101101101;
    rom[58224] = 25'b1111111111110101101101011;
    rom[58225] = 25'b1111111111110101101101000;
    rom[58226] = 25'b1111111111110101101100101;
    rom[58227] = 25'b1111111111110101101100010;
    rom[58228] = 25'b1111111111110101101011111;
    rom[58229] = 25'b1111111111110101101011100;
    rom[58230] = 25'b1111111111110101101011010;
    rom[58231] = 25'b1111111111110101101010111;
    rom[58232] = 25'b1111111111110101101010100;
    rom[58233] = 25'b1111111111110101101010001;
    rom[58234] = 25'b1111111111110101101001111;
    rom[58235] = 25'b1111111111110101101001100;
    rom[58236] = 25'b1111111111110101101001001;
    rom[58237] = 25'b1111111111110101101000110;
    rom[58238] = 25'b1111111111110101101000011;
    rom[58239] = 25'b1111111111110101101000000;
    rom[58240] = 25'b1111111111110101100111110;
    rom[58241] = 25'b1111111111110101100111011;
    rom[58242] = 25'b1111111111110101100111000;
    rom[58243] = 25'b1111111111110101100110110;
    rom[58244] = 25'b1111111111110101100110011;
    rom[58245] = 25'b1111111111110101100110001;
    rom[58246] = 25'b1111111111110101100101110;
    rom[58247] = 25'b1111111111110101100101011;
    rom[58248] = 25'b1111111111110101100101000;
    rom[58249] = 25'b1111111111110101100100110;
    rom[58250] = 25'b1111111111110101100100011;
    rom[58251] = 25'b1111111111110101100100001;
    rom[58252] = 25'b1111111111110101100011110;
    rom[58253] = 25'b1111111111110101100011100;
    rom[58254] = 25'b1111111111110101100011001;
    rom[58255] = 25'b1111111111110101100010111;
    rom[58256] = 25'b1111111111110101100010100;
    rom[58257] = 25'b1111111111110101100010001;
    rom[58258] = 25'b1111111111110101100001110;
    rom[58259] = 25'b1111111111110101100001100;
    rom[58260] = 25'b1111111111110101100001010;
    rom[58261] = 25'b1111111111110101100000111;
    rom[58262] = 25'b1111111111110101100000101;
    rom[58263] = 25'b1111111111110101100000010;
    rom[58264] = 25'b1111111111110101011111111;
    rom[58265] = 25'b1111111111110101011111101;
    rom[58266] = 25'b1111111111110101011111011;
    rom[58267] = 25'b1111111111110101011111000;
    rom[58268] = 25'b1111111111110101011110110;
    rom[58269] = 25'b1111111111110101011110011;
    rom[58270] = 25'b1111111111110101011110001;
    rom[58271] = 25'b1111111111110101011101110;
    rom[58272] = 25'b1111111111110101011101100;
    rom[58273] = 25'b1111111111110101011101010;
    rom[58274] = 25'b1111111111110101011100111;
    rom[58275] = 25'b1111111111110101011100101;
    rom[58276] = 25'b1111111111110101011100010;
    rom[58277] = 25'b1111111111110101011100000;
    rom[58278] = 25'b1111111111110101011011110;
    rom[58279] = 25'b1111111111110101011011100;
    rom[58280] = 25'b1111111111110101011011001;
    rom[58281] = 25'b1111111111110101011010111;
    rom[58282] = 25'b1111111111110101011010101;
    rom[58283] = 25'b1111111111110101011010010;
    rom[58284] = 25'b1111111111110101011010000;
    rom[58285] = 25'b1111111111110101011001101;
    rom[58286] = 25'b1111111111110101011001011;
    rom[58287] = 25'b1111111111110101011001001;
    rom[58288] = 25'b1111111111110101011000111;
    rom[58289] = 25'b1111111111110101011000100;
    rom[58290] = 25'b1111111111110101011000010;
    rom[58291] = 25'b1111111111110101011000000;
    rom[58292] = 25'b1111111111110101010111110;
    rom[58293] = 25'b1111111111110101010111011;
    rom[58294] = 25'b1111111111110101010111001;
    rom[58295] = 25'b1111111111110101010111000;
    rom[58296] = 25'b1111111111110101010110101;
    rom[58297] = 25'b1111111111110101010110011;
    rom[58298] = 25'b1111111111110101010110001;
    rom[58299] = 25'b1111111111110101010101111;
    rom[58300] = 25'b1111111111110101010101100;
    rom[58301] = 25'b1111111111110101010101010;
    rom[58302] = 25'b1111111111110101010101000;
    rom[58303] = 25'b1111111111110101010100110;
    rom[58304] = 25'b1111111111110101010100100;
    rom[58305] = 25'b1111111111110101010100010;
    rom[58306] = 25'b1111111111110101010100000;
    rom[58307] = 25'b1111111111110101010011110;
    rom[58308] = 25'b1111111111110101010011100;
    rom[58309] = 25'b1111111111110101010011010;
    rom[58310] = 25'b1111111111110101010011000;
    rom[58311] = 25'b1111111111110101010010101;
    rom[58312] = 25'b1111111111110101010010100;
    rom[58313] = 25'b1111111111110101010010010;
    rom[58314] = 25'b1111111111110101010001111;
    rom[58315] = 25'b1111111111110101010001110;
    rom[58316] = 25'b1111111111110101010001100;
    rom[58317] = 25'b1111111111110101010001001;
    rom[58318] = 25'b1111111111110101010001000;
    rom[58319] = 25'b1111111111110101010000110;
    rom[58320] = 25'b1111111111110101010000011;
    rom[58321] = 25'b1111111111110101010000010;
    rom[58322] = 25'b1111111111110101010000000;
    rom[58323] = 25'b1111111111110101001111110;
    rom[58324] = 25'b1111111111110101001111100;
    rom[58325] = 25'b1111111111110101001111010;
    rom[58326] = 25'b1111111111110101001111000;
    rom[58327] = 25'b1111111111110101001110111;
    rom[58328] = 25'b1111111111110101001110100;
    rom[58329] = 25'b1111111111110101001110011;
    rom[58330] = 25'b1111111111110101001110001;
    rom[58331] = 25'b1111111111110101001101111;
    rom[58332] = 25'b1111111111110101001101101;
    rom[58333] = 25'b1111111111110101001101011;
    rom[58334] = 25'b1111111111110101001101001;
    rom[58335] = 25'b1111111111110101001101000;
    rom[58336] = 25'b1111111111110101001100101;
    rom[58337] = 25'b1111111111110101001100100;
    rom[58338] = 25'b1111111111110101001100011;
    rom[58339] = 25'b1111111111110101001100000;
    rom[58340] = 25'b1111111111110101001011111;
    rom[58341] = 25'b1111111111110101001011101;
    rom[58342] = 25'b1111111111110101001011011;
    rom[58343] = 25'b1111111111110101001011010;
    rom[58344] = 25'b1111111111110101001011000;
    rom[58345] = 25'b1111111111110101001010110;
    rom[58346] = 25'b1111111111110101001010100;
    rom[58347] = 25'b1111111111110101001010011;
    rom[58348] = 25'b1111111111110101001010001;
    rom[58349] = 25'b1111111111110101001001111;
    rom[58350] = 25'b1111111111110101001001110;
    rom[58351] = 25'b1111111111110101001001100;
    rom[58352] = 25'b1111111111110101001001011;
    rom[58353] = 25'b1111111111110101001001000;
    rom[58354] = 25'b1111111111110101001000111;
    rom[58355] = 25'b1111111111110101001000101;
    rom[58356] = 25'b1111111111110101001000100;
    rom[58357] = 25'b1111111111110101001000010;
    rom[58358] = 25'b1111111111110101001000001;
    rom[58359] = 25'b1111111111110101000111111;
    rom[58360] = 25'b1111111111110101000111101;
    rom[58361] = 25'b1111111111110101000111100;
    rom[58362] = 25'b1111111111110101000111010;
    rom[58363] = 25'b1111111111110101000111001;
    rom[58364] = 25'b1111111111110101000110111;
    rom[58365] = 25'b1111111111110101000110110;
    rom[58366] = 25'b1111111111110101000110100;
    rom[58367] = 25'b1111111111110101000110011;
    rom[58368] = 25'b1111111111110101000110001;
    rom[58369] = 25'b1111111111110101000110000;
    rom[58370] = 25'b1111111111110101000101110;
    rom[58371] = 25'b1111111111110101000101101;
    rom[58372] = 25'b1111111111110101000101011;
    rom[58373] = 25'b1111111111110101000101010;
    rom[58374] = 25'b1111111111110101000101000;
    rom[58375] = 25'b1111111111110101000100111;
    rom[58376] = 25'b1111111111110101000100101;
    rom[58377] = 25'b1111111111110101000100100;
    rom[58378] = 25'b1111111111110101000100011;
    rom[58379] = 25'b1111111111110101000100010;
    rom[58380] = 25'b1111111111110101000100000;
    rom[58381] = 25'b1111111111110101000011111;
    rom[58382] = 25'b1111111111110101000011101;
    rom[58383] = 25'b1111111111110101000011100;
    rom[58384] = 25'b1111111111110101000011010;
    rom[58385] = 25'b1111111111110101000011001;
    rom[58386] = 25'b1111111111110101000011000;
    rom[58387] = 25'b1111111111110101000010110;
    rom[58388] = 25'b1111111111110101000010101;
    rom[58389] = 25'b1111111111110101000010100;
    rom[58390] = 25'b1111111111110101000010011;
    rom[58391] = 25'b1111111111110101000010001;
    rom[58392] = 25'b1111111111110101000010000;
    rom[58393] = 25'b1111111111110101000001111;
    rom[58394] = 25'b1111111111110101000001101;
    rom[58395] = 25'b1111111111110101000001100;
    rom[58396] = 25'b1111111111110101000001011;
    rom[58397] = 25'b1111111111110101000001010;
    rom[58398] = 25'b1111111111110101000001000;
    rom[58399] = 25'b1111111111110101000000111;
    rom[58400] = 25'b1111111111110101000000110;
    rom[58401] = 25'b1111111111110101000000101;
    rom[58402] = 25'b1111111111110101000000100;
    rom[58403] = 25'b1111111111110101000000010;
    rom[58404] = 25'b1111111111110101000000001;
    rom[58405] = 25'b1111111111110101000000000;
    rom[58406] = 25'b1111111111110100111111111;
    rom[58407] = 25'b1111111111110100111111110;
    rom[58408] = 25'b1111111111110100111111101;
    rom[58409] = 25'b1111111111110100111111011;
    rom[58410] = 25'b1111111111110100111111011;
    rom[58411] = 25'b1111111111110100111111001;
    rom[58412] = 25'b1111111111110100111111000;
    rom[58413] = 25'b1111111111110100111110111;
    rom[58414] = 25'b1111111111110100111110110;
    rom[58415] = 25'b1111111111110100111110101;
    rom[58416] = 25'b1111111111110100111110100;
    rom[58417] = 25'b1111111111110100111110011;
    rom[58418] = 25'b1111111111110100111110010;
    rom[58419] = 25'b1111111111110100111110001;
    rom[58420] = 25'b1111111111110100111101111;
    rom[58421] = 25'b1111111111110100111101111;
    rom[58422] = 25'b1111111111110100111101110;
    rom[58423] = 25'b1111111111110100111101100;
    rom[58424] = 25'b1111111111110100111101100;
    rom[58425] = 25'b1111111111110100111101011;
    rom[58426] = 25'b1111111111110100111101001;
    rom[58427] = 25'b1111111111110100111101001;
    rom[58428] = 25'b1111111111110100111101000;
    rom[58429] = 25'b1111111111110100111100111;
    rom[58430] = 25'b1111111111110100111100110;
    rom[58431] = 25'b1111111111110100111100101;
    rom[58432] = 25'b1111111111110100111100100;
    rom[58433] = 25'b1111111111110100111100011;
    rom[58434] = 25'b1111111111110100111100010;
    rom[58435] = 25'b1111111111110100111100001;
    rom[58436] = 25'b1111111111110100111100001;
    rom[58437] = 25'b1111111111110100111100000;
    rom[58438] = 25'b1111111111110100111011111;
    rom[58439] = 25'b1111111111110100111011110;
    rom[58440] = 25'b1111111111110100111011110;
    rom[58441] = 25'b1111111111110100111011100;
    rom[58442] = 25'b1111111111110100111011011;
    rom[58443] = 25'b1111111111110100111011011;
    rom[58444] = 25'b1111111111110100111011010;
    rom[58445] = 25'b1111111111110100111011001;
    rom[58446] = 25'b1111111111110100111011000;
    rom[58447] = 25'b1111111111110100111011000;
    rom[58448] = 25'b1111111111110100111010111;
    rom[58449] = 25'b1111111111110100111010110;
    rom[58450] = 25'b1111111111110100111010101;
    rom[58451] = 25'b1111111111110100111010101;
    rom[58452] = 25'b1111111111110100111010100;
    rom[58453] = 25'b1111111111110100111010011;
    rom[58454] = 25'b1111111111110100111010010;
    rom[58455] = 25'b1111111111110100111010010;
    rom[58456] = 25'b1111111111110100111010001;
    rom[58457] = 25'b1111111111110100111010000;
    rom[58458] = 25'b1111111111110100111001111;
    rom[58459] = 25'b1111111111110100111001111;
    rom[58460] = 25'b1111111111110100111001110;
    rom[58461] = 25'b1111111111110100111001101;
    rom[58462] = 25'b1111111111110100111001101;
    rom[58463] = 25'b1111111111110100111001100;
    rom[58464] = 25'b1111111111110100111001100;
    rom[58465] = 25'b1111111111110100111001011;
    rom[58466] = 25'b1111111111110100111001010;
    rom[58467] = 25'b1111111111110100111001001;
    rom[58468] = 25'b1111111111110100111001001;
    rom[58469] = 25'b1111111111110100111001001;
    rom[58470] = 25'b1111111111110100111001000;
    rom[58471] = 25'b1111111111110100111000111;
    rom[58472] = 25'b1111111111110100111000111;
    rom[58473] = 25'b1111111111110100111000110;
    rom[58474] = 25'b1111111111110100111000110;
    rom[58475] = 25'b1111111111110100111000101;
    rom[58476] = 25'b1111111111110100111000101;
    rom[58477] = 25'b1111111111110100111000100;
    rom[58478] = 25'b1111111111110100111000011;
    rom[58479] = 25'b1111111111110100111000011;
    rom[58480] = 25'b1111111111110100111000011;
    rom[58481] = 25'b1111111111110100111000010;
    rom[58482] = 25'b1111111111110100111000010;
    rom[58483] = 25'b1111111111110100111000001;
    rom[58484] = 25'b1111111111110100111000000;
    rom[58485] = 25'b1111111111110100111000000;
    rom[58486] = 25'b1111111111110100111000000;
    rom[58487] = 25'b1111111111110100111000000;
    rom[58488] = 25'b1111111111110100110111111;
    rom[58489] = 25'b1111111111110100110111110;
    rom[58490] = 25'b1111111111110100110111110;
    rom[58491] = 25'b1111111111110100110111101;
    rom[58492] = 25'b1111111111110100110111101;
    rom[58493] = 25'b1111111111110100110111101;
    rom[58494] = 25'b1111111111110100110111101;
    rom[58495] = 25'b1111111111110100110111100;
    rom[58496] = 25'b1111111111110100110111100;
    rom[58497] = 25'b1111111111110100110111011;
    rom[58498] = 25'b1111111111110100110111011;
    rom[58499] = 25'b1111111111110100110111011;
    rom[58500] = 25'b1111111111110100110111010;
    rom[58501] = 25'b1111111111110100110111010;
    rom[58502] = 25'b1111111111110100110111010;
    rom[58503] = 25'b1111111111110100110111010;
    rom[58504] = 25'b1111111111110100110111010;
    rom[58505] = 25'b1111111111110100110111001;
    rom[58506] = 25'b1111111111110100110111001;
    rom[58507] = 25'b1111111111110100110111000;
    rom[58508] = 25'b1111111111110100110111000;
    rom[58509] = 25'b1111111111110100110111000;
    rom[58510] = 25'b1111111111110100110110111;
    rom[58511] = 25'b1111111111110100110110111;
    rom[58512] = 25'b1111111111110100110110111;
    rom[58513] = 25'b1111111111110100110110111;
    rom[58514] = 25'b1111111111110100110110111;
    rom[58515] = 25'b1111111111110100110110111;
    rom[58516] = 25'b1111111111110100110110111;
    rom[58517] = 25'b1111111111110100110110111;
    rom[58518] = 25'b1111111111110100110110110;
    rom[58519] = 25'b1111111111110100110110110;
    rom[58520] = 25'b1111111111110100110110110;
    rom[58521] = 25'b1111111111110100110110110;
    rom[58522] = 25'b1111111111110100110110110;
    rom[58523] = 25'b1111111111110100110110101;
    rom[58524] = 25'b1111111111110100110110101;
    rom[58525] = 25'b1111111111110100110110101;
    rom[58526] = 25'b1111111111110100110110101;
    rom[58527] = 25'b1111111111110100110110101;
    rom[58528] = 25'b1111111111110100110110101;
    rom[58529] = 25'b1111111111110100110110101;
    rom[58530] = 25'b1111111111110100110110101;
    rom[58531] = 25'b1111111111110100110110100;
    rom[58532] = 25'b1111111111110100110110100;
    rom[58533] = 25'b1111111111110100110110100;
    rom[58534] = 25'b1111111111110100110110100;
    rom[58535] = 25'b1111111111110100110110100;
    rom[58536] = 25'b1111111111110100110110100;
    rom[58537] = 25'b1111111111110100110110100;
    rom[58538] = 25'b1111111111110100110110100;
    rom[58539] = 25'b1111111111110100110110100;
    rom[58540] = 25'b1111111111110100110110100;
    rom[58541] = 25'b1111111111110100110110100;
    rom[58542] = 25'b1111111111110100110110100;
    rom[58543] = 25'b1111111111110100110110100;
    rom[58544] = 25'b1111111111110100110110100;
    rom[58545] = 25'b1111111111110100110110101;
    rom[58546] = 25'b1111111111110100110110101;
    rom[58547] = 25'b1111111111110100110110101;
    rom[58548] = 25'b1111111111110100110110101;
    rom[58549] = 25'b1111111111110100110110101;
    rom[58550] = 25'b1111111111110100110110101;
    rom[58551] = 25'b1111111111110100110110101;
    rom[58552] = 25'b1111111111110100110110101;
    rom[58553] = 25'b1111111111110100110110110;
    rom[58554] = 25'b1111111111110100110110110;
    rom[58555] = 25'b1111111111110100110110110;
    rom[58556] = 25'b1111111111110100110110110;
    rom[58557] = 25'b1111111111110100110110110;
    rom[58558] = 25'b1111111111110100110110111;
    rom[58559] = 25'b1111111111110100110110111;
    rom[58560] = 25'b1111111111110100110110111;
    rom[58561] = 25'b1111111111110100110110111;
    rom[58562] = 25'b1111111111110100110110111;
    rom[58563] = 25'b1111111111110100110110111;
    rom[58564] = 25'b1111111111110100110110111;
    rom[58565] = 25'b1111111111110100110110111;
    rom[58566] = 25'b1111111111110100110111000;
    rom[58567] = 25'b1111111111110100110111000;
    rom[58568] = 25'b1111111111110100110111000;
    rom[58569] = 25'b1111111111110100110111001;
    rom[58570] = 25'b1111111111110100110111001;
    rom[58571] = 25'b1111111111110100110111001;
    rom[58572] = 25'b1111111111110100110111010;
    rom[58573] = 25'b1111111111110100110111010;
    rom[58574] = 25'b1111111111110100110111010;
    rom[58575] = 25'b1111111111110100110111010;
    rom[58576] = 25'b1111111111110100110111010;
    rom[58577] = 25'b1111111111110100110111011;
    rom[58578] = 25'b1111111111110100110111011;
    rom[58579] = 25'b1111111111110100110111100;
    rom[58580] = 25'b1111111111110100110111100;
    rom[58581] = 25'b1111111111110100110111101;
    rom[58582] = 25'b1111111111110100110111101;
    rom[58583] = 25'b1111111111110100110111101;
    rom[58584] = 25'b1111111111110100110111101;
    rom[58585] = 25'b1111111111110100110111110;
    rom[58586] = 25'b1111111111110100110111110;
    rom[58587] = 25'b1111111111110100110111111;
    rom[58588] = 25'b1111111111110100110111111;
    rom[58589] = 25'b1111111111110100111000000;
    rom[58590] = 25'b1111111111110100111000000;
    rom[58591] = 25'b1111111111110100111000000;
    rom[58592] = 25'b1111111111110100111000001;
    rom[58593] = 25'b1111111111110100111000001;
    rom[58594] = 25'b1111111111110100111000010;
    rom[58595] = 25'b1111111111110100111000010;
    rom[58596] = 25'b1111111111110100111000011;
    rom[58597] = 25'b1111111111110100111000011;
    rom[58598] = 25'b1111111111110100111000011;
    rom[58599] = 25'b1111111111110100111000100;
    rom[58600] = 25'b1111111111110100111000101;
    rom[58601] = 25'b1111111111110100111000101;
    rom[58602] = 25'b1111111111110100111000110;
    rom[58603] = 25'b1111111111110100111000110;
    rom[58604] = 25'b1111111111110100111000111;
    rom[58605] = 25'b1111111111110100111000111;
    rom[58606] = 25'b1111111111110100111001000;
    rom[58607] = 25'b1111111111110100111001001;
    rom[58608] = 25'b1111111111110100111001001;
    rom[58609] = 25'b1111111111110100111001001;
    rom[58610] = 25'b1111111111110100111001010;
    rom[58611] = 25'b1111111111110100111001011;
    rom[58612] = 25'b1111111111110100111001100;
    rom[58613] = 25'b1111111111110100111001100;
    rom[58614] = 25'b1111111111110100111001100;
    rom[58615] = 25'b1111111111110100111001101;
    rom[58616] = 25'b1111111111110100111001110;
    rom[58617] = 25'b1111111111110100111001111;
    rom[58618] = 25'b1111111111110100111001111;
    rom[58619] = 25'b1111111111110100111010000;
    rom[58620] = 25'b1111111111110100111010000;
    rom[58621] = 25'b1111111111110100111010001;
    rom[58622] = 25'b1111111111110100111010010;
    rom[58623] = 25'b1111111111110100111010010;
    rom[58624] = 25'b1111111111110100111010011;
    rom[58625] = 25'b1111111111110100111010100;
    rom[58626] = 25'b1111111111110100111010101;
    rom[58627] = 25'b1111111111110100111010101;
    rom[58628] = 25'b1111111111110100111010110;
    rom[58629] = 25'b1111111111110100111010111;
    rom[58630] = 25'b1111111111110100111011000;
    rom[58631] = 25'b1111111111110100111011000;
    rom[58632] = 25'b1111111111110100111011001;
    rom[58633] = 25'b1111111111110100111011010;
    rom[58634] = 25'b1111111111110100111011011;
    rom[58635] = 25'b1111111111110100111011011;
    rom[58636] = 25'b1111111111110100111011100;
    rom[58637] = 25'b1111111111110100111011101;
    rom[58638] = 25'b1111111111110100111011110;
    rom[58639] = 25'b1111111111110100111011110;
    rom[58640] = 25'b1111111111110100111011111;
    rom[58641] = 25'b1111111111110100111100001;
    rom[58642] = 25'b1111111111110100111100001;
    rom[58643] = 25'b1111111111110100111100010;
    rom[58644] = 25'b1111111111110100111100011;
    rom[58645] = 25'b1111111111110100111100011;
    rom[58646] = 25'b1111111111110100111100100;
    rom[58647] = 25'b1111111111110100111100101;
    rom[58648] = 25'b1111111111110100111100110;
    rom[58649] = 25'b1111111111110100111100111;
    rom[58650] = 25'b1111111111110100111101000;
    rom[58651] = 25'b1111111111110100111101001;
    rom[58652] = 25'b1111111111110100111101001;
    rom[58653] = 25'b1111111111110100111101011;
    rom[58654] = 25'b1111111111110100111101100;
    rom[58655] = 25'b1111111111110100111101100;
    rom[58656] = 25'b1111111111110100111101101;
    rom[58657] = 25'b1111111111110100111101111;
    rom[58658] = 25'b1111111111110100111101111;
    rom[58659] = 25'b1111111111110100111110000;
    rom[58660] = 25'b1111111111110100111110001;
    rom[58661] = 25'b1111111111110100111110010;
    rom[58662] = 25'b1111111111110100111110011;
    rom[58663] = 25'b1111111111110100111110100;
    rom[58664] = 25'b1111111111110100111110101;
    rom[58665] = 25'b1111111111110100111110110;
    rom[58666] = 25'b1111111111110100111110111;
    rom[58667] = 25'b1111111111110100111111000;
    rom[58668] = 25'b1111111111110100111111001;
    rom[58669] = 25'b1111111111110100111111011;
    rom[58670] = 25'b1111111111110100111111011;
    rom[58671] = 25'b1111111111110100111111100;
    rom[58672] = 25'b1111111111110100111111110;
    rom[58673] = 25'b1111111111110100111111110;
    rom[58674] = 25'b1111111111110101000000000;
    rom[58675] = 25'b1111111111110101000000001;
    rom[58676] = 25'b1111111111110101000000010;
    rom[58677] = 25'b1111111111110101000000011;
    rom[58678] = 25'b1111111111110101000000100;
    rom[58679] = 25'b1111111111110101000000101;
    rom[58680] = 25'b1111111111110101000000111;
    rom[58681] = 25'b1111111111110101000000111;
    rom[58682] = 25'b1111111111110101000001001;
    rom[58683] = 25'b1111111111110101000001010;
    rom[58684] = 25'b1111111111110101000001011;
    rom[58685] = 25'b1111111111110101000001100;
    rom[58686] = 25'b1111111111110101000001101;
    rom[58687] = 25'b1111111111110101000001110;
    rom[58688] = 25'b1111111111110101000010000;
    rom[58689] = 25'b1111111111110101000010001;
    rom[58690] = 25'b1111111111110101000010010;
    rom[58691] = 25'b1111111111110101000010011;
    rom[58692] = 25'b1111111111110101000010100;
    rom[58693] = 25'b1111111111110101000010110;
    rom[58694] = 25'b1111111111110101000010111;
    rom[58695] = 25'b1111111111110101000011000;
    rom[58696] = 25'b1111111111110101000011001;
    rom[58697] = 25'b1111111111110101000011011;
    rom[58698] = 25'b1111111111110101000011100;
    rom[58699] = 25'b1111111111110101000011101;
    rom[58700] = 25'b1111111111110101000011111;
    rom[58701] = 25'b1111111111110101000011111;
    rom[58702] = 25'b1111111111110101000100001;
    rom[58703] = 25'b1111111111110101000100010;
    rom[58704] = 25'b1111111111110101000100011;
    rom[58705] = 25'b1111111111110101000100100;
    rom[58706] = 25'b1111111111110101000100110;
    rom[58707] = 25'b1111111111110101000100111;
    rom[58708] = 25'b1111111111110101000101001;
    rom[58709] = 25'b1111111111110101000101010;
    rom[58710] = 25'b1111111111110101000101011;
    rom[58711] = 25'b1111111111110101000101101;
    rom[58712] = 25'b1111111111110101000101110;
    rom[58713] = 25'b1111111111110101000110000;
    rom[58714] = 25'b1111111111110101000110000;
    rom[58715] = 25'b1111111111110101000110010;
    rom[58716] = 25'b1111111111110101000110011;
    rom[58717] = 25'b1111111111110101000110101;
    rom[58718] = 25'b1111111111110101000110110;
    rom[58719] = 25'b1111111111110101000111000;
    rom[58720] = 25'b1111111111110101000111001;
    rom[58721] = 25'b1111111111110101000111010;
    rom[58722] = 25'b1111111111110101000111100;
    rom[58723] = 25'b1111111111110101000111101;
    rom[58724] = 25'b1111111111110101000111111;
    rom[58725] = 25'b1111111111110101001000000;
    rom[58726] = 25'b1111111111110101001000010;
    rom[58727] = 25'b1111111111110101001000011;
    rom[58728] = 25'b1111111111110101001000101;
    rom[58729] = 25'b1111111111110101001000110;
    rom[58730] = 25'b1111111111110101001001000;
    rom[58731] = 25'b1111111111110101001001001;
    rom[58732] = 25'b1111111111110101001001011;
    rom[58733] = 25'b1111111111110101001001100;
    rom[58734] = 25'b1111111111110101001001110;
    rom[58735] = 25'b1111111111110101001001111;
    rom[58736] = 25'b1111111111110101001010001;
    rom[58737] = 25'b1111111111110101001010010;
    rom[58738] = 25'b1111111111110101001010100;
    rom[58739] = 25'b1111111111110101001010101;
    rom[58740] = 25'b1111111111110101001010111;
    rom[58741] = 25'b1111111111110101001011000;
    rom[58742] = 25'b1111111111110101001011010;
    rom[58743] = 25'b1111111111110101001011100;
    rom[58744] = 25'b1111111111110101001011101;
    rom[58745] = 25'b1111111111110101001011111;
    rom[58746] = 25'b1111111111110101001100000;
    rom[58747] = 25'b1111111111110101001100010;
    rom[58748] = 25'b1111111111110101001100011;
    rom[58749] = 25'b1111111111110101001100101;
    rom[58750] = 25'b1111111111110101001100111;
    rom[58751] = 25'b1111111111110101001101000;
    rom[58752] = 25'b1111111111110101001101010;
    rom[58753] = 25'b1111111111110101001101011;
    rom[58754] = 25'b1111111111110101001101101;
    rom[58755] = 25'b1111111111110101001101111;
    rom[58756] = 25'b1111111111110101001110001;
    rom[58757] = 25'b1111111111110101001110010;
    rom[58758] = 25'b1111111111110101001110100;
    rom[58759] = 25'b1111111111110101001110110;
    rom[58760] = 25'b1111111111110101001110111;
    rom[58761] = 25'b1111111111110101001111001;
    rom[58762] = 25'b1111111111110101001111010;
    rom[58763] = 25'b1111111111110101001111101;
    rom[58764] = 25'b1111111111110101001111110;
    rom[58765] = 25'b1111111111110101010000000;
    rom[58766] = 25'b1111111111110101010000010;
    rom[58767] = 25'b1111111111110101010000011;
    rom[58768] = 25'b1111111111110101010000101;
    rom[58769] = 25'b1111111111110101010000111;
    rom[58770] = 25'b1111111111110101010001001;
    rom[58771] = 25'b1111111111110101010001010;
    rom[58772] = 25'b1111111111110101010001100;
    rom[58773] = 25'b1111111111110101010001110;
    rom[58774] = 25'b1111111111110101010001111;
    rom[58775] = 25'b1111111111110101010010010;
    rom[58776] = 25'b1111111111110101010010011;
    rom[58777] = 25'b1111111111110101010010101;
    rom[58778] = 25'b1111111111110101010010111;
    rom[58779] = 25'b1111111111110101010011000;
    rom[58780] = 25'b1111111111110101010011011;
    rom[58781] = 25'b1111111111110101010011100;
    rom[58782] = 25'b1111111111110101010011110;
    rom[58783] = 25'b1111111111110101010100000;
    rom[58784] = 25'b1111111111110101010100010;
    rom[58785] = 25'b1111111111110101010100100;
    rom[58786] = 25'b1111111111110101010100110;
    rom[58787] = 25'b1111111111110101010100111;
    rom[58788] = 25'b1111111111110101010101001;
    rom[58789] = 25'b1111111111110101010101011;
    rom[58790] = 25'b1111111111110101010101101;
    rom[58791] = 25'b1111111111110101010101111;
    rom[58792] = 25'b1111111111110101010110001;
    rom[58793] = 25'b1111111111110101010110010;
    rom[58794] = 25'b1111111111110101010110101;
    rom[58795] = 25'b1111111111110101010110111;
    rom[58796] = 25'b1111111111110101010111000;
    rom[58797] = 25'b1111111111110101010111011;
    rom[58798] = 25'b1111111111110101010111100;
    rom[58799] = 25'b1111111111110101010111110;
    rom[58800] = 25'b1111111111110101011000001;
    rom[58801] = 25'b1111111111110101011000010;
    rom[58802] = 25'b1111111111110101011000100;
    rom[58803] = 25'b1111111111110101011000110;
    rom[58804] = 25'b1111111111110101011001000;
    rom[58805] = 25'b1111111111110101011001010;
    rom[58806] = 25'b1111111111110101011001100;
    rom[58807] = 25'b1111111111110101011001110;
    rom[58808] = 25'b1111111111110101011010000;
    rom[58809] = 25'b1111111111110101011010011;
    rom[58810] = 25'b1111111111110101011010100;
    rom[58811] = 25'b1111111111110101011010110;
    rom[58812] = 25'b1111111111110101011011001;
    rom[58813] = 25'b1111111111110101011011010;
    rom[58814] = 25'b1111111111110101011011100;
    rom[58815] = 25'b1111111111110101011011111;
    rom[58816] = 25'b1111111111110101011100001;
    rom[58817] = 25'b1111111111110101011100010;
    rom[58818] = 25'b1111111111110101011100101;
    rom[58819] = 25'b1111111111110101011100111;
    rom[58820] = 25'b1111111111110101011101001;
    rom[58821] = 25'b1111111111110101011101011;
    rom[58822] = 25'b1111111111110101011101101;
    rom[58823] = 25'b1111111111110101011101111;
    rom[58824] = 25'b1111111111110101011110001;
    rom[58825] = 25'b1111111111110101011110011;
    rom[58826] = 25'b1111111111110101011110110;
    rom[58827] = 25'b1111111111110101011110111;
    rom[58828] = 25'b1111111111110101011111001;
    rom[58829] = 25'b1111111111110101011111100;
    rom[58830] = 25'b1111111111110101011111110;
    rom[58831] = 25'b1111111111110101100000000;
    rom[58832] = 25'b1111111111110101100000010;
    rom[58833] = 25'b1111111111110101100000101;
    rom[58834] = 25'b1111111111110101100000111;
    rom[58835] = 25'b1111111111110101100001001;
    rom[58836] = 25'b1111111111110101100001011;
    rom[58837] = 25'b1111111111110101100001101;
    rom[58838] = 25'b1111111111110101100001111;
    rom[58839] = 25'b1111111111110101100010001;
    rom[58840] = 25'b1111111111110101100010100;
    rom[58841] = 25'b1111111111110101100010110;
    rom[58842] = 25'b1111111111110101100011000;
    rom[58843] = 25'b1111111111110101100011010;
    rom[58844] = 25'b1111111111110101100011101;
    rom[58845] = 25'b1111111111110101100011111;
    rom[58846] = 25'b1111111111110101100100001;
    rom[58847] = 25'b1111111111110101100100011;
    rom[58848] = 25'b1111111111110101100100101;
    rom[58849] = 25'b1111111111110101100101000;
    rom[58850] = 25'b1111111111110101100101010;
    rom[58851] = 25'b1111111111110101100101100;
    rom[58852] = 25'b1111111111110101100101110;
    rom[58853] = 25'b1111111111110101100110001;
    rom[58854] = 25'b1111111111110101100110100;
    rom[58855] = 25'b1111111111110101100110110;
    rom[58856] = 25'b1111111111110101100111000;
    rom[58857] = 25'b1111111111110101100111010;
    rom[58858] = 25'b1111111111110101100111101;
    rom[58859] = 25'b1111111111110101100111111;
    rom[58860] = 25'b1111111111110101101000001;
    rom[58861] = 25'b1111111111110101101000011;
    rom[58862] = 25'b1111111111110101101000110;
    rom[58863] = 25'b1111111111110101101001001;
    rom[58864] = 25'b1111111111110101101001011;
    rom[58865] = 25'b1111111111110101101001101;
    rom[58866] = 25'b1111111111110101101001111;
    rom[58867] = 25'b1111111111110101101010010;
    rom[58868] = 25'b1111111111110101101010100;
    rom[58869] = 25'b1111111111110101101010111;
    rom[58870] = 25'b1111111111110101101011001;
    rom[58871] = 25'b1111111111110101101011011;
    rom[58872] = 25'b1111111111110101101011110;
    rom[58873] = 25'b1111111111110101101100000;
    rom[58874] = 25'b1111111111110101101100011;
    rom[58875] = 25'b1111111111110101101100101;
    rom[58876] = 25'b1111111111110101101100111;
    rom[58877] = 25'b1111111111110101101101001;
    rom[58878] = 25'b1111111111110101101101100;
    rom[58879] = 25'b1111111111110101101101111;
    rom[58880] = 25'b1111111111110101101110001;
    rom[58881] = 25'b1111111111110101101110100;
    rom[58882] = 25'b1111111111110101101110110;
    rom[58883] = 25'b1111111111110101101111000;
    rom[58884] = 25'b1111111111110101101111011;
    rom[58885] = 25'b1111111111110101101111110;
    rom[58886] = 25'b1111111111110101110000000;
    rom[58887] = 25'b1111111111110101110000010;
    rom[58888] = 25'b1111111111110101110000101;
    rom[58889] = 25'b1111111111110101110000111;
    rom[58890] = 25'b1111111111110101110001010;
    rom[58891] = 25'b1111111111110101110001101;
    rom[58892] = 25'b1111111111110101110001111;
    rom[58893] = 25'b1111111111110101110010010;
    rom[58894] = 25'b1111111111110101110010100;
    rom[58895] = 25'b1111111111110101110010110;
    rom[58896] = 25'b1111111111110101110011001;
    rom[58897] = 25'b1111111111110101110011100;
    rom[58898] = 25'b1111111111110101110011111;
    rom[58899] = 25'b1111111111110101110100001;
    rom[58900] = 25'b1111111111110101110100100;
    rom[58901] = 25'b1111111111110101110100110;
    rom[58902] = 25'b1111111111110101110101000;
    rom[58903] = 25'b1111111111110101110101011;
    rom[58904] = 25'b1111111111110101110101101;
    rom[58905] = 25'b1111111111110101110110000;
    rom[58906] = 25'b1111111111110101110110011;
    rom[58907] = 25'b1111111111110101110110110;
    rom[58908] = 25'b1111111111110101110111000;
    rom[58909] = 25'b1111111111110101110111011;
    rom[58910] = 25'b1111111111110101110111101;
    rom[58911] = 25'b1111111111110101111000000;
    rom[58912] = 25'b1111111111110101111000010;
    rom[58913] = 25'b1111111111110101111000101;
    rom[58914] = 25'b1111111111110101111001000;
    rom[58915] = 25'b1111111111110101111001011;
    rom[58916] = 25'b1111111111110101111001110;
    rom[58917] = 25'b1111111111110101111010000;
    rom[58918] = 25'b1111111111110101111010011;
    rom[58919] = 25'b1111111111110101111010101;
    rom[58920] = 25'b1111111111110101111011000;
    rom[58921] = 25'b1111111111110101111011010;
    rom[58922] = 25'b1111111111110101111011101;
    rom[58923] = 25'b1111111111110101111100000;
    rom[58924] = 25'b1111111111110101111100011;
    rom[58925] = 25'b1111111111110101111100110;
    rom[58926] = 25'b1111111111110101111101000;
    rom[58927] = 25'b1111111111110101111101011;
    rom[58928] = 25'b1111111111110101111101110;
    rom[58929] = 25'b1111111111110101111110000;
    rom[58930] = 25'b1111111111110101111110011;
    rom[58931] = 25'b1111111111110101111110110;
    rom[58932] = 25'b1111111111110101111111000;
    rom[58933] = 25'b1111111111110101111111011;
    rom[58934] = 25'b1111111111110101111111110;
    rom[58935] = 25'b1111111111110110000000001;
    rom[58936] = 25'b1111111111110110000000011;
    rom[58937] = 25'b1111111111110110000000110;
    rom[58938] = 25'b1111111111110110000001001;
    rom[58939] = 25'b1111111111110110000001100;
    rom[58940] = 25'b1111111111110110000001111;
    rom[58941] = 25'b1111111111110110000010010;
    rom[58942] = 25'b1111111111110110000010101;
    rom[58943] = 25'b1111111111110110000010111;
    rom[58944] = 25'b1111111111110110000011010;
    rom[58945] = 25'b1111111111110110000011101;
    rom[58946] = 25'b1111111111110110000100000;
    rom[58947] = 25'b1111111111110110000100010;
    rom[58948] = 25'b1111111111110110000100101;
    rom[58949] = 25'b1111111111110110000101000;
    rom[58950] = 25'b1111111111110110000101011;
    rom[58951] = 25'b1111111111110110000101110;
    rom[58952] = 25'b1111111111110110000110000;
    rom[58953] = 25'b1111111111110110000110011;
    rom[58954] = 25'b1111111111110110000110110;
    rom[58955] = 25'b1111111111110110000111001;
    rom[58956] = 25'b1111111111110110000111100;
    rom[58957] = 25'b1111111111110110000111111;
    rom[58958] = 25'b1111111111110110001000010;
    rom[58959] = 25'b1111111111110110001000100;
    rom[58960] = 25'b1111111111110110001000111;
    rom[58961] = 25'b1111111111110110001001010;
    rom[58962] = 25'b1111111111110110001001101;
    rom[58963] = 25'b1111111111110110001010000;
    rom[58964] = 25'b1111111111110110001010011;
    rom[58965] = 25'b1111111111110110001010110;
    rom[58966] = 25'b1111111111110110001011001;
    rom[58967] = 25'b1111111111110110001011100;
    rom[58968] = 25'b1111111111110110001011111;
    rom[58969] = 25'b1111111111110110001100010;
    rom[58970] = 25'b1111111111110110001100101;
    rom[58971] = 25'b1111111111110110001100111;
    rom[58972] = 25'b1111111111110110001101010;
    rom[58973] = 25'b1111111111110110001101101;
    rom[58974] = 25'b1111111111110110001110000;
    rom[58975] = 25'b1111111111110110001110011;
    rom[58976] = 25'b1111111111110110001110110;
    rom[58977] = 25'b1111111111110110001111001;
    rom[58978] = 25'b1111111111110110001111100;
    rom[58979] = 25'b1111111111110110001111111;
    rom[58980] = 25'b1111111111110110010000010;
    rom[58981] = 25'b1111111111110110010000101;
    rom[58982] = 25'b1111111111110110010001000;
    rom[58983] = 25'b1111111111110110010001011;
    rom[58984] = 25'b1111111111110110010001110;
    rom[58985] = 25'b1111111111110110010010001;
    rom[58986] = 25'b1111111111110110010010100;
    rom[58987] = 25'b1111111111110110010011000;
    rom[58988] = 25'b1111111111110110010011011;
    rom[58989] = 25'b1111111111110110010011110;
    rom[58990] = 25'b1111111111110110010100001;
    rom[58991] = 25'b1111111111110110010100100;
    rom[58992] = 25'b1111111111110110010100111;
    rom[58993] = 25'b1111111111110110010101010;
    rom[58994] = 25'b1111111111110110010101101;
    rom[58995] = 25'b1111111111110110010110000;
    rom[58996] = 25'b1111111111110110010110011;
    rom[58997] = 25'b1111111111110110010110110;
    rom[58998] = 25'b1111111111110110010111010;
    rom[58999] = 25'b1111111111110110010111101;
    rom[59000] = 25'b1111111111110110011000000;
    rom[59001] = 25'b1111111111110110011000011;
    rom[59002] = 25'b1111111111110110011000110;
    rom[59003] = 25'b1111111111110110011001001;
    rom[59004] = 25'b1111111111110110011001100;
    rom[59005] = 25'b1111111111110110011001111;
    rom[59006] = 25'b1111111111110110011010010;
    rom[59007] = 25'b1111111111110110011010101;
    rom[59008] = 25'b1111111111110110011011000;
    rom[59009] = 25'b1111111111110110011011100;
    rom[59010] = 25'b1111111111110110011011111;
    rom[59011] = 25'b1111111111110110011100010;
    rom[59012] = 25'b1111111111110110011100101;
    rom[59013] = 25'b1111111111110110011101000;
    rom[59014] = 25'b1111111111110110011101100;
    rom[59015] = 25'b1111111111110110011101111;
    rom[59016] = 25'b1111111111110110011110010;
    rom[59017] = 25'b1111111111110110011110101;
    rom[59018] = 25'b1111111111110110011111000;
    rom[59019] = 25'b1111111111110110011111011;
    rom[59020] = 25'b1111111111110110011111110;
    rom[59021] = 25'b1111111111110110100000001;
    rom[59022] = 25'b1111111111110110100000101;
    rom[59023] = 25'b1111111111110110100001000;
    rom[59024] = 25'b1111111111110110100001011;
    rom[59025] = 25'b1111111111110110100001111;
    rom[59026] = 25'b1111111111110110100010010;
    rom[59027] = 25'b1111111111110110100010101;
    rom[59028] = 25'b1111111111110110100011001;
    rom[59029] = 25'b1111111111110110100011100;
    rom[59030] = 25'b1111111111110110100011111;
    rom[59031] = 25'b1111111111110110100100010;
    rom[59032] = 25'b1111111111110110100100101;
    rom[59033] = 25'b1111111111110110100101000;
    rom[59034] = 25'b1111111111110110100101100;
    rom[59035] = 25'b1111111111110110100101111;
    rom[59036] = 25'b1111111111110110100110010;
    rom[59037] = 25'b1111111111110110100110110;
    rom[59038] = 25'b1111111111110110100111001;
    rom[59039] = 25'b1111111111110110100111100;
    rom[59040] = 25'b1111111111110110100111111;
    rom[59041] = 25'b1111111111110110101000010;
    rom[59042] = 25'b1111111111110110101000110;
    rom[59043] = 25'b1111111111110110101001001;
    rom[59044] = 25'b1111111111110110101001101;
    rom[59045] = 25'b1111111111110110101010000;
    rom[59046] = 25'b1111111111110110101010100;
    rom[59047] = 25'b1111111111110110101010111;
    rom[59048] = 25'b1111111111110110101011010;
    rom[59049] = 25'b1111111111110110101011101;
    rom[59050] = 25'b1111111111110110101100000;
    rom[59051] = 25'b1111111111110110101100100;
    rom[59052] = 25'b1111111111110110101100111;
    rom[59053] = 25'b1111111111110110101101011;
    rom[59054] = 25'b1111111111110110101101110;
    rom[59055] = 25'b1111111111110110101110001;
    rom[59056] = 25'b1111111111110110101110100;
    rom[59057] = 25'b1111111111110110101111000;
    rom[59058] = 25'b1111111111110110101111011;
    rom[59059] = 25'b1111111111110110101111111;
    rom[59060] = 25'b1111111111110110110000010;
    rom[59061] = 25'b1111111111110110110000110;
    rom[59062] = 25'b1111111111110110110001001;
    rom[59063] = 25'b1111111111110110110001100;
    rom[59064] = 25'b1111111111110110110001111;
    rom[59065] = 25'b1111111111110110110010011;
    rom[59066] = 25'b1111111111110110110010111;
    rom[59067] = 25'b1111111111110110110011010;
    rom[59068] = 25'b1111111111110110110011110;
    rom[59069] = 25'b1111111111110110110100001;
    rom[59070] = 25'b1111111111110110110100100;
    rom[59071] = 25'b1111111111110110110100111;
    rom[59072] = 25'b1111111111110110110101011;
    rom[59073] = 25'b1111111111110110110101111;
    rom[59074] = 25'b1111111111110110110110010;
    rom[59075] = 25'b1111111111110110110110101;
    rom[59076] = 25'b1111111111110110110111000;
    rom[59077] = 25'b1111111111110110110111100;
    rom[59078] = 25'b1111111111110110111000000;
    rom[59079] = 25'b1111111111110110111000011;
    rom[59080] = 25'b1111111111110110111000111;
    rom[59081] = 25'b1111111111110110111001010;
    rom[59082] = 25'b1111111111110110111001101;
    rom[59083] = 25'b1111111111110110111010001;
    rom[59084] = 25'b1111111111110110111010100;
    rom[59085] = 25'b1111111111110110111011000;
    rom[59086] = 25'b1111111111110110111011100;
    rom[59087] = 25'b1111111111110110111011111;
    rom[59088] = 25'b1111111111110110111100010;
    rom[59089] = 25'b1111111111110110111100110;
    rom[59090] = 25'b1111111111110110111101010;
    rom[59091] = 25'b1111111111110110111101101;
    rom[59092] = 25'b1111111111110110111110000;
    rom[59093] = 25'b1111111111110110111110100;
    rom[59094] = 25'b1111111111110110111110111;
    rom[59095] = 25'b1111111111110110111111011;
    rom[59096] = 25'b1111111111110110111111111;
    rom[59097] = 25'b1111111111110111000000010;
    rom[59098] = 25'b1111111111110111000000101;
    rom[59099] = 25'b1111111111110111000001001;
    rom[59100] = 25'b1111111111110111000001101;
    rom[59101] = 25'b1111111111110111000010001;
    rom[59102] = 25'b1111111111110111000010100;
    rom[59103] = 25'b1111111111110111000010111;
    rom[59104] = 25'b1111111111110111000011011;
    rom[59105] = 25'b1111111111110111000011111;
    rom[59106] = 25'b1111111111110111000100010;
    rom[59107] = 25'b1111111111110111000100110;
    rom[59108] = 25'b1111111111110111000101001;
    rom[59109] = 25'b1111111111110111000101101;
    rom[59110] = 25'b1111111111110111000110001;
    rom[59111] = 25'b1111111111110111000110100;
    rom[59112] = 25'b1111111111110111000110111;
    rom[59113] = 25'b1111111111110111000111011;
    rom[59114] = 25'b1111111111110111000111111;
    rom[59115] = 25'b1111111111110111001000011;
    rom[59116] = 25'b1111111111110111001000110;
    rom[59117] = 25'b1111111111110111001001001;
    rom[59118] = 25'b1111111111110111001001101;
    rom[59119] = 25'b1111111111110111001010001;
    rom[59120] = 25'b1111111111110111001010101;
    rom[59121] = 25'b1111111111110111001011000;
    rom[59122] = 25'b1111111111110111001011100;
    rom[59123] = 25'b1111111111110111001011111;
    rom[59124] = 25'b1111111111110111001100011;
    rom[59125] = 25'b1111111111110111001100111;
    rom[59126] = 25'b1111111111110111001101010;
    rom[59127] = 25'b1111111111110111001101110;
    rom[59128] = 25'b1111111111110111001110010;
    rom[59129] = 25'b1111111111110111001110101;
    rom[59130] = 25'b1111111111110111001111001;
    rom[59131] = 25'b1111111111110111001111101;
    rom[59132] = 25'b1111111111110111010000000;
    rom[59133] = 25'b1111111111110111010000100;
    rom[59134] = 25'b1111111111110111010000111;
    rom[59135] = 25'b1111111111110111010001011;
    rom[59136] = 25'b1111111111110111010001111;
    rom[59137] = 25'b1111111111110111010010011;
    rom[59138] = 25'b1111111111110111010010110;
    rom[59139] = 25'b1111111111110111010011010;
    rom[59140] = 25'b1111111111110111010011110;
    rom[59141] = 25'b1111111111110111010100010;
    rom[59142] = 25'b1111111111110111010100101;
    rom[59143] = 25'b1111111111110111010101001;
    rom[59144] = 25'b1111111111110111010101101;
    rom[59145] = 25'b1111111111110111010110000;
    rom[59146] = 25'b1111111111110111010110100;
    rom[59147] = 25'b1111111111110111010111000;
    rom[59148] = 25'b1111111111110111010111100;
    rom[59149] = 25'b1111111111110111010111111;
    rom[59150] = 25'b1111111111110111011000011;
    rom[59151] = 25'b1111111111110111011000111;
    rom[59152] = 25'b1111111111110111011001011;
    rom[59153] = 25'b1111111111110111011001110;
    rom[59154] = 25'b1111111111110111011010010;
    rom[59155] = 25'b1111111111110111011010110;
    rom[59156] = 25'b1111111111110111011011010;
    rom[59157] = 25'b1111111111110111011011101;
    rom[59158] = 25'b1111111111110111011100001;
    rom[59159] = 25'b1111111111110111011100101;
    rom[59160] = 25'b1111111111110111011101001;
    rom[59161] = 25'b1111111111110111011101100;
    rom[59162] = 25'b1111111111110111011110000;
    rom[59163] = 25'b1111111111110111011110100;
    rom[59164] = 25'b1111111111110111011110111;
    rom[59165] = 25'b1111111111110111011111011;
    rom[59166] = 25'b1111111111110111100000000;
    rom[59167] = 25'b1111111111110111100000011;
    rom[59168] = 25'b1111111111110111100000111;
    rom[59169] = 25'b1111111111110111100001011;
    rom[59170] = 25'b1111111111110111100001111;
    rom[59171] = 25'b1111111111110111100010010;
    rom[59172] = 25'b1111111111110111100010110;
    rom[59173] = 25'b1111111111110111100011010;
    rom[59174] = 25'b1111111111110111100011110;
    rom[59175] = 25'b1111111111110111100100001;
    rom[59176] = 25'b1111111111110111100100110;
    rom[59177] = 25'b1111111111110111100101010;
    rom[59178] = 25'b1111111111110111100101101;
    rom[59179] = 25'b1111111111110111100110001;
    rom[59180] = 25'b1111111111110111100110101;
    rom[59181] = 25'b1111111111110111100111000;
    rom[59182] = 25'b1111111111110111100111100;
    rom[59183] = 25'b1111111111110111101000001;
    rom[59184] = 25'b1111111111110111101000100;
    rom[59185] = 25'b1111111111110111101001000;
    rom[59186] = 25'b1111111111110111101001100;
    rom[59187] = 25'b1111111111110111101010000;
    rom[59188] = 25'b1111111111110111101010011;
    rom[59189] = 25'b1111111111110111101011000;
    rom[59190] = 25'b1111111111110111101011100;
    rom[59191] = 25'b1111111111110111101011111;
    rom[59192] = 25'b1111111111110111101100011;
    rom[59193] = 25'b1111111111110111101100111;
    rom[59194] = 25'b1111111111110111101101011;
    rom[59195] = 25'b1111111111110111101101111;
    rom[59196] = 25'b1111111111110111101110011;
    rom[59197] = 25'b1111111111110111101110110;
    rom[59198] = 25'b1111111111110111101111011;
    rom[59199] = 25'b1111111111110111101111111;
    rom[59200] = 25'b1111111111110111110000010;
    rom[59201] = 25'b1111111111110111110000110;
    rom[59202] = 25'b1111111111110111110001010;
    rom[59203] = 25'b1111111111110111110001110;
    rom[59204] = 25'b1111111111110111110010010;
    rom[59205] = 25'b1111111111110111110010110;
    rom[59206] = 25'b1111111111110111110011010;
    rom[59207] = 25'b1111111111110111110011110;
    rom[59208] = 25'b1111111111110111110100010;
    rom[59209] = 25'b1111111111110111110100110;
    rom[59210] = 25'b1111111111110111110101010;
    rom[59211] = 25'b1111111111110111110101110;
    rom[59212] = 25'b1111111111110111110110001;
    rom[59213] = 25'b1111111111110111110110101;
    rom[59214] = 25'b1111111111110111110111010;
    rom[59215] = 25'b1111111111110111110111101;
    rom[59216] = 25'b1111111111110111111000001;
    rom[59217] = 25'b1111111111110111111000110;
    rom[59218] = 25'b1111111111110111111001001;
    rom[59219] = 25'b1111111111110111111001101;
    rom[59220] = 25'b1111111111110111111010010;
    rom[59221] = 25'b1111111111110111111010101;
    rom[59222] = 25'b1111111111110111111011001;
    rom[59223] = 25'b1111111111110111111011110;
    rom[59224] = 25'b1111111111110111111100001;
    rom[59225] = 25'b1111111111110111111100101;
    rom[59226] = 25'b1111111111110111111101010;
    rom[59227] = 25'b1111111111110111111101101;
    rom[59228] = 25'b1111111111110111111110001;
    rom[59229] = 25'b1111111111110111111110101;
    rom[59230] = 25'b1111111111110111111111001;
    rom[59231] = 25'b1111111111110111111111101;
    rom[59232] = 25'b1111111111111000000000001;
    rom[59233] = 25'b1111111111111000000000101;
    rom[59234] = 25'b1111111111111000000001010;
    rom[59235] = 25'b1111111111111000000001101;
    rom[59236] = 25'b1111111111111000000010001;
    rom[59237] = 25'b1111111111111000000010110;
    rom[59238] = 25'b1111111111111000000011001;
    rom[59239] = 25'b1111111111111000000011101;
    rom[59240] = 25'b1111111111111000000100010;
    rom[59241] = 25'b1111111111111000000100101;
    rom[59242] = 25'b1111111111111000000101010;
    rom[59243] = 25'b1111111111111000000101101;
    rom[59244] = 25'b1111111111111000000110001;
    rom[59245] = 25'b1111111111111000000110110;
    rom[59246] = 25'b1111111111111000000111001;
    rom[59247] = 25'b1111111111111000000111110;
    rom[59248] = 25'b1111111111111000001000010;
    rom[59249] = 25'b1111111111111000001000110;
    rom[59250] = 25'b1111111111111000001001010;
    rom[59251] = 25'b1111111111111000001001110;
    rom[59252] = 25'b1111111111111000001010010;
    rom[59253] = 25'b1111111111111000001010110;
    rom[59254] = 25'b1111111111111000001011010;
    rom[59255] = 25'b1111111111111000001011110;
    rom[59256] = 25'b1111111111111000001100011;
    rom[59257] = 25'b1111111111111000001100110;
    rom[59258] = 25'b1111111111111000001101011;
    rom[59259] = 25'b1111111111111000001101110;
    rom[59260] = 25'b1111111111111000001110011;
    rom[59261] = 25'b1111111111111000001110111;
    rom[59262] = 25'b1111111111111000001111011;
    rom[59263] = 25'b1111111111111000001111111;
    rom[59264] = 25'b1111111111111000010000011;
    rom[59265] = 25'b1111111111111000010000111;
    rom[59266] = 25'b1111111111111000010001100;
    rom[59267] = 25'b1111111111111000010001111;
    rom[59268] = 25'b1111111111111000010010100;
    rom[59269] = 25'b1111111111111000010011000;
    rom[59270] = 25'b1111111111111000010011100;
    rom[59271] = 25'b1111111111111000010100000;
    rom[59272] = 25'b1111111111111000010100100;
    rom[59273] = 25'b1111111111111000010101000;
    rom[59274] = 25'b1111111111111000010101100;
    rom[59275] = 25'b1111111111111000010110000;
    rom[59276] = 25'b1111111111111000010110101;
    rom[59277] = 25'b1111111111111000010111000;
    rom[59278] = 25'b1111111111111000010111101;
    rom[59279] = 25'b1111111111111000011000001;
    rom[59280] = 25'b1111111111111000011000101;
    rom[59281] = 25'b1111111111111000011001001;
    rom[59282] = 25'b1111111111111000011001101;
    rom[59283] = 25'b1111111111111000011010010;
    rom[59284] = 25'b1111111111111000011010110;
    rom[59285] = 25'b1111111111111000011011010;
    rom[59286] = 25'b1111111111111000011011110;
    rom[59287] = 25'b1111111111111000011100010;
    rom[59288] = 25'b1111111111111000011100110;
    rom[59289] = 25'b1111111111111000011101011;
    rom[59290] = 25'b1111111111111000011101111;
    rom[59291] = 25'b1111111111111000011110011;
    rom[59292] = 25'b1111111111111000011110111;
    rom[59293] = 25'b1111111111111000011111011;
    rom[59294] = 25'b1111111111111000011111111;
    rom[59295] = 25'b1111111111111000100000011;
    rom[59296] = 25'b1111111111111000100001000;
    rom[59297] = 25'b1111111111111000100001100;
    rom[59298] = 25'b1111111111111000100010000;
    rom[59299] = 25'b1111111111111000100010100;
    rom[59300] = 25'b1111111111111000100011001;
    rom[59301] = 25'b1111111111111000100011101;
    rom[59302] = 25'b1111111111111000100100001;
    rom[59303] = 25'b1111111111111000100100101;
    rom[59304] = 25'b1111111111111000100101001;
    rom[59305] = 25'b1111111111111000100101110;
    rom[59306] = 25'b1111111111111000100110001;
    rom[59307] = 25'b1111111111111000100110110;
    rom[59308] = 25'b1111111111111000100111010;
    rom[59309] = 25'b1111111111111000100111110;
    rom[59310] = 25'b1111111111111000101000011;
    rom[59311] = 25'b1111111111111000101000110;
    rom[59312] = 25'b1111111111111000101001011;
    rom[59313] = 25'b1111111111111000101001111;
    rom[59314] = 25'b1111111111111000101010011;
    rom[59315] = 25'b1111111111111000101011000;
    rom[59316] = 25'b1111111111111000101011100;
    rom[59317] = 25'b1111111111111000101100000;
    rom[59318] = 25'b1111111111111000101100100;
    rom[59319] = 25'b1111111111111000101101001;
    rom[59320] = 25'b1111111111111000101101101;
    rom[59321] = 25'b1111111111111000101110001;
    rom[59322] = 25'b1111111111111000101110101;
    rom[59323] = 25'b1111111111111000101111001;
    rom[59324] = 25'b1111111111111000101111110;
    rom[59325] = 25'b1111111111111000110000010;
    rom[59326] = 25'b1111111111111000110000111;
    rom[59327] = 25'b1111111111111000110001010;
    rom[59328] = 25'b1111111111111000110001111;
    rom[59329] = 25'b1111111111111000110010011;
    rom[59330] = 25'b1111111111111000110010111;
    rom[59331] = 25'b1111111111111000110011100;
    rom[59332] = 25'b1111111111111000110100000;
    rom[59333] = 25'b1111111111111000110100101;
    rom[59334] = 25'b1111111111111000110101000;
    rom[59335] = 25'b1111111111111000110101101;
    rom[59336] = 25'b1111111111111000110110001;
    rom[59337] = 25'b1111111111111000110110101;
    rom[59338] = 25'b1111111111111000110111001;
    rom[59339] = 25'b1111111111111000110111110;
    rom[59340] = 25'b1111111111111000111000010;
    rom[59341] = 25'b1111111111111000111000110;
    rom[59342] = 25'b1111111111111000111001011;
    rom[59343] = 25'b1111111111111000111001111;
    rom[59344] = 25'b1111111111111000111010100;
    rom[59345] = 25'b1111111111111000111010111;
    rom[59346] = 25'b1111111111111000111011100;
    rom[59347] = 25'b1111111111111000111100000;
    rom[59348] = 25'b1111111111111000111100101;
    rom[59349] = 25'b1111111111111000111101001;
    rom[59350] = 25'b1111111111111000111101101;
    rom[59351] = 25'b1111111111111000111110001;
    rom[59352] = 25'b1111111111111000111110110;
    rom[59353] = 25'b1111111111111000111111010;
    rom[59354] = 25'b1111111111111000111111110;
    rom[59355] = 25'b1111111111111001000000011;
    rom[59356] = 25'b1111111111111001000000111;
    rom[59357] = 25'b1111111111111001000001011;
    rom[59358] = 25'b1111111111111001000001111;
    rom[59359] = 25'b1111111111111001000010100;
    rom[59360] = 25'b1111111111111001000011000;
    rom[59361] = 25'b1111111111111001000011101;
    rom[59362] = 25'b1111111111111001000100001;
    rom[59363] = 25'b1111111111111001000100101;
    rom[59364] = 25'b1111111111111001000101010;
    rom[59365] = 25'b1111111111111001000101110;
    rom[59366] = 25'b1111111111111001000110010;
    rom[59367] = 25'b1111111111111001000110110;
    rom[59368] = 25'b1111111111111001000111011;
    rom[59369] = 25'b1111111111111001000111111;
    rom[59370] = 25'b1111111111111001001000100;
    rom[59371] = 25'b1111111111111001001001000;
    rom[59372] = 25'b1111111111111001001001100;
    rom[59373] = 25'b1111111111111001001010000;
    rom[59374] = 25'b1111111111111001001010101;
    rom[59375] = 25'b1111111111111001001011001;
    rom[59376] = 25'b1111111111111001001011110;
    rom[59377] = 25'b1111111111111001001100010;
    rom[59378] = 25'b1111111111111001001100110;
    rom[59379] = 25'b1111111111111001001101011;
    rom[59380] = 25'b1111111111111001001101111;
    rom[59381] = 25'b1111111111111001001110011;
    rom[59382] = 25'b1111111111111001001111000;
    rom[59383] = 25'b1111111111111001001111100;
    rom[59384] = 25'b1111111111111001010000000;
    rom[59385] = 25'b1111111111111001010000101;
    rom[59386] = 25'b1111111111111001010001001;
    rom[59387] = 25'b1111111111111001010001110;
    rom[59388] = 25'b1111111111111001010010010;
    rom[59389] = 25'b1111111111111001010010111;
    rom[59390] = 25'b1111111111111001010011011;
    rom[59391] = 25'b1111111111111001010011111;
    rom[59392] = 25'b1111111111111001010100011;
    rom[59393] = 25'b1111111111111001010101000;
    rom[59394] = 25'b1111111111111001010101100;
    rom[59395] = 25'b1111111111111001010110001;
    rom[59396] = 25'b1111111111111001010110101;
    rom[59397] = 25'b1111111111111001010111010;
    rom[59398] = 25'b1111111111111001010111110;
    rom[59399] = 25'b1111111111111001011000010;
    rom[59400] = 25'b1111111111111001011000110;
    rom[59401] = 25'b1111111111111001011001011;
    rom[59402] = 25'b1111111111111001011001111;
    rom[59403] = 25'b1111111111111001011010100;
    rom[59404] = 25'b1111111111111001011011000;
    rom[59405] = 25'b1111111111111001011011101;
    rom[59406] = 25'b1111111111111001011100001;
    rom[59407] = 25'b1111111111111001011100110;
    rom[59408] = 25'b1111111111111001011101010;
    rom[59409] = 25'b1111111111111001011101110;
    rom[59410] = 25'b1111111111111001011110010;
    rom[59411] = 25'b1111111111111001011110111;
    rom[59412] = 25'b1111111111111001011111011;
    rom[59413] = 25'b1111111111111001100000000;
    rom[59414] = 25'b1111111111111001100000100;
    rom[59415] = 25'b1111111111111001100001001;
    rom[59416] = 25'b1111111111111001100001101;
    rom[59417] = 25'b1111111111111001100010010;
    rom[59418] = 25'b1111111111111001100010110;
    rom[59419] = 25'b1111111111111001100011011;
    rom[59420] = 25'b1111111111111001100011111;
    rom[59421] = 25'b1111111111111001100100011;
    rom[59422] = 25'b1111111111111001100101000;
    rom[59423] = 25'b1111111111111001100101100;
    rom[59424] = 25'b1111111111111001100110000;
    rom[59425] = 25'b1111111111111001100110101;
    rom[59426] = 25'b1111111111111001100111001;
    rom[59427] = 25'b1111111111111001100111110;
    rom[59428] = 25'b1111111111111001101000010;
    rom[59429] = 25'b1111111111111001101000111;
    rom[59430] = 25'b1111111111111001101001011;
    rom[59431] = 25'b1111111111111001101010000;
    rom[59432] = 25'b1111111111111001101010100;
    rom[59433] = 25'b1111111111111001101011001;
    rom[59434] = 25'b1111111111111001101011101;
    rom[59435] = 25'b1111111111111001101100010;
    rom[59436] = 25'b1111111111111001101100110;
    rom[59437] = 25'b1111111111111001101101010;
    rom[59438] = 25'b1111111111111001101101111;
    rom[59439] = 25'b1111111111111001101110011;
    rom[59440] = 25'b1111111111111001101110111;
    rom[59441] = 25'b1111111111111001101111100;
    rom[59442] = 25'b1111111111111001110000000;
    rom[59443] = 25'b1111111111111001110000101;
    rom[59444] = 25'b1111111111111001110001001;
    rom[59445] = 25'b1111111111111001110001110;
    rom[59446] = 25'b1111111111111001110010010;
    rom[59447] = 25'b1111111111111001110010111;
    rom[59448] = 25'b1111111111111001110011011;
    rom[59449] = 25'b1111111111111001110100000;
    rom[59450] = 25'b1111111111111001110100100;
    rom[59451] = 25'b1111111111111001110101001;
    rom[59452] = 25'b1111111111111001110101101;
    rom[59453] = 25'b1111111111111001110110010;
    rom[59454] = 25'b1111111111111001110110110;
    rom[59455] = 25'b1111111111111001110111011;
    rom[59456] = 25'b1111111111111001110111111;
    rom[59457] = 25'b1111111111111001111000100;
    rom[59458] = 25'b1111111111111001111001000;
    rom[59459] = 25'b1111111111111001111001101;
    rom[59460] = 25'b1111111111111001111010001;
    rom[59461] = 25'b1111111111111001111010110;
    rom[59462] = 25'b1111111111111001111011010;
    rom[59463] = 25'b1111111111111001111011111;
    rom[59464] = 25'b1111111111111001111100011;
    rom[59465] = 25'b1111111111111001111101000;
    rom[59466] = 25'b1111111111111001111101100;
    rom[59467] = 25'b1111111111111001111110000;
    rom[59468] = 25'b1111111111111001111110101;
    rom[59469] = 25'b1111111111111001111111001;
    rom[59470] = 25'b1111111111111001111111110;
    rom[59471] = 25'b1111111111111010000000010;
    rom[59472] = 25'b1111111111111010000000111;
    rom[59473] = 25'b1111111111111010000001011;
    rom[59474] = 25'b1111111111111010000010000;
    rom[59475] = 25'b1111111111111010000010100;
    rom[59476] = 25'b1111111111111010000011001;
    rom[59477] = 25'b1111111111111010000011101;
    rom[59478] = 25'b1111111111111010000100010;
    rom[59479] = 25'b1111111111111010000100110;
    rom[59480] = 25'b1111111111111010000101011;
    rom[59481] = 25'b1111111111111010000101111;
    rom[59482] = 25'b1111111111111010000110100;
    rom[59483] = 25'b1111111111111010000111000;
    rom[59484] = 25'b1111111111111010000111101;
    rom[59485] = 25'b1111111111111010001000001;
    rom[59486] = 25'b1111111111111010001000110;
    rom[59487] = 25'b1111111111111010001001010;
    rom[59488] = 25'b1111111111111010001001111;
    rom[59489] = 25'b1111111111111010001010011;
    rom[59490] = 25'b1111111111111010001011000;
    rom[59491] = 25'b1111111111111010001011100;
    rom[59492] = 25'b1111111111111010001100001;
    rom[59493] = 25'b1111111111111010001100110;
    rom[59494] = 25'b1111111111111010001101010;
    rom[59495] = 25'b1111111111111010001101111;
    rom[59496] = 25'b1111111111111010001110011;
    rom[59497] = 25'b1111111111111010001111000;
    rom[59498] = 25'b1111111111111010001111100;
    rom[59499] = 25'b1111111111111010010000001;
    rom[59500] = 25'b1111111111111010010000101;
    rom[59501] = 25'b1111111111111010010001010;
    rom[59502] = 25'b1111111111111010010001110;
    rom[59503] = 25'b1111111111111010010010011;
    rom[59504] = 25'b1111111111111010010010111;
    rom[59505] = 25'b1111111111111010010011100;
    rom[59506] = 25'b1111111111111010010100000;
    rom[59507] = 25'b1111111111111010010100101;
    rom[59508] = 25'b1111111111111010010101001;
    rom[59509] = 25'b1111111111111010010101110;
    rom[59510] = 25'b1111111111111010010110010;
    rom[59511] = 25'b1111111111111010010110110;
    rom[59512] = 25'b1111111111111010010111100;
    rom[59513] = 25'b1111111111111010011000000;
    rom[59514] = 25'b1111111111111010011000101;
    rom[59515] = 25'b1111111111111010011001001;
    rom[59516] = 25'b1111111111111010011001110;
    rom[59517] = 25'b1111111111111010011010010;
    rom[59518] = 25'b1111111111111010011010111;
    rom[59519] = 25'b1111111111111010011011011;
    rom[59520] = 25'b1111111111111010011100000;
    rom[59521] = 25'b1111111111111010011100100;
    rom[59522] = 25'b1111111111111010011101001;
    rom[59523] = 25'b1111111111111010011101101;
    rom[59524] = 25'b1111111111111010011110001;
    rom[59525] = 25'b1111111111111010011110110;
    rom[59526] = 25'b1111111111111010011111011;
    rom[59527] = 25'b1111111111111010100000000;
    rom[59528] = 25'b1111111111111010100000100;
    rom[59529] = 25'b1111111111111010100001001;
    rom[59530] = 25'b1111111111111010100001101;
    rom[59531] = 25'b1111111111111010100010010;
    rom[59532] = 25'b1111111111111010100010110;
    rom[59533] = 25'b1111111111111010100011011;
    rom[59534] = 25'b1111111111111010100011111;
    rom[59535] = 25'b1111111111111010100100100;
    rom[59536] = 25'b1111111111111010100101000;
    rom[59537] = 25'b1111111111111010100101101;
    rom[59538] = 25'b1111111111111010100110001;
    rom[59539] = 25'b1111111111111010100110110;
    rom[59540] = 25'b1111111111111010100111011;
    rom[59541] = 25'b1111111111111010100111111;
    rom[59542] = 25'b1111111111111010101000100;
    rom[59543] = 25'b1111111111111010101001000;
    rom[59544] = 25'b1111111111111010101001101;
    rom[59545] = 25'b1111111111111010101010001;
    rom[59546] = 25'b1111111111111010101010110;
    rom[59547] = 25'b1111111111111010101011010;
    rom[59548] = 25'b1111111111111010101011111;
    rom[59549] = 25'b1111111111111010101100011;
    rom[59550] = 25'b1111111111111010101101000;
    rom[59551] = 25'b1111111111111010101101101;
    rom[59552] = 25'b1111111111111010101110001;
    rom[59553] = 25'b1111111111111010101110110;
    rom[59554] = 25'b1111111111111010101111010;
    rom[59555] = 25'b1111111111111010101111111;
    rom[59556] = 25'b1111111111111010110000011;
    rom[59557] = 25'b1111111111111010110001000;
    rom[59558] = 25'b1111111111111010110001100;
    rom[59559] = 25'b1111111111111010110010001;
    rom[59560] = 25'b1111111111111010110010110;
    rom[59561] = 25'b1111111111111010110011010;
    rom[59562] = 25'b1111111111111010110011111;
    rom[59563] = 25'b1111111111111010110100011;
    rom[59564] = 25'b1111111111111010110101000;
    rom[59565] = 25'b1111111111111010110101100;
    rom[59566] = 25'b1111111111111010110110001;
    rom[59567] = 25'b1111111111111010110110101;
    rom[59568] = 25'b1111111111111010110111010;
    rom[59569] = 25'b1111111111111010110111110;
    rom[59570] = 25'b1111111111111010111000011;
    rom[59571] = 25'b1111111111111010111001000;
    rom[59572] = 25'b1111111111111010111001100;
    rom[59573] = 25'b1111111111111010111010001;
    rom[59574] = 25'b1111111111111010111010101;
    rom[59575] = 25'b1111111111111010111011010;
    rom[59576] = 25'b1111111111111010111011110;
    rom[59577] = 25'b1111111111111010111100011;
    rom[59578] = 25'b1111111111111010111100111;
    rom[59579] = 25'b1111111111111010111101101;
    rom[59580] = 25'b1111111111111010111110001;
    rom[59581] = 25'b1111111111111010111110101;
    rom[59582] = 25'b1111111111111010111111010;
    rom[59583] = 25'b1111111111111010111111110;
    rom[59584] = 25'b1111111111111011000000011;
    rom[59585] = 25'b1111111111111011000000111;
    rom[59586] = 25'b1111111111111011000001100;
    rom[59587] = 25'b1111111111111011000010000;
    rom[59588] = 25'b1111111111111011000010110;
    rom[59589] = 25'b1111111111111011000011010;
    rom[59590] = 25'b1111111111111011000011111;
    rom[59591] = 25'b1111111111111011000100011;
    rom[59592] = 25'b1111111111111011000101000;
    rom[59593] = 25'b1111111111111011000101100;
    rom[59594] = 25'b1111111111111011000110001;
    rom[59595] = 25'b1111111111111011000110101;
    rom[59596] = 25'b1111111111111011000111001;
    rom[59597] = 25'b1111111111111011000111111;
    rom[59598] = 25'b1111111111111011001000011;
    rom[59599] = 25'b1111111111111011001001000;
    rom[59600] = 25'b1111111111111011001001100;
    rom[59601] = 25'b1111111111111011001010001;
    rom[59602] = 25'b1111111111111011001010101;
    rom[59603] = 25'b1111111111111011001011010;
    rom[59604] = 25'b1111111111111011001011110;
    rom[59605] = 25'b1111111111111011001100011;
    rom[59606] = 25'b1111111111111011001101000;
    rom[59607] = 25'b1111111111111011001101100;
    rom[59608] = 25'b1111111111111011001110001;
    rom[59609] = 25'b1111111111111011001110101;
    rom[59610] = 25'b1111111111111011001111010;
    rom[59611] = 25'b1111111111111011001111110;
    rom[59612] = 25'b1111111111111011010000011;
    rom[59613] = 25'b1111111111111011010000111;
    rom[59614] = 25'b1111111111111011010001100;
    rom[59615] = 25'b1111111111111011010010001;
    rom[59616] = 25'b1111111111111011010010101;
    rom[59617] = 25'b1111111111111011010011010;
    rom[59618] = 25'b1111111111111011010011110;
    rom[59619] = 25'b1111111111111011010100011;
    rom[59620] = 25'b1111111111111011010100111;
    rom[59621] = 25'b1111111111111011010101100;
    rom[59622] = 25'b1111111111111011010110000;
    rom[59623] = 25'b1111111111111011010110101;
    rom[59624] = 25'b1111111111111011010111010;
    rom[59625] = 25'b1111111111111011010111110;
    rom[59626] = 25'b1111111111111011011000011;
    rom[59627] = 25'b1111111111111011011000111;
    rom[59628] = 25'b1111111111111011011001100;
    rom[59629] = 25'b1111111111111011011010000;
    rom[59630] = 25'b1111111111111011011010101;
    rom[59631] = 25'b1111111111111011011011001;
    rom[59632] = 25'b1111111111111011011011111;
    rom[59633] = 25'b1111111111111011011100011;
    rom[59634] = 25'b1111111111111011011101000;
    rom[59635] = 25'b1111111111111011011101100;
    rom[59636] = 25'b1111111111111011011110001;
    rom[59637] = 25'b1111111111111011011110101;
    rom[59638] = 25'b1111111111111011011111001;
    rom[59639] = 25'b1111111111111011011111110;
    rom[59640] = 25'b1111111111111011100000011;
    rom[59641] = 25'b1111111111111011100001000;
    rom[59642] = 25'b1111111111111011100001100;
    rom[59643] = 25'b1111111111111011100010001;
    rom[59644] = 25'b1111111111111011100010101;
    rom[59645] = 25'b1111111111111011100011010;
    rom[59646] = 25'b1111111111111011100011110;
    rom[59647] = 25'b1111111111111011100100011;
    rom[59648] = 25'b1111111111111011100100111;
    rom[59649] = 25'b1111111111111011100101100;
    rom[59650] = 25'b1111111111111011100110001;
    rom[59651] = 25'b1111111111111011100110101;
    rom[59652] = 25'b1111111111111011100111010;
    rom[59653] = 25'b1111111111111011100111110;
    rom[59654] = 25'b1111111111111011101000011;
    rom[59655] = 25'b1111111111111011101000111;
    rom[59656] = 25'b1111111111111011101001100;
    rom[59657] = 25'b1111111111111011101010000;
    rom[59658] = 25'b1111111111111011101010101;
    rom[59659] = 25'b1111111111111011101011010;
    rom[59660] = 25'b1111111111111011101011110;
    rom[59661] = 25'b1111111111111011101100011;
    rom[59662] = 25'b1111111111111011101100111;
    rom[59663] = 25'b1111111111111011101101100;
    rom[59664] = 25'b1111111111111011101110000;
    rom[59665] = 25'b1111111111111011101110101;
    rom[59666] = 25'b1111111111111011101111001;
    rom[59667] = 25'b1111111111111011101111110;
    rom[59668] = 25'b1111111111111011110000011;
    rom[59669] = 25'b1111111111111011110000111;
    rom[59670] = 25'b1111111111111011110001100;
    rom[59671] = 25'b1111111111111011110010000;
    rom[59672] = 25'b1111111111111011110010101;
    rom[59673] = 25'b1111111111111011110011001;
    rom[59674] = 25'b1111111111111011110011110;
    rom[59675] = 25'b1111111111111011110100010;
    rom[59676] = 25'b1111111111111011110100111;
    rom[59677] = 25'b1111111111111011110101100;
    rom[59678] = 25'b1111111111111011110110001;
    rom[59679] = 25'b1111111111111011110110101;
    rom[59680] = 25'b1111111111111011110111001;
    rom[59681] = 25'b1111111111111011110111110;
    rom[59682] = 25'b1111111111111011111000010;
    rom[59683] = 25'b1111111111111011111000111;
    rom[59684] = 25'b1111111111111011111001011;
    rom[59685] = 25'b1111111111111011111010000;
    rom[59686] = 25'b1111111111111011111010100;
    rom[59687] = 25'b1111111111111011111011010;
    rom[59688] = 25'b1111111111111011111011110;
    rom[59689] = 25'b1111111111111011111100011;
    rom[59690] = 25'b1111111111111011111100111;
    rom[59691] = 25'b1111111111111011111101100;
    rom[59692] = 25'b1111111111111011111110000;
    rom[59693] = 25'b1111111111111011111110101;
    rom[59694] = 25'b1111111111111011111111001;
    rom[59695] = 25'b1111111111111011111111101;
    rom[59696] = 25'b1111111111111100000000010;
    rom[59697] = 25'b1111111111111100000000111;
    rom[59698] = 25'b1111111111111100000001100;
    rom[59699] = 25'b1111111111111100000010000;
    rom[59700] = 25'b1111111111111100000010101;
    rom[59701] = 25'b1111111111111100000011001;
    rom[59702] = 25'b1111111111111100000011110;
    rom[59703] = 25'b1111111111111100000100010;
    rom[59704] = 25'b1111111111111100000100111;
    rom[59705] = 25'b1111111111111100000101011;
    rom[59706] = 25'b1111111111111100000110000;
    rom[59707] = 25'b1111111111111100000110100;
    rom[59708] = 25'b1111111111111100000111000;
    rom[59709] = 25'b1111111111111100000111110;
    rom[59710] = 25'b1111111111111100001000010;
    rom[59711] = 25'b1111111111111100001000111;
    rom[59712] = 25'b1111111111111100001001011;
    rom[59713] = 25'b1111111111111100001010000;
    rom[59714] = 25'b1111111111111100001010100;
    rom[59715] = 25'b1111111111111100001011001;
    rom[59716] = 25'b1111111111111100001011101;
    rom[59717] = 25'b1111111111111100001100010;
    rom[59718] = 25'b1111111111111100001100110;
    rom[59719] = 25'b1111111111111100001101011;
    rom[59720] = 25'b1111111111111100001101111;
    rom[59721] = 25'b1111111111111100001110100;
    rom[59722] = 25'b1111111111111100001111001;
    rom[59723] = 25'b1111111111111100001111101;
    rom[59724] = 25'b1111111111111100010000010;
    rom[59725] = 25'b1111111111111100010000110;
    rom[59726] = 25'b1111111111111100010001011;
    rom[59727] = 25'b1111111111111100010001111;
    rom[59728] = 25'b1111111111111100010010100;
    rom[59729] = 25'b1111111111111100010011000;
    rom[59730] = 25'b1111111111111100010011101;
    rom[59731] = 25'b1111111111111100010100001;
    rom[59732] = 25'b1111111111111100010100110;
    rom[59733] = 25'b1111111111111100010101010;
    rom[59734] = 25'b1111111111111100010101111;
    rom[59735] = 25'b1111111111111100010110011;
    rom[59736] = 25'b1111111111111100010110111;
    rom[59737] = 25'b1111111111111100010111100;
    rom[59738] = 25'b1111111111111100011000001;
    rom[59739] = 25'b1111111111111100011000110;
    rom[59740] = 25'b1111111111111100011001010;
    rom[59741] = 25'b1111111111111100011001111;
    rom[59742] = 25'b1111111111111100011010011;
    rom[59743] = 25'b1111111111111100011011000;
    rom[59744] = 25'b1111111111111100011011100;
    rom[59745] = 25'b1111111111111100011100001;
    rom[59746] = 25'b1111111111111100011100101;
    rom[59747] = 25'b1111111111111100011101010;
    rom[59748] = 25'b1111111111111100011101110;
    rom[59749] = 25'b1111111111111100011110011;
    rom[59750] = 25'b1111111111111100011110111;
    rom[59751] = 25'b1111111111111100011111011;
    rom[59752] = 25'b1111111111111100100000000;
    rom[59753] = 25'b1111111111111100100000100;
    rom[59754] = 25'b1111111111111100100001001;
    rom[59755] = 25'b1111111111111100100001101;
    rom[59756] = 25'b1111111111111100100010010;
    rom[59757] = 25'b1111111111111100100010110;
    rom[59758] = 25'b1111111111111100100011011;
    rom[59759] = 25'b1111111111111100100011111;
    rom[59760] = 25'b1111111111111100100100100;
    rom[59761] = 25'b1111111111111100100101000;
    rom[59762] = 25'b1111111111111100100101110;
    rom[59763] = 25'b1111111111111100100110010;
    rom[59764] = 25'b1111111111111100100110111;
    rom[59765] = 25'b1111111111111100100111011;
    rom[59766] = 25'b1111111111111100100111111;
    rom[59767] = 25'b1111111111111100101000100;
    rom[59768] = 25'b1111111111111100101001000;
    rom[59769] = 25'b1111111111111100101001101;
    rom[59770] = 25'b1111111111111100101010001;
    rom[59771] = 25'b1111111111111100101010110;
    rom[59772] = 25'b1111111111111100101011010;
    rom[59773] = 25'b1111111111111100101011111;
    rom[59774] = 25'b1111111111111100101100011;
    rom[59775] = 25'b1111111111111100101101000;
    rom[59776] = 25'b1111111111111100101101100;
    rom[59777] = 25'b1111111111111100101110001;
    rom[59778] = 25'b1111111111111100101110101;
    rom[59779] = 25'b1111111111111100101111010;
    rom[59780] = 25'b1111111111111100101111110;
    rom[59781] = 25'b1111111111111100110000011;
    rom[59782] = 25'b1111111111111100110000111;
    rom[59783] = 25'b1111111111111100110001100;
    rom[59784] = 25'b1111111111111100110010000;
    rom[59785] = 25'b1111111111111100110010101;
    rom[59786] = 25'b1111111111111100110011001;
    rom[59787] = 25'b1111111111111100110011110;
    rom[59788] = 25'b1111111111111100110100010;
    rom[59789] = 25'b1111111111111100110100111;
    rom[59790] = 25'b1111111111111100110101011;
    rom[59791] = 25'b1111111111111100110110000;
    rom[59792] = 25'b1111111111111100110110100;
    rom[59793] = 25'b1111111111111100110111000;
    rom[59794] = 25'b1111111111111100110111101;
    rom[59795] = 25'b1111111111111100111000001;
    rom[59796] = 25'b1111111111111100111000110;
    rom[59797] = 25'b1111111111111100111001010;
    rom[59798] = 25'b1111111111111100111001111;
    rom[59799] = 25'b1111111111111100111010011;
    rom[59800] = 25'b1111111111111100111011000;
    rom[59801] = 25'b1111111111111100111011100;
    rom[59802] = 25'b1111111111111100111100001;
    rom[59803] = 25'b1111111111111100111100101;
    rom[59804] = 25'b1111111111111100111101001;
    rom[59805] = 25'b1111111111111100111101110;
    rom[59806] = 25'b1111111111111100111110010;
    rom[59807] = 25'b1111111111111100111110111;
    rom[59808] = 25'b1111111111111100111111011;
    rom[59809] = 25'b1111111111111100111111111;
    rom[59810] = 25'b1111111111111101000000100;
    rom[59811] = 25'b1111111111111101000001000;
    rom[59812] = 25'b1111111111111101000001101;
    rom[59813] = 25'b1111111111111101000010001;
    rom[59814] = 25'b1111111111111101000010110;
    rom[59815] = 25'b1111111111111101000011010;
    rom[59816] = 25'b1111111111111101000011111;
    rom[59817] = 25'b1111111111111101000100011;
    rom[59818] = 25'b1111111111111101000101000;
    rom[59819] = 25'b1111111111111101000101100;
    rom[59820] = 25'b1111111111111101000110001;
    rom[59821] = 25'b1111111111111101000110101;
    rom[59822] = 25'b1111111111111101000111010;
    rom[59823] = 25'b1111111111111101000111110;
    rom[59824] = 25'b1111111111111101001000011;
    rom[59825] = 25'b1111111111111101001000110;
    rom[59826] = 25'b1111111111111101001001011;
    rom[59827] = 25'b1111111111111101001001111;
    rom[59828] = 25'b1111111111111101001010100;
    rom[59829] = 25'b1111111111111101001011000;
    rom[59830] = 25'b1111111111111101001011101;
    rom[59831] = 25'b1111111111111101001100001;
    rom[59832] = 25'b1111111111111101001100110;
    rom[59833] = 25'b1111111111111101001101010;
    rom[59834] = 25'b1111111111111101001101111;
    rom[59835] = 25'b1111111111111101001110011;
    rom[59836] = 25'b1111111111111101001111000;
    rom[59837] = 25'b1111111111111101001111100;
    rom[59838] = 25'b1111111111111101010000000;
    rom[59839] = 25'b1111111111111101010000100;
    rom[59840] = 25'b1111111111111101010001001;
    rom[59841] = 25'b1111111111111101010001101;
    rom[59842] = 25'b1111111111111101010010010;
    rom[59843] = 25'b1111111111111101010010110;
    rom[59844] = 25'b1111111111111101010011011;
    rom[59845] = 25'b1111111111111101010011111;
    rom[59846] = 25'b1111111111111101010100100;
    rom[59847] = 25'b1111111111111101010101000;
    rom[59848] = 25'b1111111111111101010101100;
    rom[59849] = 25'b1111111111111101010110001;
    rom[59850] = 25'b1111111111111101010110101;
    rom[59851] = 25'b1111111111111101010111001;
    rom[59852] = 25'b1111111111111101010111110;
    rom[59853] = 25'b1111111111111101011000010;
    rom[59854] = 25'b1111111111111101011000111;
    rom[59855] = 25'b1111111111111101011001011;
    rom[59856] = 25'b1111111111111101011010000;
    rom[59857] = 25'b1111111111111101011010100;
    rom[59858] = 25'b1111111111111101011011000;
    rom[59859] = 25'b1111111111111101011011101;
    rom[59860] = 25'b1111111111111101011100001;
    rom[59861] = 25'b1111111111111101011100110;
    rom[59862] = 25'b1111111111111101011101010;
    rom[59863] = 25'b1111111111111101011101111;
    rom[59864] = 25'b1111111111111101011110011;
    rom[59865] = 25'b1111111111111101011110111;
    rom[59866] = 25'b1111111111111101011111011;
    rom[59867] = 25'b1111111111111101100000000;
    rom[59868] = 25'b1111111111111101100000100;
    rom[59869] = 25'b1111111111111101100001001;
    rom[59870] = 25'b1111111111111101100001101;
    rom[59871] = 25'b1111111111111101100010010;
    rom[59872] = 25'b1111111111111101100010101;
    rom[59873] = 25'b1111111111111101100011010;
    rom[59874] = 25'b1111111111111101100011110;
    rom[59875] = 25'b1111111111111101100100011;
    rom[59876] = 25'b1111111111111101100100111;
    rom[59877] = 25'b1111111111111101100101100;
    rom[59878] = 25'b1111111111111101100110000;
    rom[59879] = 25'b1111111111111101100110100;
    rom[59880] = 25'b1111111111111101100111001;
    rom[59881] = 25'b1111111111111101100111101;
    rom[59882] = 25'b1111111111111101101000001;
    rom[59883] = 25'b1111111111111101101000110;
    rom[59884] = 25'b1111111111111101101001010;
    rom[59885] = 25'b1111111111111101101001110;
    rom[59886] = 25'b1111111111111101101010011;
    rom[59887] = 25'b1111111111111101101010111;
    rom[59888] = 25'b1111111111111101101011100;
    rom[59889] = 25'b1111111111111101101011111;
    rom[59890] = 25'b1111111111111101101100100;
    rom[59891] = 25'b1111111111111101101101000;
    rom[59892] = 25'b1111111111111101101101101;
    rom[59893] = 25'b1111111111111101101110001;
    rom[59894] = 25'b1111111111111101101110101;
    rom[59895] = 25'b1111111111111101101111010;
    rom[59896] = 25'b1111111111111101101111110;
    rom[59897] = 25'b1111111111111101110000010;
    rom[59898] = 25'b1111111111111101110000111;
    rom[59899] = 25'b1111111111111101110001011;
    rom[59900] = 25'b1111111111111101110001111;
    rom[59901] = 25'b1111111111111101110010100;
    rom[59902] = 25'b1111111111111101110011000;
    rom[59903] = 25'b1111111111111101110011101;
    rom[59904] = 25'b1111111111111101110100000;
    rom[59905] = 25'b1111111111111101110100101;
    rom[59906] = 25'b1111111111111101110101001;
    rom[59907] = 25'b1111111111111101110101110;
    rom[59908] = 25'b1111111111111101110110010;
    rom[59909] = 25'b1111111111111101110110110;
    rom[59910] = 25'b1111111111111101110111010;
    rom[59911] = 25'b1111111111111101110111111;
    rom[59912] = 25'b1111111111111101111000011;
    rom[59913] = 25'b1111111111111101111000111;
    rom[59914] = 25'b1111111111111101111001100;
    rom[59915] = 25'b1111111111111101111010000;
    rom[59916] = 25'b1111111111111101111010100;
    rom[59917] = 25'b1111111111111101111011000;
    rom[59918] = 25'b1111111111111101111011101;
    rom[59919] = 25'b1111111111111101111100001;
    rom[59920] = 25'b1111111111111101111100101;
    rom[59921] = 25'b1111111111111101111101010;
    rom[59922] = 25'b1111111111111101111101110;
    rom[59923] = 25'b1111111111111101111110011;
    rom[59924] = 25'b1111111111111101111110110;
    rom[59925] = 25'b1111111111111101111111011;
    rom[59926] = 25'b1111111111111101111111111;
    rom[59927] = 25'b1111111111111110000000011;
    rom[59928] = 25'b1111111111111110000000111;
    rom[59929] = 25'b1111111111111110000001100;
    rom[59930] = 25'b1111111111111110000010000;
    rom[59931] = 25'b1111111111111110000010100;
    rom[59932] = 25'b1111111111111110000011001;
    rom[59933] = 25'b1111111111111110000011101;
    rom[59934] = 25'b1111111111111110000100001;
    rom[59935] = 25'b1111111111111110000100101;
    rom[59936] = 25'b1111111111111110000101010;
    rom[59937] = 25'b1111111111111110000101110;
    rom[59938] = 25'b1111111111111110000110010;
    rom[59939] = 25'b1111111111111110000110111;
    rom[59940] = 25'b1111111111111110000111011;
    rom[59941] = 25'b1111111111111110000111111;
    rom[59942] = 25'b1111111111111110001000011;
    rom[59943] = 25'b1111111111111110001001000;
    rom[59944] = 25'b1111111111111110001001011;
    rom[59945] = 25'b1111111111111110001010000;
    rom[59946] = 25'b1111111111111110001010100;
    rom[59947] = 25'b1111111111111110001011000;
    rom[59948] = 25'b1111111111111110001011101;
    rom[59949] = 25'b1111111111111110001100001;
    rom[59950] = 25'b1111111111111110001100101;
    rom[59951] = 25'b1111111111111110001101001;
    rom[59952] = 25'b1111111111111110001101110;
    rom[59953] = 25'b1111111111111110001110010;
    rom[59954] = 25'b1111111111111110001110110;
    rom[59955] = 25'b1111111111111110001111011;
    rom[59956] = 25'b1111111111111110001111110;
    rom[59957] = 25'b1111111111111110010000011;
    rom[59958] = 25'b1111111111111110010000111;
    rom[59959] = 25'b1111111111111110010001011;
    rom[59960] = 25'b1111111111111110010001111;
    rom[59961] = 25'b1111111111111110010010100;
    rom[59962] = 25'b1111111111111110010011000;
    rom[59963] = 25'b1111111111111110010011100;
    rom[59964] = 25'b1111111111111110010100000;
    rom[59965] = 25'b1111111111111110010100100;
    rom[59966] = 25'b1111111111111110010101001;
    rom[59967] = 25'b1111111111111110010101101;
    rom[59968] = 25'b1111111111111110010110001;
    rom[59969] = 25'b1111111111111110010110101;
    rom[59970] = 25'b1111111111111110010111001;
    rom[59971] = 25'b1111111111111110010111110;
    rom[59972] = 25'b1111111111111110011000001;
    rom[59973] = 25'b1111111111111110011000110;
    rom[59974] = 25'b1111111111111110011001010;
    rom[59975] = 25'b1111111111111110011001110;
    rom[59976] = 25'b1111111111111110011010011;
    rom[59977] = 25'b1111111111111110011010110;
    rom[59978] = 25'b1111111111111110011011011;
    rom[59979] = 25'b1111111111111110011011111;
    rom[59980] = 25'b1111111111111110011100011;
    rom[59981] = 25'b1111111111111110011101000;
    rom[59982] = 25'b1111111111111110011101011;
    rom[59983] = 25'b1111111111111110011110000;
    rom[59984] = 25'b1111111111111110011110100;
    rom[59985] = 25'b1111111111111110011111000;
    rom[59986] = 25'b1111111111111110011111100;
    rom[59987] = 25'b1111111111111110100000000;
    rom[59988] = 25'b1111111111111110100000101;
    rom[59989] = 25'b1111111111111110100001000;
    rom[59990] = 25'b1111111111111110100001101;
    rom[59991] = 25'b1111111111111110100010001;
    rom[59992] = 25'b1111111111111110100010101;
    rom[59993] = 25'b1111111111111110100011001;
    rom[59994] = 25'b1111111111111110100011101;
    rom[59995] = 25'b1111111111111110100100001;
    rom[59996] = 25'b1111111111111110100100110;
    rom[59997] = 25'b1111111111111110100101010;
    rom[59998] = 25'b1111111111111110100101110;
    rom[59999] = 25'b1111111111111110100110010;
    rom[60000] = 25'b1111111111111110100110110;
    rom[60001] = 25'b1111111111111110100111011;
    rom[60002] = 25'b1111111111111110100111110;
    rom[60003] = 25'b1111111111111110101000011;
    rom[60004] = 25'b1111111111111110101000110;
    rom[60005] = 25'b1111111111111110101001011;
    rom[60006] = 25'b1111111111111110101001111;
    rom[60007] = 25'b1111111111111110101010011;
    rom[60008] = 25'b1111111111111110101010111;
    rom[60009] = 25'b1111111111111110101011011;
    rom[60010] = 25'b1111111111111110101011111;
    rom[60011] = 25'b1111111111111110101100100;
    rom[60012] = 25'b1111111111111110101100111;
    rom[60013] = 25'b1111111111111110101101100;
    rom[60014] = 25'b1111111111111110101110000;
    rom[60015] = 25'b1111111111111110101110100;
    rom[60016] = 25'b1111111111111110101111000;
    rom[60017] = 25'b1111111111111110101111100;
    rom[60018] = 25'b1111111111111110110000000;
    rom[60019] = 25'b1111111111111110110000100;
    rom[60020] = 25'b1111111111111110110001000;
    rom[60021] = 25'b1111111111111110110001100;
    rom[60022] = 25'b1111111111111110110010000;
    rom[60023] = 25'b1111111111111110110010100;
    rom[60024] = 25'b1111111111111110110011001;
    rom[60025] = 25'b1111111111111110110011100;
    rom[60026] = 25'b1111111111111110110100001;
    rom[60027] = 25'b1111111111111110110100101;
    rom[60028] = 25'b1111111111111110110101001;
    rom[60029] = 25'b1111111111111110110101101;
    rom[60030] = 25'b1111111111111110110110001;
    rom[60031] = 25'b1111111111111110110110101;
    rom[60032] = 25'b1111111111111110110111001;
    rom[60033] = 25'b1111111111111110110111101;
    rom[60034] = 25'b1111111111111110111000001;
    rom[60035] = 25'b1111111111111110111000101;
    rom[60036] = 25'b1111111111111110111001001;
    rom[60037] = 25'b1111111111111110111001101;
    rom[60038] = 25'b1111111111111110111010001;
    rom[60039] = 25'b1111111111111110111010101;
    rom[60040] = 25'b1111111111111110111011010;
    rom[60041] = 25'b1111111111111110111011101;
    rom[60042] = 25'b1111111111111110111100001;
    rom[60043] = 25'b1111111111111110111100110;
    rom[60044] = 25'b1111111111111110111101001;
    rom[60045] = 25'b1111111111111110111101110;
    rom[60046] = 25'b1111111111111110111110010;
    rom[60047] = 25'b1111111111111110111110101;
    rom[60048] = 25'b1111111111111110111111010;
    rom[60049] = 25'b1111111111111110111111101;
    rom[60050] = 25'b1111111111111111000000010;
    rom[60051] = 25'b1111111111111111000000110;
    rom[60052] = 25'b1111111111111111000001001;
    rom[60053] = 25'b1111111111111111000001110;
    rom[60054] = 25'b1111111111111111000010010;
    rom[60055] = 25'b1111111111111111000010101;
    rom[60056] = 25'b1111111111111111000011010;
    rom[60057] = 25'b1111111111111111000011110;
    rom[60058] = 25'b1111111111111111000100001;
    rom[60059] = 25'b1111111111111111000100110;
    rom[60060] = 25'b1111111111111111000101010;
    rom[60061] = 25'b1111111111111111000101101;
    rom[60062] = 25'b1111111111111111000110010;
    rom[60063] = 25'b1111111111111111000110110;
    rom[60064] = 25'b1111111111111111000111001;
    rom[60065] = 25'b1111111111111111000111110;
    rom[60066] = 25'b1111111111111111001000001;
    rom[60067] = 25'b1111111111111111001000101;
    rom[60068] = 25'b1111111111111111001001010;
    rom[60069] = 25'b1111111111111111001001101;
    rom[60070] = 25'b1111111111111111001010001;
    rom[60071] = 25'b1111111111111111001010110;
    rom[60072] = 25'b1111111111111111001011001;
    rom[60073] = 25'b1111111111111111001011101;
    rom[60074] = 25'b1111111111111111001100001;
    rom[60075] = 25'b1111111111111111001100101;
    rom[60076] = 25'b1111111111111111001101001;
    rom[60077] = 25'b1111111111111111001101101;
    rom[60078] = 25'b1111111111111111001110001;
    rom[60079] = 25'b1111111111111111001110101;
    rom[60080] = 25'b1111111111111111001111001;
    rom[60081] = 25'b1111111111111111001111101;
    rom[60082] = 25'b1111111111111111010000001;
    rom[60083] = 25'b1111111111111111010000101;
    rom[60084] = 25'b1111111111111111010001000;
    rom[60085] = 25'b1111111111111111010001100;
    rom[60086] = 25'b1111111111111111010010001;
    rom[60087] = 25'b1111111111111111010010100;
    rom[60088] = 25'b1111111111111111010011000;
    rom[60089] = 25'b1111111111111111010011100;
    rom[60090] = 25'b1111111111111111010100000;
    rom[60091] = 25'b1111111111111111010100100;
    rom[60092] = 25'b1111111111111111010101000;
    rom[60093] = 25'b1111111111111111010101100;
    rom[60094] = 25'b1111111111111111010110000;
    rom[60095] = 25'b1111111111111111010110100;
    rom[60096] = 25'b1111111111111111010111000;
    rom[60097] = 25'b1111111111111111010111011;
    rom[60098] = 25'b1111111111111111010111111;
    rom[60099] = 25'b1111111111111111011000011;
    rom[60100] = 25'b1111111111111111011000111;
    rom[60101] = 25'b1111111111111111011001011;
    rom[60102] = 25'b1111111111111111011001111;
    rom[60103] = 25'b1111111111111111011010010;
    rom[60104] = 25'b1111111111111111011010111;
    rom[60105] = 25'b1111111111111111011011011;
    rom[60106] = 25'b1111111111111111011011110;
    rom[60107] = 25'b1111111111111111011100010;
    rom[60108] = 25'b1111111111111111011100110;
    rom[60109] = 25'b1111111111111111011101010;
    rom[60110] = 25'b1111111111111111011101110;
    rom[60111] = 25'b1111111111111111011110010;
    rom[60112] = 25'b1111111111111111011110110;
    rom[60113] = 25'b1111111111111111011111001;
    rom[60114] = 25'b1111111111111111011111101;
    rom[60115] = 25'b1111111111111111100000001;
    rom[60116] = 25'b1111111111111111100000101;
    rom[60117] = 25'b1111111111111111100001001;
    rom[60118] = 25'b1111111111111111100001101;
    rom[60119] = 25'b1111111111111111100010000;
    rom[60120] = 25'b1111111111111111100010100;
    rom[60121] = 25'b1111111111111111100011000;
    rom[60122] = 25'b1111111111111111100011100;
    rom[60123] = 25'b1111111111111111100100000;
    rom[60124] = 25'b1111111111111111100100100;
    rom[60125] = 25'b1111111111111111100101000;
    rom[60126] = 25'b1111111111111111100101011;
    rom[60127] = 25'b1111111111111111100101111;
    rom[60128] = 25'b1111111111111111100110011;
    rom[60129] = 25'b1111111111111111100110111;
    rom[60130] = 25'b1111111111111111100111010;
    rom[60131] = 25'b1111111111111111100111110;
    rom[60132] = 25'b1111111111111111101000010;
    rom[60133] = 25'b1111111111111111101000110;
    rom[60134] = 25'b1111111111111111101001010;
    rom[60135] = 25'b1111111111111111101001110;
    rom[60136] = 25'b1111111111111111101010001;
    rom[60137] = 25'b1111111111111111101010101;
    rom[60138] = 25'b1111111111111111101011001;
    rom[60139] = 25'b1111111111111111101011101;
    rom[60140] = 25'b1111111111111111101100000;
    rom[60141] = 25'b1111111111111111101100100;
    rom[60142] = 25'b1111111111111111101101000;
    rom[60143] = 25'b1111111111111111101101100;
    rom[60144] = 25'b1111111111111111101101111;
    rom[60145] = 25'b1111111111111111101110011;
    rom[60146] = 25'b1111111111111111101110111;
    rom[60147] = 25'b1111111111111111101111011;
    rom[60148] = 25'b1111111111111111101111111;
    rom[60149] = 25'b1111111111111111110000011;
    rom[60150] = 25'b1111111111111111110000110;
    rom[60151] = 25'b1111111111111111110001010;
    rom[60152] = 25'b1111111111111111110001110;
    rom[60153] = 25'b1111111111111111110010010;
    rom[60154] = 25'b1111111111111111110010101;
    rom[60155] = 25'b1111111111111111110011001;
    rom[60156] = 25'b1111111111111111110011101;
    rom[60157] = 25'b1111111111111111110100001;
    rom[60158] = 25'b1111111111111111110100100;
    rom[60159] = 25'b1111111111111111110101000;
    rom[60160] = 25'b1111111111111111110101100;
    rom[60161] = 25'b1111111111111111110110000;
    rom[60162] = 25'b1111111111111111110110011;
    rom[60163] = 25'b1111111111111111110110111;
    rom[60164] = 25'b1111111111111111110111011;
    rom[60165] = 25'b1111111111111111110111110;
    rom[60166] = 25'b1111111111111111111000001;
    rom[60167] = 25'b1111111111111111111000101;
    rom[60168] = 25'b1111111111111111111001001;
    rom[60169] = 25'b1111111111111111111001101;
    rom[60170] = 25'b1111111111111111111010000;
    rom[60171] = 25'b1111111111111111111010100;
    rom[60172] = 25'b1111111111111111111011000;
    rom[60173] = 25'b1111111111111111111011100;
    rom[60174] = 25'b1111111111111111111011111;
    rom[60175] = 25'b1111111111111111111100011;
    rom[60176] = 25'b1111111111111111111100111;
    rom[60177] = 25'b1111111111111111111101011;
    rom[60178] = 25'b1111111111111111111101110;
    rom[60179] = 25'b1111111111111111111110010;
    rom[60180] = 25'b1111111111111111111110110;
    rom[60181] = 25'b1111111111111111111111001;
    rom[60182] = 25'b1111111111111111111111101;
    rom[60183] = 25'b0000000000000000000000000;
    rom[60184] = 25'b0000000000000000000000011;
    rom[60185] = 25'b0000000000000000000000111;
    rom[60186] = 25'b0000000000000000000001011;
    rom[60187] = 25'b0000000000000000000001110;
    rom[60188] = 25'b0000000000000000000010010;
    rom[60189] = 25'b0000000000000000000010110;
    rom[60190] = 25'b0000000000000000000011001;
    rom[60191] = 25'b0000000000000000000011101;
    rom[60192] = 25'b0000000000000000000100000;
    rom[60193] = 25'b0000000000000000000100100;
    rom[60194] = 25'b0000000000000000000101000;
    rom[60195] = 25'b0000000000000000000101100;
    rom[60196] = 25'b0000000000000000000101111;
    rom[60197] = 25'b0000000000000000000110010;
    rom[60198] = 25'b0000000000000000000110110;
    rom[60199] = 25'b0000000000000000000111010;
    rom[60200] = 25'b0000000000000000000111110;
    rom[60201] = 25'b0000000000000000001000001;
    rom[60202] = 25'b0000000000000000001000101;
    rom[60203] = 25'b0000000000000000001001000;
    rom[60204] = 25'b0000000000000000001001100;
    rom[60205] = 25'b0000000000000000001001111;
    rom[60206] = 25'b0000000000000000001010011;
    rom[60207] = 25'b0000000000000000001010111;
    rom[60208] = 25'b0000000000000000001011010;
    rom[60209] = 25'b0000000000000000001011110;
    rom[60210] = 25'b0000000000000000001100001;
    rom[60211] = 25'b0000000000000000001100101;
    rom[60212] = 25'b0000000000000000001101001;
    rom[60213] = 25'b0000000000000000001101100;
    rom[60214] = 25'b0000000000000000001110000;
    rom[60215] = 25'b0000000000000000001110011;
    rom[60216] = 25'b0000000000000000001110111;
    rom[60217] = 25'b0000000000000000001111010;
    rom[60218] = 25'b0000000000000000001111110;
    rom[60219] = 25'b0000000000000000010000001;
    rom[60220] = 25'b0000000000000000010000101;
    rom[60221] = 25'b0000000000000000010001000;
    rom[60222] = 25'b0000000000000000010001100;
    rom[60223] = 25'b0000000000000000010010000;
    rom[60224] = 25'b0000000000000000010010011;
    rom[60225] = 25'b0000000000000000010010110;
    rom[60226] = 25'b0000000000000000010011010;
    rom[60227] = 25'b0000000000000000010011110;
    rom[60228] = 25'b0000000000000000010100010;
    rom[60229] = 25'b0000000000000000010100101;
    rom[60230] = 25'b0000000000000000010101000;
    rom[60231] = 25'b0000000000000000010101100;
    rom[60232] = 25'b0000000000000000010101111;
    rom[60233] = 25'b0000000000000000010110011;
    rom[60234] = 25'b0000000000000000010110111;
    rom[60235] = 25'b0000000000000000010111010;
    rom[60236] = 25'b0000000000000000010111101;
    rom[60237] = 25'b0000000000000000011000001;
    rom[60238] = 25'b0000000000000000011000101;
    rom[60239] = 25'b0000000000000000011001000;
    rom[60240] = 25'b0000000000000000011001011;
    rom[60241] = 25'b0000000000000000011001111;
    rom[60242] = 25'b0000000000000000011010010;
    rom[60243] = 25'b0000000000000000011010110;
    rom[60244] = 25'b0000000000000000011011010;
    rom[60245] = 25'b0000000000000000011011101;
    rom[60246] = 25'b0000000000000000011100000;
    rom[60247] = 25'b0000000000000000011100100;
    rom[60248] = 25'b0000000000000000011100111;
    rom[60249] = 25'b0000000000000000011101011;
    rom[60250] = 25'b0000000000000000011101110;
    rom[60251] = 25'b0000000000000000011110010;
    rom[60252] = 25'b0000000000000000011110101;
    rom[60253] = 25'b0000000000000000011111000;
    rom[60254] = 25'b0000000000000000011111100;
    rom[60255] = 25'b0000000000000000100000000;
    rom[60256] = 25'b0000000000000000100000011;
    rom[60257] = 25'b0000000000000000100000110;
    rom[60258] = 25'b0000000000000000100001001;
    rom[60259] = 25'b0000000000000000100001101;
    rom[60260] = 25'b0000000000000000100010000;
    rom[60261] = 25'b0000000000000000100010100;
    rom[60262] = 25'b0000000000000000100011000;
    rom[60263] = 25'b0000000000000000100011011;
    rom[60264] = 25'b0000000000000000100011110;
    rom[60265] = 25'b0000000000000000100100001;
    rom[60266] = 25'b0000000000000000100100101;
    rom[60267] = 25'b0000000000000000100101000;
    rom[60268] = 25'b0000000000000000100101100;
    rom[60269] = 25'b0000000000000000100110000;
    rom[60270] = 25'b0000000000000000100110011;
    rom[60271] = 25'b0000000000000000100110110;
    rom[60272] = 25'b0000000000000000100111001;
    rom[60273] = 25'b0000000000000000100111101;
    rom[60274] = 25'b0000000000000000101000000;
    rom[60275] = 25'b0000000000000000101000100;
    rom[60276] = 25'b0000000000000000101000111;
    rom[60277] = 25'b0000000000000000101001010;
    rom[60278] = 25'b0000000000000000101001101;
    rom[60279] = 25'b0000000000000000101010001;
    rom[60280] = 25'b0000000000000000101010100;
    rom[60281] = 25'b0000000000000000101011000;
    rom[60282] = 25'b0000000000000000101011011;
    rom[60283] = 25'b0000000000000000101011111;
    rom[60284] = 25'b0000000000000000101100010;
    rom[60285] = 25'b0000000000000000101100101;
    rom[60286] = 25'b0000000000000000101101000;
    rom[60287] = 25'b0000000000000000101101100;
    rom[60288] = 25'b0000000000000000101101111;
    rom[60289] = 25'b0000000000000000101110011;
    rom[60290] = 25'b0000000000000000101110110;
    rom[60291] = 25'b0000000000000000101111010;
    rom[60292] = 25'b0000000000000000101111101;
    rom[60293] = 25'b0000000000000000110000000;
    rom[60294] = 25'b0000000000000000110000011;
    rom[60295] = 25'b0000000000000000110000110;
    rom[60296] = 25'b0000000000000000110001010;
    rom[60297] = 25'b0000000000000000110001101;
    rom[60298] = 25'b0000000000000000110010001;
    rom[60299] = 25'b0000000000000000110010100;
    rom[60300] = 25'b0000000000000000110010111;
    rom[60301] = 25'b0000000000000000110011010;
    rom[60302] = 25'b0000000000000000110011101;
    rom[60303] = 25'b0000000000000000110100001;
    rom[60304] = 25'b0000000000000000110100100;
    rom[60305] = 25'b0000000000000000110101000;
    rom[60306] = 25'b0000000000000000110101011;
    rom[60307] = 25'b0000000000000000110101110;
    rom[60308] = 25'b0000000000000000110110010;
    rom[60309] = 25'b0000000000000000110110101;
    rom[60310] = 25'b0000000000000000110111000;
    rom[60311] = 25'b0000000000000000110111011;
    rom[60312] = 25'b0000000000000000110111110;
    rom[60313] = 25'b0000000000000000111000010;
    rom[60314] = 25'b0000000000000000111000101;
    rom[60315] = 25'b0000000000000000111001000;
    rom[60316] = 25'b0000000000000000111001100;
    rom[60317] = 25'b0000000000000000111001111;
    rom[60318] = 25'b0000000000000000111010010;
    rom[60319] = 25'b0000000000000000111010101;
    rom[60320] = 25'b0000000000000000111011000;
    rom[60321] = 25'b0000000000000000111011011;
    rom[60322] = 25'b0000000000000000111011111;
    rom[60323] = 25'b0000000000000000111100010;
    rom[60324] = 25'b0000000000000000111100101;
    rom[60325] = 25'b0000000000000000111101001;
    rom[60326] = 25'b0000000000000000111101100;
    rom[60327] = 25'b0000000000000000111101111;
    rom[60328] = 25'b0000000000000000111110010;
    rom[60329] = 25'b0000000000000000111110110;
    rom[60330] = 25'b0000000000000000111111001;
    rom[60331] = 25'b0000000000000000111111100;
    rom[60332] = 25'b0000000000000000111111111;
    rom[60333] = 25'b0000000000000001000000010;
    rom[60334] = 25'b0000000000000001000000101;
    rom[60335] = 25'b0000000000000001000001000;
    rom[60336] = 25'b0000000000000001000001100;
    rom[60337] = 25'b0000000000000001000001111;
    rom[60338] = 25'b0000000000000001000010010;
    rom[60339] = 25'b0000000000000001000010101;
    rom[60340] = 25'b0000000000000001000011001;
    rom[60341] = 25'b0000000000000001000011100;
    rom[60342] = 25'b0000000000000001000011111;
    rom[60343] = 25'b0000000000000001000100010;
    rom[60344] = 25'b0000000000000001000100101;
    rom[60345] = 25'b0000000000000001000101000;
    rom[60346] = 25'b0000000000000001000101011;
    rom[60347] = 25'b0000000000000001000101110;
    rom[60348] = 25'b0000000000000001000110001;
    rom[60349] = 25'b0000000000000001000110101;
    rom[60350] = 25'b0000000000000001000111000;
    rom[60351] = 25'b0000000000000001000111011;
    rom[60352] = 25'b0000000000000001000111110;
    rom[60353] = 25'b0000000000000001001000001;
    rom[60354] = 25'b0000000000000001001000101;
    rom[60355] = 25'b0000000000000001001001000;
    rom[60356] = 25'b0000000000000001001001011;
    rom[60357] = 25'b0000000000000001001001110;
    rom[60358] = 25'b0000000000000001001010001;
    rom[60359] = 25'b0000000000000001001010100;
    rom[60360] = 25'b0000000000000001001010111;
    rom[60361] = 25'b0000000000000001001011010;
    rom[60362] = 25'b0000000000000001001011101;
    rom[60363] = 25'b0000000000000001001100000;
    rom[60364] = 25'b0000000000000001001100011;
    rom[60365] = 25'b0000000000000001001100110;
    rom[60366] = 25'b0000000000000001001101001;
    rom[60367] = 25'b0000000000000001001101101;
    rom[60368] = 25'b0000000000000001001110000;
    rom[60369] = 25'b0000000000000001001110011;
    rom[60370] = 25'b0000000000000001001110110;
    rom[60371] = 25'b0000000000000001001111001;
    rom[60372] = 25'b0000000000000001001111100;
    rom[60373] = 25'b0000000000000001001111111;
    rom[60374] = 25'b0000000000000001010000010;
    rom[60375] = 25'b0000000000000001010000101;
    rom[60376] = 25'b0000000000000001010001000;
    rom[60377] = 25'b0000000000000001010001011;
    rom[60378] = 25'b0000000000000001010001111;
    rom[60379] = 25'b0000000000000001010010010;
    rom[60380] = 25'b0000000000000001010010101;
    rom[60381] = 25'b0000000000000001010011000;
    rom[60382] = 25'b0000000000000001010011011;
    rom[60383] = 25'b0000000000000001010011110;
    rom[60384] = 25'b0000000000000001010100001;
    rom[60385] = 25'b0000000000000001010100100;
    rom[60386] = 25'b0000000000000001010100111;
    rom[60387] = 25'b0000000000000001010101010;
    rom[60388] = 25'b0000000000000001010101101;
    rom[60389] = 25'b0000000000000001010110000;
    rom[60390] = 25'b0000000000000001010110011;
    rom[60391] = 25'b0000000000000001010110110;
    rom[60392] = 25'b0000000000000001010111001;
    rom[60393] = 25'b0000000000000001010111100;
    rom[60394] = 25'b0000000000000001010111111;
    rom[60395] = 25'b0000000000000001011000010;
    rom[60396] = 25'b0000000000000001011000100;
    rom[60397] = 25'b0000000000000001011000111;
    rom[60398] = 25'b0000000000000001011001010;
    rom[60399] = 25'b0000000000000001011001101;
    rom[60400] = 25'b0000000000000001011010000;
    rom[60401] = 25'b0000000000000001011010011;
    rom[60402] = 25'b0000000000000001011010110;
    rom[60403] = 25'b0000000000000001011011001;
    rom[60404] = 25'b0000000000000001011011100;
    rom[60405] = 25'b0000000000000001011011111;
    rom[60406] = 25'b0000000000000001011100010;
    rom[60407] = 25'b0000000000000001011100101;
    rom[60408] = 25'b0000000000000001011101000;
    rom[60409] = 25'b0000000000000001011101011;
    rom[60410] = 25'b0000000000000001011101110;
    rom[60411] = 25'b0000000000000001011110001;
    rom[60412] = 25'b0000000000000001011110100;
    rom[60413] = 25'b0000000000000001011110111;
    rom[60414] = 25'b0000000000000001011111010;
    rom[60415] = 25'b0000000000000001011111101;
    rom[60416] = 25'b0000000000000001100000000;
    rom[60417] = 25'b0000000000000001100000011;
    rom[60418] = 25'b0000000000000001100000101;
    rom[60419] = 25'b0000000000000001100001000;
    rom[60420] = 25'b0000000000000001100001011;
    rom[60421] = 25'b0000000000000001100001110;
    rom[60422] = 25'b0000000000000001100010001;
    rom[60423] = 25'b0000000000000001100010100;
    rom[60424] = 25'b0000000000000001100010111;
    rom[60425] = 25'b0000000000000001100011010;
    rom[60426] = 25'b0000000000000001100011101;
    rom[60427] = 25'b0000000000000001100011111;
    rom[60428] = 25'b0000000000000001100100010;
    rom[60429] = 25'b0000000000000001100100101;
    rom[60430] = 25'b0000000000000001100101000;
    rom[60431] = 25'b0000000000000001100101011;
    rom[60432] = 25'b0000000000000001100101110;
    rom[60433] = 25'b0000000000000001100110000;
    rom[60434] = 25'b0000000000000001100110011;
    rom[60435] = 25'b0000000000000001100110110;
    rom[60436] = 25'b0000000000000001100111001;
    rom[60437] = 25'b0000000000000001100111100;
    rom[60438] = 25'b0000000000000001100111110;
    rom[60439] = 25'b0000000000000001101000001;
    rom[60440] = 25'b0000000000000001101000100;
    rom[60441] = 25'b0000000000000001101000111;
    rom[60442] = 25'b0000000000000001101001010;
    rom[60443] = 25'b0000000000000001101001100;
    rom[60444] = 25'b0000000000000001101001111;
    rom[60445] = 25'b0000000000000001101010010;
    rom[60446] = 25'b0000000000000001101010101;
    rom[60447] = 25'b0000000000000001101011000;
    rom[60448] = 25'b0000000000000001101011011;
    rom[60449] = 25'b0000000000000001101011110;
    rom[60450] = 25'b0000000000000001101100001;
    rom[60451] = 25'b0000000000000001101100011;
    rom[60452] = 25'b0000000000000001101100110;
    rom[60453] = 25'b0000000000000001101101001;
    rom[60454] = 25'b0000000000000001101101011;
    rom[60455] = 25'b0000000000000001101101110;
    rom[60456] = 25'b0000000000000001101110001;
    rom[60457] = 25'b0000000000000001101110100;
    rom[60458] = 25'b0000000000000001101110110;
    rom[60459] = 25'b0000000000000001101111001;
    rom[60460] = 25'b0000000000000001101111100;
    rom[60461] = 25'b0000000000000001101111111;
    rom[60462] = 25'b0000000000000001110000010;
    rom[60463] = 25'b0000000000000001110000100;
    rom[60464] = 25'b0000000000000001110000111;
    rom[60465] = 25'b0000000000000001110001010;
    rom[60466] = 25'b0000000000000001110001101;
    rom[60467] = 25'b0000000000000001110001111;
    rom[60468] = 25'b0000000000000001110010010;
    rom[60469] = 25'b0000000000000001110010101;
    rom[60470] = 25'b0000000000000001110010111;
    rom[60471] = 25'b0000000000000001110011010;
    rom[60472] = 25'b0000000000000001110011101;
    rom[60473] = 25'b0000000000000001110011111;
    rom[60474] = 25'b0000000000000001110100010;
    rom[60475] = 25'b0000000000000001110100101;
    rom[60476] = 25'b0000000000000001110101000;
    rom[60477] = 25'b0000000000000001110101011;
    rom[60478] = 25'b0000000000000001110101101;
    rom[60479] = 25'b0000000000000001110110000;
    rom[60480] = 25'b0000000000000001110110010;
    rom[60481] = 25'b0000000000000001110110101;
    rom[60482] = 25'b0000000000000001110111000;
    rom[60483] = 25'b0000000000000001110111010;
    rom[60484] = 25'b0000000000000001110111101;
    rom[60485] = 25'b0000000000000001111000000;
    rom[60486] = 25'b0000000000000001111000011;
    rom[60487] = 25'b0000000000000001111000101;
    rom[60488] = 25'b0000000000000001111001000;
    rom[60489] = 25'b0000000000000001111001011;
    rom[60490] = 25'b0000000000000001111001101;
    rom[60491] = 25'b0000000000000001111010000;
    rom[60492] = 25'b0000000000000001111010010;
    rom[60493] = 25'b0000000000000001111010101;
    rom[60494] = 25'b0000000000000001111010111;
    rom[60495] = 25'b0000000000000001111011010;
    rom[60496] = 25'b0000000000000001111011101;
    rom[60497] = 25'b0000000000000001111100000;
    rom[60498] = 25'b0000000000000001111100010;
    rom[60499] = 25'b0000000000000001111100101;
    rom[60500] = 25'b0000000000000001111100111;
    rom[60501] = 25'b0000000000000001111101010;
    rom[60502] = 25'b0000000000000001111101100;
    rom[60503] = 25'b0000000000000001111101111;
    rom[60504] = 25'b0000000000000001111110010;
    rom[60505] = 25'b0000000000000001111110101;
    rom[60506] = 25'b0000000000000001111110111;
    rom[60507] = 25'b0000000000000001111111010;
    rom[60508] = 25'b0000000000000001111111100;
    rom[60509] = 25'b0000000000000001111111111;
    rom[60510] = 25'b0000000000000010000000001;
    rom[60511] = 25'b0000000000000010000000100;
    rom[60512] = 25'b0000000000000010000000110;
    rom[60513] = 25'b0000000000000010000001001;
    rom[60514] = 25'b0000000000000010000001100;
    rom[60515] = 25'b0000000000000010000001110;
    rom[60516] = 25'b0000000000000010000010001;
    rom[60517] = 25'b0000000000000010000010011;
    rom[60518] = 25'b0000000000000010000010110;
    rom[60519] = 25'b0000000000000010000011000;
    rom[60520] = 25'b0000000000000010000011011;
    rom[60521] = 25'b0000000000000010000011110;
    rom[60522] = 25'b0000000000000010000100000;
    rom[60523] = 25'b0000000000000010000100011;
    rom[60524] = 25'b0000000000000010000100101;
    rom[60525] = 25'b0000000000000010000100111;
    rom[60526] = 25'b0000000000000010000101010;
    rom[60527] = 25'b0000000000000010000101101;
    rom[60528] = 25'b0000000000000010000101111;
    rom[60529] = 25'b0000000000000010000110010;
    rom[60530] = 25'b0000000000000010000110100;
    rom[60531] = 25'b0000000000000010000110110;
    rom[60532] = 25'b0000000000000010000111001;
    rom[60533] = 25'b0000000000000010000111100;
    rom[60534] = 25'b0000000000000010000111110;
    rom[60535] = 25'b0000000000000010001000001;
    rom[60536] = 25'b0000000000000010001000011;
    rom[60537] = 25'b0000000000000010001000101;
    rom[60538] = 25'b0000000000000010001001000;
    rom[60539] = 25'b0000000000000010001001010;
    rom[60540] = 25'b0000000000000010001001101;
    rom[60541] = 25'b0000000000000010001010000;
    rom[60542] = 25'b0000000000000010001010010;
    rom[60543] = 25'b0000000000000010001010100;
    rom[60544] = 25'b0000000000000010001010111;
    rom[60545] = 25'b0000000000000010001011001;
    rom[60546] = 25'b0000000000000010001011100;
    rom[60547] = 25'b0000000000000010001011110;
    rom[60548] = 25'b0000000000000010001100001;
    rom[60549] = 25'b0000000000000010001100011;
    rom[60550] = 25'b0000000000000010001100101;
    rom[60551] = 25'b0000000000000010001101000;
    rom[60552] = 25'b0000000000000010001101011;
    rom[60553] = 25'b0000000000000010001101101;
    rom[60554] = 25'b0000000000000010001101111;
    rom[60555] = 25'b0000000000000010001110001;
    rom[60556] = 25'b0000000000000010001110100;
    rom[60557] = 25'b0000000000000010001110111;
    rom[60558] = 25'b0000000000000010001111001;
    rom[60559] = 25'b0000000000000010001111011;
    rom[60560] = 25'b0000000000000010001111101;
    rom[60561] = 25'b0000000000000010010000000;
    rom[60562] = 25'b0000000000000010010000011;
    rom[60563] = 25'b0000000000000010010000101;
    rom[60564] = 25'b0000000000000010010000111;
    rom[60565] = 25'b0000000000000010010001001;
    rom[60566] = 25'b0000000000000010010001100;
    rom[60567] = 25'b0000000000000010010001110;
    rom[60568] = 25'b0000000000000010010010001;
    rom[60569] = 25'b0000000000000010010010011;
    rom[60570] = 25'b0000000000000010010010101;
    rom[60571] = 25'b0000000000000010010010111;
    rom[60572] = 25'b0000000000000010010011010;
    rom[60573] = 25'b0000000000000010010011101;
    rom[60574] = 25'b0000000000000010010011111;
    rom[60575] = 25'b0000000000000010010100001;
    rom[60576] = 25'b0000000000000010010100011;
    rom[60577] = 25'b0000000000000010010100110;
    rom[60578] = 25'b0000000000000010010101000;
    rom[60579] = 25'b0000000000000010010101010;
    rom[60580] = 25'b0000000000000010010101101;
    rom[60581] = 25'b0000000000000010010101111;
    rom[60582] = 25'b0000000000000010010110010;
    rom[60583] = 25'b0000000000000010010110100;
    rom[60584] = 25'b0000000000000010010110110;
    rom[60585] = 25'b0000000000000010010111000;
    rom[60586] = 25'b0000000000000010010111011;
    rom[60587] = 25'b0000000000000010010111101;
    rom[60588] = 25'b0000000000000010010111111;
    rom[60589] = 25'b0000000000000010011000001;
    rom[60590] = 25'b0000000000000010011000100;
    rom[60591] = 25'b0000000000000010011000110;
    rom[60592] = 25'b0000000000000010011001001;
    rom[60593] = 25'b0000000000000010011001011;
    rom[60594] = 25'b0000000000000010011001101;
    rom[60595] = 25'b0000000000000010011001111;
    rom[60596] = 25'b0000000000000010011010010;
    rom[60597] = 25'b0000000000000010011010100;
    rom[60598] = 25'b0000000000000010011010110;
    rom[60599] = 25'b0000000000000010011011000;
    rom[60600] = 25'b0000000000000010011011011;
    rom[60601] = 25'b0000000000000010011011101;
    rom[60602] = 25'b0000000000000010011011111;
    rom[60603] = 25'b0000000000000010011100001;
    rom[60604] = 25'b0000000000000010011100100;
    rom[60605] = 25'b0000000000000010011100110;
    rom[60606] = 25'b0000000000000010011101000;
    rom[60607] = 25'b0000000000000010011101010;
    rom[60608] = 25'b0000000000000010011101101;
    rom[60609] = 25'b0000000000000010011101111;
    rom[60610] = 25'b0000000000000010011110001;
    rom[60611] = 25'b0000000000000010011110011;
    rom[60612] = 25'b0000000000000010011110110;
    rom[60613] = 25'b0000000000000010011111000;
    rom[60614] = 25'b0000000000000010011111001;
    rom[60615] = 25'b0000000000000010011111100;
    rom[60616] = 25'b0000000000000010011111110;
    rom[60617] = 25'b0000000000000010100000000;
    rom[60618] = 25'b0000000000000010100000010;
    rom[60619] = 25'b0000000000000010100000101;
    rom[60620] = 25'b0000000000000010100000111;
    rom[60621] = 25'b0000000000000010100001001;
    rom[60622] = 25'b0000000000000010100001011;
    rom[60623] = 25'b0000000000000010100001101;
    rom[60624] = 25'b0000000000000010100010000;
    rom[60625] = 25'b0000000000000010100010010;
    rom[60626] = 25'b0000000000000010100010011;
    rom[60627] = 25'b0000000000000010100010110;
    rom[60628] = 25'b0000000000000010100011000;
    rom[60629] = 25'b0000000000000010100011010;
    rom[60630] = 25'b0000000000000010100011100;
    rom[60631] = 25'b0000000000000010100011111;
    rom[60632] = 25'b0000000000000010100100001;
    rom[60633] = 25'b0000000000000010100100010;
    rom[60634] = 25'b0000000000000010100100101;
    rom[60635] = 25'b0000000000000010100100111;
    rom[60636] = 25'b0000000000000010100101001;
    rom[60637] = 25'b0000000000000010100101011;
    rom[60638] = 25'b0000000000000010100101110;
    rom[60639] = 25'b0000000000000010100101111;
    rom[60640] = 25'b0000000000000010100110001;
    rom[60641] = 25'b0000000000000010100110100;
    rom[60642] = 25'b0000000000000010100110110;
    rom[60643] = 25'b0000000000000010100111000;
    rom[60644] = 25'b0000000000000010100111010;
    rom[60645] = 25'b0000000000000010100111100;
    rom[60646] = 25'b0000000000000010100111110;
    rom[60647] = 25'b0000000000000010101000000;
    rom[60648] = 25'b0000000000000010101000011;
    rom[60649] = 25'b0000000000000010101000100;
    rom[60650] = 25'b0000000000000010101000110;
    rom[60651] = 25'b0000000000000010101001000;
    rom[60652] = 25'b0000000000000010101001011;
    rom[60653] = 25'b0000000000000010101001100;
    rom[60654] = 25'b0000000000000010101001110;
    rom[60655] = 25'b0000000000000010101010001;
    rom[60656] = 25'b0000000000000010101010011;
    rom[60657] = 25'b0000000000000010101010100;
    rom[60658] = 25'b0000000000000010101010111;
    rom[60659] = 25'b0000000000000010101011001;
    rom[60660] = 25'b0000000000000010101011011;
    rom[60661] = 25'b0000000000000010101011101;
    rom[60662] = 25'b0000000000000010101011111;
    rom[60663] = 25'b0000000000000010101100001;
    rom[60664] = 25'b0000000000000010101100011;
    rom[60665] = 25'b0000000000000010101100101;
    rom[60666] = 25'b0000000000000010101100111;
    rom[60667] = 25'b0000000000000010101101001;
    rom[60668] = 25'b0000000000000010101101011;
    rom[60669] = 25'b0000000000000010101101101;
    rom[60670] = 25'b0000000000000010101101111;
    rom[60671] = 25'b0000000000000010101110001;
    rom[60672] = 25'b0000000000000010101110011;
    rom[60673] = 25'b0000000000000010101110101;
    rom[60674] = 25'b0000000000000010101110111;
    rom[60675] = 25'b0000000000000010101111001;
    rom[60676] = 25'b0000000000000010101111011;
    rom[60677] = 25'b0000000000000010101111101;
    rom[60678] = 25'b0000000000000010101111111;
    rom[60679] = 25'b0000000000000010110000001;
    rom[60680] = 25'b0000000000000010110000011;
    rom[60681] = 25'b0000000000000010110000100;
    rom[60682] = 25'b0000000000000010110000111;
    rom[60683] = 25'b0000000000000010110001001;
    rom[60684] = 25'b0000000000000010110001010;
    rom[60685] = 25'b0000000000000010110001100;
    rom[60686] = 25'b0000000000000010110001110;
    rom[60687] = 25'b0000000000000010110010000;
    rom[60688] = 25'b0000000000000010110010010;
    rom[60689] = 25'b0000000000000010110010100;
    rom[60690] = 25'b0000000000000010110010110;
    rom[60691] = 25'b0000000000000010110011000;
    rom[60692] = 25'b0000000000000010110011010;
    rom[60693] = 25'b0000000000000010110011011;
    rom[60694] = 25'b0000000000000010110011110;
    rom[60695] = 25'b0000000000000010110011111;
    rom[60696] = 25'b0000000000000010110100001;
    rom[60697] = 25'b0000000000000010110100100;
    rom[60698] = 25'b0000000000000010110100101;
    rom[60699] = 25'b0000000000000010110100111;
    rom[60700] = 25'b0000000000000010110101001;
    rom[60701] = 25'b0000000000000010110101011;
    rom[60702] = 25'b0000000000000010110101101;
    rom[60703] = 25'b0000000000000010110101111;
    rom[60704] = 25'b0000000000000010110110000;
    rom[60705] = 25'b0000000000000010110110011;
    rom[60706] = 25'b0000000000000010110110100;
    rom[60707] = 25'b0000000000000010110110110;
    rom[60708] = 25'b0000000000000010110111000;
    rom[60709] = 25'b0000000000000010110111010;
    rom[60710] = 25'b0000000000000010110111100;
    rom[60711] = 25'b0000000000000010110111110;
    rom[60712] = 25'b0000000000000010110111111;
    rom[60713] = 25'b0000000000000010111000001;
    rom[60714] = 25'b0000000000000010111000011;
    rom[60715] = 25'b0000000000000010111000101;
    rom[60716] = 25'b0000000000000010111000111;
    rom[60717] = 25'b0000000000000010111001000;
    rom[60718] = 25'b0000000000000010111001010;
    rom[60719] = 25'b0000000000000010111001100;
    rom[60720] = 25'b0000000000000010111001101;
    rom[60721] = 25'b0000000000000010111010000;
    rom[60722] = 25'b0000000000000010111010001;
    rom[60723] = 25'b0000000000000010111010011;
    rom[60724] = 25'b0000000000000010111010101;
    rom[60725] = 25'b0000000000000010111010111;
    rom[60726] = 25'b0000000000000010111011001;
    rom[60727] = 25'b0000000000000010111011010;
    rom[60728] = 25'b0000000000000010111011100;
    rom[60729] = 25'b0000000000000010111011110;
    rom[60730] = 25'b0000000000000010111011111;
    rom[60731] = 25'b0000000000000010111100010;
    rom[60732] = 25'b0000000000000010111100011;
    rom[60733] = 25'b0000000000000010111100101;
    rom[60734] = 25'b0000000000000010111100111;
    rom[60735] = 25'b0000000000000010111101000;
    rom[60736] = 25'b0000000000000010111101011;
    rom[60737] = 25'b0000000000000010111101100;
    rom[60738] = 25'b0000000000000010111101110;
    rom[60739] = 25'b0000000000000010111110000;
    rom[60740] = 25'b0000000000000010111110001;
    rom[60741] = 25'b0000000000000010111110011;
    rom[60742] = 25'b0000000000000010111110100;
    rom[60743] = 25'b0000000000000010111110111;
    rom[60744] = 25'b0000000000000010111111000;
    rom[60745] = 25'b0000000000000010111111010;
    rom[60746] = 25'b0000000000000010111111100;
    rom[60747] = 25'b0000000000000010111111101;
    rom[60748] = 25'b0000000000000010111111111;
    rom[60749] = 25'b0000000000000011000000001;
    rom[60750] = 25'b0000000000000011000000011;
    rom[60751] = 25'b0000000000000011000000100;
    rom[60752] = 25'b0000000000000011000000110;
    rom[60753] = 25'b0000000000000011000001000;
    rom[60754] = 25'b0000000000000011000001001;
    rom[60755] = 25'b0000000000000011000001011;
    rom[60756] = 25'b0000000000000011000001100;
    rom[60757] = 25'b0000000000000011000001110;
    rom[60758] = 25'b0000000000000011000010000;
    rom[60759] = 25'b0000000000000011000010001;
    rom[60760] = 25'b0000000000000011000010011;
    rom[60761] = 25'b0000000000000011000010100;
    rom[60762] = 25'b0000000000000011000010111;
    rom[60763] = 25'b0000000000000011000011000;
    rom[60764] = 25'b0000000000000011000011010;
    rom[60765] = 25'b0000000000000011000011011;
    rom[60766] = 25'b0000000000000011000011101;
    rom[60767] = 25'b0000000000000011000011111;
    rom[60768] = 25'b0000000000000011000100000;
    rom[60769] = 25'b0000000000000011000100010;
    rom[60770] = 25'b0000000000000011000100011;
    rom[60771] = 25'b0000000000000011000100101;
    rom[60772] = 25'b0000000000000011000100111;
    rom[60773] = 25'b0000000000000011000101001;
    rom[60774] = 25'b0000000000000011000101010;
    rom[60775] = 25'b0000000000000011000101100;
    rom[60776] = 25'b0000000000000011000101101;
    rom[60777] = 25'b0000000000000011000101111;
    rom[60778] = 25'b0000000000000011000110000;
    rom[60779] = 25'b0000000000000011000110010;
    rom[60780] = 25'b0000000000000011000110100;
    rom[60781] = 25'b0000000000000011000110101;
    rom[60782] = 25'b0000000000000011000110111;
    rom[60783] = 25'b0000000000000011000111000;
    rom[60784] = 25'b0000000000000011000111010;
    rom[60785] = 25'b0000000000000011000111011;
    rom[60786] = 25'b0000000000000011000111101;
    rom[60787] = 25'b0000000000000011000111110;
    rom[60788] = 25'b0000000000000011001000000;
    rom[60789] = 25'b0000000000000011001000010;
    rom[60790] = 25'b0000000000000011001000100;
    rom[60791] = 25'b0000000000000011001000101;
    rom[60792] = 25'b0000000000000011001000111;
    rom[60793] = 25'b0000000000000011001001000;
    rom[60794] = 25'b0000000000000011001001001;
    rom[60795] = 25'b0000000000000011001001011;
    rom[60796] = 25'b0000000000000011001001100;
    rom[60797] = 25'b0000000000000011001001110;
    rom[60798] = 25'b0000000000000011001001111;
    rom[60799] = 25'b0000000000000011001010001;
    rom[60800] = 25'b0000000000000011001010010;
    rom[60801] = 25'b0000000000000011001010100;
    rom[60802] = 25'b0000000000000011001010101;
    rom[60803] = 25'b0000000000000011001010111;
    rom[60804] = 25'b0000000000000011001011000;
    rom[60805] = 25'b0000000000000011001011010;
    rom[60806] = 25'b0000000000000011001011011;
    rom[60807] = 25'b0000000000000011001011101;
    rom[60808] = 25'b0000000000000011001011110;
    rom[60809] = 25'b0000000000000011001100000;
    rom[60810] = 25'b0000000000000011001100001;
    rom[60811] = 25'b0000000000000011001100011;
    rom[60812] = 25'b0000000000000011001100100;
    rom[60813] = 25'b0000000000000011001100110;
    rom[60814] = 25'b0000000000000011001100111;
    rom[60815] = 25'b0000000000000011001101001;
    rom[60816] = 25'b0000000000000011001101010;
    rom[60817] = 25'b0000000000000011001101100;
    rom[60818] = 25'b0000000000000011001101101;
    rom[60819] = 25'b0000000000000011001101111;
    rom[60820] = 25'b0000000000000011001110000;
    rom[60821] = 25'b0000000000000011001110010;
    rom[60822] = 25'b0000000000000011001110011;
    rom[60823] = 25'b0000000000000011001110100;
    rom[60824] = 25'b0000000000000011001110110;
    rom[60825] = 25'b0000000000000011001110111;
    rom[60826] = 25'b0000000000000011001111001;
    rom[60827] = 25'b0000000000000011001111010;
    rom[60828] = 25'b0000000000000011001111100;
    rom[60829] = 25'b0000000000000011001111101;
    rom[60830] = 25'b0000000000000011001111111;
    rom[60831] = 25'b0000000000000011010000000;
    rom[60832] = 25'b0000000000000011010000001;
    rom[60833] = 25'b0000000000000011010000010;
    rom[60834] = 25'b0000000000000011010000100;
    rom[60835] = 25'b0000000000000011010000101;
    rom[60836] = 25'b0000000000000011010000111;
    rom[60837] = 25'b0000000000000011010001000;
    rom[60838] = 25'b0000000000000011010001010;
    rom[60839] = 25'b0000000000000011010001010;
    rom[60840] = 25'b0000000000000011010001100;
    rom[60841] = 25'b0000000000000011010001101;
    rom[60842] = 25'b0000000000000011010001111;
    rom[60843] = 25'b0000000000000011010010000;
    rom[60844] = 25'b0000000000000011010010001;
    rom[60845] = 25'b0000000000000011010010011;
    rom[60846] = 25'b0000000000000011010010100;
    rom[60847] = 25'b0000000000000011010010110;
    rom[60848] = 25'b0000000000000011010010111;
    rom[60849] = 25'b0000000000000011010011000;
    rom[60850] = 25'b0000000000000011010011001;
    rom[60851] = 25'b0000000000000011010011011;
    rom[60852] = 25'b0000000000000011010011100;
    rom[60853] = 25'b0000000000000011010011110;
    rom[60854] = 25'b0000000000000011010011111;
    rom[60855] = 25'b0000000000000011010100000;
    rom[60856] = 25'b0000000000000011010100010;
    rom[60857] = 25'b0000000000000011010100011;
    rom[60858] = 25'b0000000000000011010100100;
    rom[60859] = 25'b0000000000000011010100101;
    rom[60860] = 25'b0000000000000011010100111;
    rom[60861] = 25'b0000000000000011010101000;
    rom[60862] = 25'b0000000000000011010101001;
    rom[60863] = 25'b0000000000000011010101011;
    rom[60864] = 25'b0000000000000011010101100;
    rom[60865] = 25'b0000000000000011010101101;
    rom[60866] = 25'b0000000000000011010101110;
    rom[60867] = 25'b0000000000000011010110000;
    rom[60868] = 25'b0000000000000011010110001;
    rom[60869] = 25'b0000000000000011010110010;
    rom[60870] = 25'b0000000000000011010110100;
    rom[60871] = 25'b0000000000000011010110101;
    rom[60872] = 25'b0000000000000011010110110;
    rom[60873] = 25'b0000000000000011010110111;
    rom[60874] = 25'b0000000000000011010111001;
    rom[60875] = 25'b0000000000000011010111010;
    rom[60876] = 25'b0000000000000011010111011;
    rom[60877] = 25'b0000000000000011010111101;
    rom[60878] = 25'b0000000000000011010111101;
    rom[60879] = 25'b0000000000000011010111111;
    rom[60880] = 25'b0000000000000011011000000;
    rom[60881] = 25'b0000000000000011011000001;
    rom[60882] = 25'b0000000000000011011000011;
    rom[60883] = 25'b0000000000000011011000011;
    rom[60884] = 25'b0000000000000011011000101;
    rom[60885] = 25'b0000000000000011011000110;
    rom[60886] = 25'b0000000000000011011000111;
    rom[60887] = 25'b0000000000000011011001000;
    rom[60888] = 25'b0000000000000011011001001;
    rom[60889] = 25'b0000000000000011011001011;
    rom[60890] = 25'b0000000000000011011001100;
    rom[60891] = 25'b0000000000000011011001101;
    rom[60892] = 25'b0000000000000011011001110;
    rom[60893] = 25'b0000000000000011011001111;
    rom[60894] = 25'b0000000000000011011010001;
    rom[60895] = 25'b0000000000000011011010001;
    rom[60896] = 25'b0000000000000011011010011;
    rom[60897] = 25'b0000000000000011011010100;
    rom[60898] = 25'b0000000000000011011010101;
    rom[60899] = 25'b0000000000000011011010111;
    rom[60900] = 25'b0000000000000011011010111;
    rom[60901] = 25'b0000000000000011011011001;
    rom[60902] = 25'b0000000000000011011011010;
    rom[60903] = 25'b0000000000000011011011011;
    rom[60904] = 25'b0000000000000011011011100;
    rom[60905] = 25'b0000000000000011011011101;
    rom[60906] = 25'b0000000000000011011011110;
    rom[60907] = 25'b0000000000000011011100000;
    rom[60908] = 25'b0000000000000011011100000;
    rom[60909] = 25'b0000000000000011011100010;
    rom[60910] = 25'b0000000000000011011100011;
    rom[60911] = 25'b0000000000000011011100100;
    rom[60912] = 25'b0000000000000011011100101;
    rom[60913] = 25'b0000000000000011011100110;
    rom[60914] = 25'b0000000000000011011100111;
    rom[60915] = 25'b0000000000000011011101001;
    rom[60916] = 25'b0000000000000011011101001;
    rom[60917] = 25'b0000000000000011011101011;
    rom[60918] = 25'b0000000000000011011101100;
    rom[60919] = 25'b0000000000000011011101101;
    rom[60920] = 25'b0000000000000011011101110;
    rom[60921] = 25'b0000000000000011011101111;
    rom[60922] = 25'b0000000000000011011110000;
    rom[60923] = 25'b0000000000000011011110001;
    rom[60924] = 25'b0000000000000011011110010;
    rom[60925] = 25'b0000000000000011011110011;
    rom[60926] = 25'b0000000000000011011110101;
    rom[60927] = 25'b0000000000000011011110101;
    rom[60928] = 25'b0000000000000011011110110;
    rom[60929] = 25'b0000000000000011011111000;
    rom[60930] = 25'b0000000000000011011111000;
    rom[60931] = 25'b0000000000000011011111010;
    rom[60932] = 25'b0000000000000011011111011;
    rom[60933] = 25'b0000000000000011011111011;
    rom[60934] = 25'b0000000000000011011111101;
    rom[60935] = 25'b0000000000000011011111110;
    rom[60936] = 25'b0000000000000011011111111;
    rom[60937] = 25'b0000000000000011100000000;
    rom[60938] = 25'b0000000000000011100000001;
    rom[60939] = 25'b0000000000000011100000010;
    rom[60940] = 25'b0000000000000011100000011;
    rom[60941] = 25'b0000000000000011100000100;
    rom[60942] = 25'b0000000000000011100000101;
    rom[60943] = 25'b0000000000000011100000110;
    rom[60944] = 25'b0000000000000011100000111;
    rom[60945] = 25'b0000000000000011100001000;
    rom[60946] = 25'b0000000000000011100001001;
    rom[60947] = 25'b0000000000000011100001001;
    rom[60948] = 25'b0000000000000011100001011;
    rom[60949] = 25'b0000000000000011100001100;
    rom[60950] = 25'b0000000000000011100001100;
    rom[60951] = 25'b0000000000000011100001110;
    rom[60952] = 25'b0000000000000011100001111;
    rom[60953] = 25'b0000000000000011100001111;
    rom[60954] = 25'b0000000000000011100010000;
    rom[60955] = 25'b0000000000000011100010010;
    rom[60956] = 25'b0000000000000011100010010;
    rom[60957] = 25'b0000000000000011100010011;
    rom[60958] = 25'b0000000000000011100010101;
    rom[60959] = 25'b0000000000000011100010101;
    rom[60960] = 25'b0000000000000011100010110;
    rom[60961] = 25'b0000000000000011100010111;
    rom[60962] = 25'b0000000000000011100011000;
    rom[60963] = 25'b0000000000000011100011001;
    rom[60964] = 25'b0000000000000011100011010;
    rom[60965] = 25'b0000000000000011100011011;
    rom[60966] = 25'b0000000000000011100011100;
    rom[60967] = 25'b0000000000000011100011101;
    rom[60968] = 25'b0000000000000011100011110;
    rom[60969] = 25'b0000000000000011100011110;
    rom[60970] = 25'b0000000000000011100011111;
    rom[60971] = 25'b0000000000000011100100001;
    rom[60972] = 25'b0000000000000011100100001;
    rom[60973] = 25'b0000000000000011100100010;
    rom[60974] = 25'b0000000000000011100100011;
    rom[60975] = 25'b0000000000000011100100100;
    rom[60976] = 25'b0000000000000011100100101;
    rom[60977] = 25'b0000000000000011100100110;
    rom[60978] = 25'b0000000000000011100100111;
    rom[60979] = 25'b0000000000000011100100111;
    rom[60980] = 25'b0000000000000011100101000;
    rom[60981] = 25'b0000000000000011100101001;
    rom[60982] = 25'b0000000000000011100101010;
    rom[60983] = 25'b0000000000000011100101011;
    rom[60984] = 25'b0000000000000011100101100;
    rom[60985] = 25'b0000000000000011100101101;
    rom[60986] = 25'b0000000000000011100101101;
    rom[60987] = 25'b0000000000000011100101110;
    rom[60988] = 25'b0000000000000011100101111;
    rom[60989] = 25'b0000000000000011100110000;
    rom[60990] = 25'b0000000000000011100110001;
    rom[60991] = 25'b0000000000000011100110010;
    rom[60992] = 25'b0000000000000011100110011;
    rom[60993] = 25'b0000000000000011100110011;
    rom[60994] = 25'b0000000000000011100110100;
    rom[60995] = 25'b0000000000000011100110101;
    rom[60996] = 25'b0000000000000011100110110;
    rom[60997] = 25'b0000000000000011100110110;
    rom[60998] = 25'b0000000000000011100110111;
    rom[60999] = 25'b0000000000000011100111001;
    rom[61000] = 25'b0000000000000011100111001;
    rom[61001] = 25'b0000000000000011100111010;
    rom[61002] = 25'b0000000000000011100111011;
    rom[61003] = 25'b0000000000000011100111100;
    rom[61004] = 25'b0000000000000011100111100;
    rom[61005] = 25'b0000000000000011100111101;
    rom[61006] = 25'b0000000000000011100111110;
    rom[61007] = 25'b0000000000000011100111111;
    rom[61008] = 25'b0000000000000011100111111;
    rom[61009] = 25'b0000000000000011101000000;
    rom[61010] = 25'b0000000000000011101000001;
    rom[61011] = 25'b0000000000000011101000010;
    rom[61012] = 25'b0000000000000011101000010;
    rom[61013] = 25'b0000000000000011101000011;
    rom[61014] = 25'b0000000000000011101000100;
    rom[61015] = 25'b0000000000000011101000101;
    rom[61016] = 25'b0000000000000011101000101;
    rom[61017] = 25'b0000000000000011101000110;
    rom[61018] = 25'b0000000000000011101000111;
    rom[61019] = 25'b0000000000000011101001000;
    rom[61020] = 25'b0000000000000011101001000;
    rom[61021] = 25'b0000000000000011101001001;
    rom[61022] = 25'b0000000000000011101001010;
    rom[61023] = 25'b0000000000000011101001010;
    rom[61024] = 25'b0000000000000011101001011;
    rom[61025] = 25'b0000000000000011101001100;
    rom[61026] = 25'b0000000000000011101001101;
    rom[61027] = 25'b0000000000000011101001101;
    rom[61028] = 25'b0000000000000011101001110;
    rom[61029] = 25'b0000000000000011101001111;
    rom[61030] = 25'b0000000000000011101010000;
    rom[61031] = 25'b0000000000000011101010000;
    rom[61032] = 25'b0000000000000011101010001;
    rom[61033] = 25'b0000000000000011101010001;
    rom[61034] = 25'b0000000000000011101010010;
    rom[61035] = 25'b0000000000000011101010011;
    rom[61036] = 25'b0000000000000011101010011;
    rom[61037] = 25'b0000000000000011101010100;
    rom[61038] = 25'b0000000000000011101010101;
    rom[61039] = 25'b0000000000000011101010110;
    rom[61040] = 25'b0000000000000011101010110;
    rom[61041] = 25'b0000000000000011101010111;
    rom[61042] = 25'b0000000000000011101011000;
    rom[61043] = 25'b0000000000000011101011000;
    rom[61044] = 25'b0000000000000011101011001;
    rom[61045] = 25'b0000000000000011101011001;
    rom[61046] = 25'b0000000000000011101011010;
    rom[61047] = 25'b0000000000000011101011011;
    rom[61048] = 25'b0000000000000011101011100;
    rom[61049] = 25'b0000000000000011101011100;
    rom[61050] = 25'b0000000000000011101011100;
    rom[61051] = 25'b0000000000000011101011101;
    rom[61052] = 25'b0000000000000011101011110;
    rom[61053] = 25'b0000000000000011101011111;
    rom[61054] = 25'b0000000000000011101011111;
    rom[61055] = 25'b0000000000000011101100000;
    rom[61056] = 25'b0000000000000011101100000;
    rom[61057] = 25'b0000000000000011101100001;
    rom[61058] = 25'b0000000000000011101100010;
    rom[61059] = 25'b0000000000000011101100010;
    rom[61060] = 25'b0000000000000011101100011;
    rom[61061] = 25'b0000000000000011101100011;
    rom[61062] = 25'b0000000000000011101100100;
    rom[61063] = 25'b0000000000000011101100101;
    rom[61064] = 25'b0000000000000011101100101;
    rom[61065] = 25'b0000000000000011101100110;
    rom[61066] = 25'b0000000000000011101100110;
    rom[61067] = 25'b0000000000000011101100111;
    rom[61068] = 25'b0000000000000011101101000;
    rom[61069] = 25'b0000000000000011101101000;
    rom[61070] = 25'b0000000000000011101101000;
    rom[61071] = 25'b0000000000000011101101001;
    rom[61072] = 25'b0000000000000011101101010;
    rom[61073] = 25'b0000000000000011101101011;
    rom[61074] = 25'b0000000000000011101101011;
    rom[61075] = 25'b0000000000000011101101011;
    rom[61076] = 25'b0000000000000011101101100;
    rom[61077] = 25'b0000000000000011101101101;
    rom[61078] = 25'b0000000000000011101101101;
    rom[61079] = 25'b0000000000000011101101110;
    rom[61080] = 25'b0000000000000011101101110;
    rom[61081] = 25'b0000000000000011101101110;
    rom[61082] = 25'b0000000000000011101101111;
    rom[61083] = 25'b0000000000000011101110000;
    rom[61084] = 25'b0000000000000011101110001;
    rom[61085] = 25'b0000000000000011101110001;
    rom[61086] = 25'b0000000000000011101110001;
    rom[61087] = 25'b0000000000000011101110010;
    rom[61088] = 25'b0000000000000011101110010;
    rom[61089] = 25'b0000000000000011101110011;
    rom[61090] = 25'b0000000000000011101110100;
    rom[61091] = 25'b0000000000000011101110100;
    rom[61092] = 25'b0000000000000011101110100;
    rom[61093] = 25'b0000000000000011101110101;
    rom[61094] = 25'b0000000000000011101110101;
    rom[61095] = 25'b0000000000000011101110110;
    rom[61096] = 25'b0000000000000011101110111;
    rom[61097] = 25'b0000000000000011101110111;
    rom[61098] = 25'b0000000000000011101110111;
    rom[61099] = 25'b0000000000000011101110111;
    rom[61100] = 25'b0000000000000011101111000;
    rom[61101] = 25'b0000000000000011101111001;
    rom[61102] = 25'b0000000000000011101111001;
    rom[61103] = 25'b0000000000000011101111010;
    rom[61104] = 25'b0000000000000011101111010;
    rom[61105] = 25'b0000000000000011101111010;
    rom[61106] = 25'b0000000000000011101111011;
    rom[61107] = 25'b0000000000000011101111011;
    rom[61108] = 25'b0000000000000011101111100;
    rom[61109] = 25'b0000000000000011101111100;
    rom[61110] = 25'b0000000000000011101111101;
    rom[61111] = 25'b0000000000000011101111101;
    rom[61112] = 25'b0000000000000011101111101;
    rom[61113] = 25'b0000000000000011101111110;
    rom[61114] = 25'b0000000000000011101111110;
    rom[61115] = 25'b0000000000000011101111111;
    rom[61116] = 25'b0000000000000011101111111;
    rom[61117] = 25'b0000000000000011110000000;
    rom[61118] = 25'b0000000000000011110000000;
    rom[61119] = 25'b0000000000000011110000000;
    rom[61120] = 25'b0000000000000011110000001;
    rom[61121] = 25'b0000000000000011110000001;
    rom[61122] = 25'b0000000000000011110000010;
    rom[61123] = 25'b0000000000000011110000010;
    rom[61124] = 25'b0000000000000011110000011;
    rom[61125] = 25'b0000000000000011110000011;
    rom[61126] = 25'b0000000000000011110000011;
    rom[61127] = 25'b0000000000000011110000011;
    rom[61128] = 25'b0000000000000011110000100;
    rom[61129] = 25'b0000000000000011110000100;
    rom[61130] = 25'b0000000000000011110000101;
    rom[61131] = 25'b0000000000000011110000101;
    rom[61132] = 25'b0000000000000011110000110;
    rom[61133] = 25'b0000000000000011110000110;
    rom[61134] = 25'b0000000000000011110000110;
    rom[61135] = 25'b0000000000000011110000110;
    rom[61136] = 25'b0000000000000011110000111;
    rom[61137] = 25'b0000000000000011110000111;
    rom[61138] = 25'b0000000000000011110001000;
    rom[61139] = 25'b0000000000000011110001000;
    rom[61140] = 25'b0000000000000011110001000;
    rom[61141] = 25'b0000000000000011110001001;
    rom[61142] = 25'b0000000000000011110001001;
    rom[61143] = 25'b0000000000000011110001001;
    rom[61144] = 25'b0000000000000011110001001;
    rom[61145] = 25'b0000000000000011110001010;
    rom[61146] = 25'b0000000000000011110001010;
    rom[61147] = 25'b0000000000000011110001010;
    rom[61148] = 25'b0000000000000011110001011;
    rom[61149] = 25'b0000000000000011110001011;
    rom[61150] = 25'b0000000000000011110001011;
    rom[61151] = 25'b0000000000000011110001011;
    rom[61152] = 25'b0000000000000011110001100;
    rom[61153] = 25'b0000000000000011110001100;
    rom[61154] = 25'b0000000000000011110001100;
    rom[61155] = 25'b0000000000000011110001101;
    rom[61156] = 25'b0000000000000011110001101;
    rom[61157] = 25'b0000000000000011110001101;
    rom[61158] = 25'b0000000000000011110001110;
    rom[61159] = 25'b0000000000000011110001110;
    rom[61160] = 25'b0000000000000011110001110;
    rom[61161] = 25'b0000000000000011110001110;
    rom[61162] = 25'b0000000000000011110001110;
    rom[61163] = 25'b0000000000000011110001111;
    rom[61164] = 25'b0000000000000011110001111;
    rom[61165] = 25'b0000000000000011110001111;
    rom[61166] = 25'b0000000000000011110010000;
    rom[61167] = 25'b0000000000000011110010000;
    rom[61168] = 25'b0000000000000011110010000;
    rom[61169] = 25'b0000000000000011110010001;
    rom[61170] = 25'b0000000000000011110010001;
    rom[61171] = 25'b0000000000000011110010001;
    rom[61172] = 25'b0000000000000011110010001;
    rom[61173] = 25'b0000000000000011110010001;
    rom[61174] = 25'b0000000000000011110010001;
    rom[61175] = 25'b0000000000000011110010010;
    rom[61176] = 25'b0000000000000011110010010;
    rom[61177] = 25'b0000000000000011110010010;
    rom[61178] = 25'b0000000000000011110010010;
    rom[61179] = 25'b0000000000000011110010011;
    rom[61180] = 25'b0000000000000011110010011;
    rom[61181] = 25'b0000000000000011110010011;
    rom[61182] = 25'b0000000000000011110010100;
    rom[61183] = 25'b0000000000000011110010100;
    rom[61184] = 25'b0000000000000011110010100;
    rom[61185] = 25'b0000000000000011110010100;
    rom[61186] = 25'b0000000000000011110010100;
    rom[61187] = 25'b0000000000000011110010100;
    rom[61188] = 25'b0000000000000011110010100;
    rom[61189] = 25'b0000000000000011110010100;
    rom[61190] = 25'b0000000000000011110010101;
    rom[61191] = 25'b0000000000000011110010101;
    rom[61192] = 25'b0000000000000011110010101;
    rom[61193] = 25'b0000000000000011110010101;
    rom[61194] = 25'b0000000000000011110010110;
    rom[61195] = 25'b0000000000000011110010110;
    rom[61196] = 25'b0000000000000011110010110;
    rom[61197] = 25'b0000000000000011110010110;
    rom[61198] = 25'b0000000000000011110010110;
    rom[61199] = 25'b0000000000000011110010111;
    rom[61200] = 25'b0000000000000011110010111;
    rom[61201] = 25'b0000000000000011110010111;
    rom[61202] = 25'b0000000000000011110010111;
    rom[61203] = 25'b0000000000000011110010111;
    rom[61204] = 25'b0000000000000011110010111;
    rom[61205] = 25'b0000000000000011110010111;
    rom[61206] = 25'b0000000000000011110010111;
    rom[61207] = 25'b0000000000000011110010111;
    rom[61208] = 25'b0000000000000011110010111;
    rom[61209] = 25'b0000000000000011110010111;
    rom[61210] = 25'b0000000000000011110011000;
    rom[61211] = 25'b0000000000000011110011000;
    rom[61212] = 25'b0000000000000011110011000;
    rom[61213] = 25'b0000000000000011110011000;
    rom[61214] = 25'b0000000000000011110011000;
    rom[61215] = 25'b0000000000000011110011000;
    rom[61216] = 25'b0000000000000011110011001;
    rom[61217] = 25'b0000000000000011110011001;
    rom[61218] = 25'b0000000000000011110011001;
    rom[61219] = 25'b0000000000000011110011001;
    rom[61220] = 25'b0000000000000011110011001;
    rom[61221] = 25'b0000000000000011110011001;
    rom[61222] = 25'b0000000000000011110011001;
    rom[61223] = 25'b0000000000000011110011001;
    rom[61224] = 25'b0000000000000011110011001;
    rom[61225] = 25'b0000000000000011110011010;
    rom[61226] = 25'b0000000000000011110011010;
    rom[61227] = 25'b0000000000000011110011010;
    rom[61228] = 25'b0000000000000011110011010;
    rom[61229] = 25'b0000000000000011110011010;
    rom[61230] = 25'b0000000000000011110011010;
    rom[61231] = 25'b0000000000000011110011010;
    rom[61232] = 25'b0000000000000011110011010;
    rom[61233] = 25'b0000000000000011110011010;
    rom[61234] = 25'b0000000000000011110011010;
    rom[61235] = 25'b0000000000000011110011010;
    rom[61236] = 25'b0000000000000011110011010;
    rom[61237] = 25'b0000000000000011110011010;
    rom[61238] = 25'b0000000000000011110011010;
    rom[61239] = 25'b0000000000000011110011010;
    rom[61240] = 25'b0000000000000011110011010;
    rom[61241] = 25'b0000000000000011110011010;
    rom[61242] = 25'b0000000000000011110011010;
    rom[61243] = 25'b0000000000000011110011010;
    rom[61244] = 25'b0000000000000011110011010;
    rom[61245] = 25'b0000000000000011110011010;
    rom[61246] = 25'b0000000000000011110011010;
    rom[61247] = 25'b0000000000000011110011010;
    rom[61248] = 25'b0000000000000011110011010;
    rom[61249] = 25'b0000000000000011110011010;
    rom[61250] = 25'b0000000000000011110011010;
    rom[61251] = 25'b0000000000000011110011010;
    rom[61252] = 25'b0000000000000011110011010;
    rom[61253] = 25'b0000000000000011110011010;
    rom[61254] = 25'b0000000000000011110011010;
    rom[61255] = 25'b0000000000000011110011010;
    rom[61256] = 25'b0000000000000011110011010;
    rom[61257] = 25'b0000000000000011110011010;
    rom[61258] = 25'b0000000000000011110011010;
    rom[61259] = 25'b0000000000000011110011010;
    rom[61260] = 25'b0000000000000011110011010;
    rom[61261] = 25'b0000000000000011110011010;
    rom[61262] = 25'b0000000000000011110011010;
    rom[61263] = 25'b0000000000000011110011010;
    rom[61264] = 25'b0000000000000011110011010;
    rom[61265] = 25'b0000000000000011110011010;
    rom[61266] = 25'b0000000000000011110011010;
    rom[61267] = 25'b0000000000000011110011010;
    rom[61268] = 25'b0000000000000011110011010;
    rom[61269] = 25'b0000000000000011110011010;
    rom[61270] = 25'b0000000000000011110011010;
    rom[61271] = 25'b0000000000000011110011010;
    rom[61272] = 25'b0000000000000011110011010;
    rom[61273] = 25'b0000000000000011110011010;
    rom[61274] = 25'b0000000000000011110011010;
    rom[61275] = 25'b0000000000000011110011010;
    rom[61276] = 25'b0000000000000011110011001;
    rom[61277] = 25'b0000000000000011110011001;
    rom[61278] = 25'b0000000000000011110011001;
    rom[61279] = 25'b0000000000000011110011001;
    rom[61280] = 25'b0000000000000011110011001;
    rom[61281] = 25'b0000000000000011110011001;
    rom[61282] = 25'b0000000000000011110011001;
    rom[61283] = 25'b0000000000000011110011001;
    rom[61284] = 25'b0000000000000011110011001;
    rom[61285] = 25'b0000000000000011110011000;
    rom[61286] = 25'b0000000000000011110011000;
    rom[61287] = 25'b0000000000000011110011000;
    rom[61288] = 25'b0000000000000011110011000;
    rom[61289] = 25'b0000000000000011110011000;
    rom[61290] = 25'b0000000000000011110011000;
    rom[61291] = 25'b0000000000000011110010111;
    rom[61292] = 25'b0000000000000011110010111;
    rom[61293] = 25'b0000000000000011110010111;
    rom[61294] = 25'b0000000000000011110010111;
    rom[61295] = 25'b0000000000000011110010111;
    rom[61296] = 25'b0000000000000011110010111;
    rom[61297] = 25'b0000000000000011110010111;
    rom[61298] = 25'b0000000000000011110010111;
    rom[61299] = 25'b0000000000000011110010111;
    rom[61300] = 25'b0000000000000011110010111;
    rom[61301] = 25'b0000000000000011110010111;
    rom[61302] = 25'b0000000000000011110010111;
    rom[61303] = 25'b0000000000000011110010110;
    rom[61304] = 25'b0000000000000011110010110;
    rom[61305] = 25'b0000000000000011110010110;
    rom[61306] = 25'b0000000000000011110010110;
    rom[61307] = 25'b0000000000000011110010101;
    rom[61308] = 25'b0000000000000011110010101;
    rom[61309] = 25'b0000000000000011110010101;
    rom[61310] = 25'b0000000000000011110010101;
    rom[61311] = 25'b0000000000000011110010101;
    rom[61312] = 25'b0000000000000011110010100;
    rom[61313] = 25'b0000000000000011110010100;
    rom[61314] = 25'b0000000000000011110010100;
    rom[61315] = 25'b0000000000000011110010100;
    rom[61316] = 25'b0000000000000011110010100;
    rom[61317] = 25'b0000000000000011110010100;
    rom[61318] = 25'b0000000000000011110010100;
    rom[61319] = 25'b0000000000000011110010100;
    rom[61320] = 25'b0000000000000011110010011;
    rom[61321] = 25'b0000000000000011110010011;
    rom[61322] = 25'b0000000000000011110010011;
    rom[61323] = 25'b0000000000000011110010010;
    rom[61324] = 25'b0000000000000011110010010;
    rom[61325] = 25'b0000000000000011110010010;
    rom[61326] = 25'b0000000000000011110010010;
    rom[61327] = 25'b0000000000000011110010001;
    rom[61328] = 25'b0000000000000011110010001;
    rom[61329] = 25'b0000000000000011110010001;
    rom[61330] = 25'b0000000000000011110010001;
    rom[61331] = 25'b0000000000000011110010001;
    rom[61332] = 25'b0000000000000011110010001;
    rom[61333] = 25'b0000000000000011110010001;
    rom[61334] = 25'b0000000000000011110010000;
    rom[61335] = 25'b0000000000000011110010000;
    rom[61336] = 25'b0000000000000011110010000;
    rom[61337] = 25'b0000000000000011110001111;
    rom[61338] = 25'b0000000000000011110001111;
    rom[61339] = 25'b0000000000000011110001111;
    rom[61340] = 25'b0000000000000011110001110;
    rom[61341] = 25'b0000000000000011110001110;
    rom[61342] = 25'b0000000000000011110001110;
    rom[61343] = 25'b0000000000000011110001110;
    rom[61344] = 25'b0000000000000011110001110;
    rom[61345] = 25'b0000000000000011110001101;
    rom[61346] = 25'b0000000000000011110001101;
    rom[61347] = 25'b0000000000000011110001101;
    rom[61348] = 25'b0000000000000011110001100;
    rom[61349] = 25'b0000000000000011110001100;
    rom[61350] = 25'b0000000000000011110001100;
    rom[61351] = 25'b0000000000000011110001011;
    rom[61352] = 25'b0000000000000011110001011;
    rom[61353] = 25'b0000000000000011110001011;
    rom[61354] = 25'b0000000000000011110001011;
    rom[61355] = 25'b0000000000000011110001011;
    rom[61356] = 25'b0000000000000011110001010;
    rom[61357] = 25'b0000000000000011110001010;
    rom[61358] = 25'b0000000000000011110001001;
    rom[61359] = 25'b0000000000000011110001001;
    rom[61360] = 25'b0000000000000011110001001;
    rom[61361] = 25'b0000000000000011110001001;
    rom[61362] = 25'b0000000000000011110001001;
    rom[61363] = 25'b0000000000000011110001000;
    rom[61364] = 25'b0000000000000011110001000;
    rom[61365] = 25'b0000000000000011110001000;
    rom[61366] = 25'b0000000000000011110000111;
    rom[61367] = 25'b0000000000000011110000111;
    rom[61368] = 25'b0000000000000011110000110;
    rom[61369] = 25'b0000000000000011110000110;
    rom[61370] = 25'b0000000000000011110000110;
    rom[61371] = 25'b0000000000000011110000110;
    rom[61372] = 25'b0000000000000011110000101;
    rom[61373] = 25'b0000000000000011110000101;
    rom[61374] = 25'b0000000000000011110000101;
    rom[61375] = 25'b0000000000000011110000100;
    rom[61376] = 25'b0000000000000011110000100;
    rom[61377] = 25'b0000000000000011110000011;
    rom[61378] = 25'b0000000000000011110000011;
    rom[61379] = 25'b0000000000000011110000011;
    rom[61380] = 25'b0000000000000011110000011;
    rom[61381] = 25'b0000000000000011110000010;
    rom[61382] = 25'b0000000000000011110000010;
    rom[61383] = 25'b0000000000000011110000001;
    rom[61384] = 25'b0000000000000011110000001;
    rom[61385] = 25'b0000000000000011110000000;
    rom[61386] = 25'b0000000000000011110000000;
    rom[61387] = 25'b0000000000000011110000000;
    rom[61388] = 25'b0000000000000011110000000;
    rom[61389] = 25'b0000000000000011101111111;
    rom[61390] = 25'b0000000000000011101111111;
    rom[61391] = 25'b0000000000000011101111110;
    rom[61392] = 25'b0000000000000011101111110;
    rom[61393] = 25'b0000000000000011101111101;
    rom[61394] = 25'b0000000000000011101111101;
    rom[61395] = 25'b0000000000000011101111101;
    rom[61396] = 25'b0000000000000011101111101;
    rom[61397] = 25'b0000000000000011101111100;
    rom[61398] = 25'b0000000000000011101111011;
    rom[61399] = 25'b0000000000000011101111011;
    rom[61400] = 25'b0000000000000011101111010;
    rom[61401] = 25'b0000000000000011101111010;
    rom[61402] = 25'b0000000000000011101111010;
    rom[61403] = 25'b0000000000000011101111010;
    rom[61404] = 25'b0000000000000011101111001;
    rom[61405] = 25'b0000000000000011101111001;
    rom[61406] = 25'b0000000000000011101111000;
    rom[61407] = 25'b0000000000000011101110111;
    rom[61408] = 25'b0000000000000011101110111;
    rom[61409] = 25'b0000000000000011101110111;
    rom[61410] = 25'b0000000000000011101110111;
    rom[61411] = 25'b0000000000000011101110110;
    rom[61412] = 25'b0000000000000011101110110;
    rom[61413] = 25'b0000000000000011101110101;
    rom[61414] = 25'b0000000000000011101110100;
    rom[61415] = 25'b0000000000000011101110100;
    rom[61416] = 25'b0000000000000011101110100;
    rom[61417] = 25'b0000000000000011101110100;
    rom[61418] = 25'b0000000000000011101110011;
    rom[61419] = 25'b0000000000000011101110010;
    rom[61420] = 25'b0000000000000011101110010;
    rom[61421] = 25'b0000000000000011101110001;
    rom[61422] = 25'b0000000000000011101110001;
    rom[61423] = 25'b0000000000000011101110001;
    rom[61424] = 25'b0000000000000011101110000;
    rom[61425] = 25'b0000000000000011101110000;
    rom[61426] = 25'b0000000000000011101101111;
    rom[61427] = 25'b0000000000000011101101110;
    rom[61428] = 25'b0000000000000011101101110;
    rom[61429] = 25'b0000000000000011101101110;
    rom[61430] = 25'b0000000000000011101101101;
    rom[61431] = 25'b0000000000000011101101101;
    rom[61432] = 25'b0000000000000011101101100;
    rom[61433] = 25'b0000000000000011101101011;
    rom[61434] = 25'b0000000000000011101101011;
    rom[61435] = 25'b0000000000000011101101011;
    rom[61436] = 25'b0000000000000011101101010;
    rom[61437] = 25'b0000000000000011101101010;
    rom[61438] = 25'b0000000000000011101101001;
    rom[61439] = 25'b0000000000000011101101000;
    rom[61440] = 25'b0000000000000011101101000;
    rom[61441] = 25'b0000000000000011101101000;
    rom[61442] = 25'b0000000000000011101100111;
    rom[61443] = 25'b0000000000000011101100111;
    rom[61444] = 25'b0000000000000011101100110;
    rom[61445] = 25'b0000000000000011101100101;
    rom[61446] = 25'b0000000000000011101100101;
    rom[61447] = 25'b0000000000000011101100101;
    rom[61448] = 25'b0000000000000011101100100;
    rom[61449] = 25'b0000000000000011101100011;
    rom[61450] = 25'b0000000000000011101100011;
    rom[61451] = 25'b0000000000000011101100010;
    rom[61452] = 25'b0000000000000011101100010;
    rom[61453] = 25'b0000000000000011101100001;
    rom[61454] = 25'b0000000000000011101100001;
    rom[61455] = 25'b0000000000000011101100000;
    rom[61456] = 25'b0000000000000011101011111;
    rom[61457] = 25'b0000000000000011101011111;
    rom[61458] = 25'b0000000000000011101011111;
    rom[61459] = 25'b0000000000000011101011110;
    rom[61460] = 25'b0000000000000011101011101;
    rom[61461] = 25'b0000000000000011101011101;
    rom[61462] = 25'b0000000000000011101011100;
    rom[61463] = 25'b0000000000000011101011100;
    rom[61464] = 25'b0000000000000011101011011;
    rom[61465] = 25'b0000000000000011101011011;
    rom[61466] = 25'b0000000000000011101011010;
    rom[61467] = 25'b0000000000000011101011001;
    rom[61468] = 25'b0000000000000011101011001;
    rom[61469] = 25'b0000000000000011101011000;
    rom[61470] = 25'b0000000000000011101011000;
    rom[61471] = 25'b0000000000000011101010111;
    rom[61472] = 25'b0000000000000011101010110;
    rom[61473] = 25'b0000000000000011101010110;
    rom[61474] = 25'b0000000000000011101010110;
    rom[61475] = 25'b0000000000000011101010101;
    rom[61476] = 25'b0000000000000011101010100;
    rom[61477] = 25'b0000000000000011101010011;
    rom[61478] = 25'b0000000000000011101010011;
    rom[61479] = 25'b0000000000000011101010011;
    rom[61480] = 25'b0000000000000011101010010;
    rom[61481] = 25'b0000000000000011101010001;
    rom[61482] = 25'b0000000000000011101010000;
    rom[61483] = 25'b0000000000000011101010000;
    rom[61484] = 25'b0000000000000011101001111;
    rom[61485] = 25'b0000000000000011101001111;
    rom[61486] = 25'b0000000000000011101001110;
    rom[61487] = 25'b0000000000000011101001101;
    rom[61488] = 25'b0000000000000011101001101;
    rom[61489] = 25'b0000000000000011101001100;
    rom[61490] = 25'b0000000000000011101001011;
    rom[61491] = 25'b0000000000000011101001011;
    rom[61492] = 25'b0000000000000011101001010;
    rom[61493] = 25'b0000000000000011101001010;
    rom[61494] = 25'b0000000000000011101001001;
    rom[61495] = 25'b0000000000000011101001000;
    rom[61496] = 25'b0000000000000011101001000;
    rom[61497] = 25'b0000000000000011101000111;
    rom[61498] = 25'b0000000000000011101000111;
    rom[61499] = 25'b0000000000000011101000110;
    rom[61500] = 25'b0000000000000011101000101;
    rom[61501] = 25'b0000000000000011101000101;
    rom[61502] = 25'b0000000000000011101000100;
    rom[61503] = 25'b0000000000000011101000011;
    rom[61504] = 25'b0000000000000011101000010;
    rom[61505] = 25'b0000000000000011101000010;
    rom[61506] = 25'b0000000000000011101000010;
    rom[61507] = 25'b0000000000000011101000001;
    rom[61508] = 25'b0000000000000011101000000;
    rom[61509] = 25'b0000000000000011100111111;
    rom[61510] = 25'b0000000000000011100111111;
    rom[61511] = 25'b0000000000000011100111110;
    rom[61512] = 25'b0000000000000011100111101;
    rom[61513] = 25'b0000000000000011100111100;
    rom[61514] = 25'b0000000000000011100111100;
    rom[61515] = 25'b0000000000000011100111011;
    rom[61516] = 25'b0000000000000011100111010;
    rom[61517] = 25'b0000000000000011100111010;
    rom[61518] = 25'b0000000000000011100111001;
    rom[61519] = 25'b0000000000000011100111001;
    rom[61520] = 25'b0000000000000011100111000;
    rom[61521] = 25'b0000000000000011100110111;
    rom[61522] = 25'b0000000000000011100110110;
    rom[61523] = 25'b0000000000000011100110110;
    rom[61524] = 25'b0000000000000011100110101;
    rom[61525] = 25'b0000000000000011100110100;
    rom[61526] = 25'b0000000000000011100110011;
    rom[61527] = 25'b0000000000000011100110011;
    rom[61528] = 25'b0000000000000011100110010;
    rom[61529] = 25'b0000000000000011100110001;
    rom[61530] = 25'b0000000000000011100110000;
    rom[61531] = 25'b0000000000000011100110000;
    rom[61532] = 25'b0000000000000011100101111;
    rom[61533] = 25'b0000000000000011100101110;
    rom[61534] = 25'b0000000000000011100101101;
    rom[61535] = 25'b0000000000000011100101101;
    rom[61536] = 25'b0000000000000011100101100;
    rom[61537] = 25'b0000000000000011100101100;
    rom[61538] = 25'b0000000000000011100101011;
    rom[61539] = 25'b0000000000000011100101010;
    rom[61540] = 25'b0000000000000011100101010;
    rom[61541] = 25'b0000000000000011100101001;
    rom[61542] = 25'b0000000000000011100101000;
    rom[61543] = 25'b0000000000000011100100111;
    rom[61544] = 25'b0000000000000011100100111;
    rom[61545] = 25'b0000000000000011100100110;
    rom[61546] = 25'b0000000000000011100100101;
    rom[61547] = 25'b0000000000000011100100100;
    rom[61548] = 25'b0000000000000011100100100;
    rom[61549] = 25'b0000000000000011100100011;
    rom[61550] = 25'b0000000000000011100100001;
    rom[61551] = 25'b0000000000000011100100001;
    rom[61552] = 25'b0000000000000011100100000;
    rom[61553] = 25'b0000000000000011100011111;
    rom[61554] = 25'b0000000000000011100011110;
    rom[61555] = 25'b0000000000000011100011110;
    rom[61556] = 25'b0000000000000011100011101;
    rom[61557] = 25'b0000000000000011100011100;
    rom[61558] = 25'b0000000000000011100011011;
    rom[61559] = 25'b0000000000000011100011011;
    rom[61560] = 25'b0000000000000011100011010;
    rom[61561] = 25'b0000000000000011100011001;
    rom[61562] = 25'b0000000000000011100011000;
    rom[61563] = 25'b0000000000000011100011000;
    rom[61564] = 25'b0000000000000011100010111;
    rom[61565] = 25'b0000000000000011100010110;
    rom[61566] = 25'b0000000000000011100010101;
    rom[61567] = 25'b0000000000000011100010101;
    rom[61568] = 25'b0000000000000011100010100;
    rom[61569] = 25'b0000000000000011100010011;
    rom[61570] = 25'b0000000000000011100010010;
    rom[61571] = 25'b0000000000000011100010001;
    rom[61572] = 25'b0000000000000011100010000;
    rom[61573] = 25'b0000000000000011100001111;
    rom[61574] = 25'b0000000000000011100001111;
    rom[61575] = 25'b0000000000000011100001110;
    rom[61576] = 25'b0000000000000011100001101;
    rom[61577] = 25'b0000000000000011100001100;
    rom[61578] = 25'b0000000000000011100001100;
    rom[61579] = 25'b0000000000000011100001011;
    rom[61580] = 25'b0000000000000011100001010;
    rom[61581] = 25'b0000000000000011100001001;
    rom[61582] = 25'b0000000000000011100001000;
    rom[61583] = 25'b0000000000000011100000111;
    rom[61584] = 25'b0000000000000011100000111;
    rom[61585] = 25'b0000000000000011100000110;
    rom[61586] = 25'b0000000000000011100000101;
    rom[61587] = 25'b0000000000000011100000100;
    rom[61588] = 25'b0000000000000011100000100;
    rom[61589] = 25'b0000000000000011100000011;
    rom[61590] = 25'b0000000000000011100000001;
    rom[61591] = 25'b0000000000000011100000001;
    rom[61592] = 25'b0000000000000011100000000;
    rom[61593] = 25'b0000000000000011011111111;
    rom[61594] = 25'b0000000000000011011111110;
    rom[61595] = 25'b0000000000000011011111110;
    rom[61596] = 25'b0000000000000011011111101;
    rom[61597] = 25'b0000000000000011011111100;
    rom[61598] = 25'b0000000000000011011111011;
    rom[61599] = 25'b0000000000000011011111010;
    rom[61600] = 25'b0000000000000011011111001;
    rom[61601] = 25'b0000000000000011011111000;
    rom[61602] = 25'b0000000000000011011111000;
    rom[61603] = 25'b0000000000000011011110111;
    rom[61604] = 25'b0000000000000011011110101;
    rom[61605] = 25'b0000000000000011011110101;
    rom[61606] = 25'b0000000000000011011110100;
    rom[61607] = 25'b0000000000000011011110011;
    rom[61608] = 25'b0000000000000011011110010;
    rom[61609] = 25'b0000000000000011011110010;
    rom[61610] = 25'b0000000000000011011110000;
    rom[61611] = 25'b0000000000000011011101111;
    rom[61612] = 25'b0000000000000011011101111;
    rom[61613] = 25'b0000000000000011011101110;
    rom[61614] = 25'b0000000000000011011101101;
    rom[61615] = 25'b0000000000000011011101100;
    rom[61616] = 25'b0000000000000011011101011;
    rom[61617] = 25'b0000000000000011011101010;
    rom[61618] = 25'b0000000000000011011101001;
    rom[61619] = 25'b0000000000000011011101001;
    rom[61620] = 25'b0000000000000011011100111;
    rom[61621] = 25'b0000000000000011011100110;
    rom[61622] = 25'b0000000000000011011100110;
    rom[61623] = 25'b0000000000000011011100101;
    rom[61624] = 25'b0000000000000011011100100;
    rom[61625] = 25'b0000000000000011011100011;
    rom[61626] = 25'b0000000000000011011100010;
    rom[61627] = 25'b0000000000000011011100001;
    rom[61628] = 25'b0000000000000011011100000;
    rom[61629] = 25'b0000000000000011011011111;
    rom[61630] = 25'b0000000000000011011011110;
    rom[61631] = 25'b0000000000000011011011101;
    rom[61632] = 25'b0000000000000011011011101;
    rom[61633] = 25'b0000000000000011011011100;
    rom[61634] = 25'b0000000000000011011011010;
    rom[61635] = 25'b0000000000000011011011010;
    rom[61636] = 25'b0000000000000011011011001;
    rom[61637] = 25'b0000000000000011011011000;
    rom[61638] = 25'b0000000000000011011010111;
    rom[61639] = 25'b0000000000000011011010110;
    rom[61640] = 25'b0000000000000011011010101;
    rom[61641] = 25'b0000000000000011011010100;
    rom[61642] = 25'b0000000000000011011010011;
    rom[61643] = 25'b0000000000000011011010010;
    rom[61644] = 25'b0000000000000011011010001;
    rom[61645] = 25'b0000000000000011011010000;
    rom[61646] = 25'b0000000000000011011001111;
    rom[61647] = 25'b0000000000000011011001110;
    rom[61648] = 25'b0000000000000011011001110;
    rom[61649] = 25'b0000000000000011011001100;
    rom[61650] = 25'b0000000000000011011001011;
    rom[61651] = 25'b0000000000000011011001011;
    rom[61652] = 25'b0000000000000011011001010;
    rom[61653] = 25'b0000000000000011011001000;
    rom[61654] = 25'b0000000000000011011001000;
    rom[61655] = 25'b0000000000000011011000111;
    rom[61656] = 25'b0000000000000011011000110;
    rom[61657] = 25'b0000000000000011011000101;
    rom[61658] = 25'b0000000000000011011000100;
    rom[61659] = 25'b0000000000000011011000011;
    rom[61660] = 25'b0000000000000011011000010;
    rom[61661] = 25'b0000000000000011011000001;
    rom[61662] = 25'b0000000000000011011000000;
    rom[61663] = 25'b0000000000000011010111111;
    rom[61664] = 25'b0000000000000011010111110;
    rom[61665] = 25'b0000000000000011010111101;
    rom[61666] = 25'b0000000000000011010111100;
    rom[61667] = 25'b0000000000000011010111011;
    rom[61668] = 25'b0000000000000011010111010;
    rom[61669] = 25'b0000000000000011010111001;
    rom[61670] = 25'b0000000000000011010111000;
    rom[61671] = 25'b0000000000000011010110111;
    rom[61672] = 25'b0000000000000011010110110;
    rom[61673] = 25'b0000000000000011010110101;
    rom[61674] = 25'b0000000000000011010110100;
    rom[61675] = 25'b0000000000000011010110011;
    rom[61676] = 25'b0000000000000011010110010;
    rom[61677] = 25'b0000000000000011010110001;
    rom[61678] = 25'b0000000000000011010110000;
    rom[61679] = 25'b0000000000000011010101111;
    rom[61680] = 25'b0000000000000011010101110;
    rom[61681] = 25'b0000000000000011010101101;
    rom[61682] = 25'b0000000000000011010101100;
    rom[61683] = 25'b0000000000000011010101011;
    rom[61684] = 25'b0000000000000011010101010;
    rom[61685] = 25'b0000000000000011010101001;
    rom[61686] = 25'b0000000000000011010101000;
    rom[61687] = 25'b0000000000000011010100111;
    rom[61688] = 25'b0000000000000011010100110;
    rom[61689] = 25'b0000000000000011010100101;
    rom[61690] = 25'b0000000000000011010100100;
    rom[61691] = 25'b0000000000000011010100011;
    rom[61692] = 25'b0000000000000011010100010;
    rom[61693] = 25'b0000000000000011010100001;
    rom[61694] = 25'b0000000000000011010011111;
    rom[61695] = 25'b0000000000000011010011111;
    rom[61696] = 25'b0000000000000011010011110;
    rom[61697] = 25'b0000000000000011010011100;
    rom[61698] = 25'b0000000000000011010011100;
    rom[61699] = 25'b0000000000000011010011010;
    rom[61700] = 25'b0000000000000011010011001;
    rom[61701] = 25'b0000000000000011010011001;
    rom[61702] = 25'b0000000000000011010010111;
    rom[61703] = 25'b0000000000000011010010110;
    rom[61704] = 25'b0000000000000011010010101;
    rom[61705] = 25'b0000000000000011010010100;
    rom[61706] = 25'b0000000000000011010010011;
    rom[61707] = 25'b0000000000000011010010010;
    rom[61708] = 25'b0000000000000011010010001;
    rom[61709] = 25'b0000000000000011010010000;
    rom[61710] = 25'b0000000000000011010001111;
    rom[61711] = 25'b0000000000000011010001110;
    rom[61712] = 25'b0000000000000011010001101;
    rom[61713] = 25'b0000000000000011010001100;
    rom[61714] = 25'b0000000000000011010001010;
    rom[61715] = 25'b0000000000000011010001010;
    rom[61716] = 25'b0000000000000011010001000;
    rom[61717] = 25'b0000000000000011010001000;
    rom[61718] = 25'b0000000000000011010000111;
    rom[61719] = 25'b0000000000000011010000101;
    rom[61720] = 25'b0000000000000011010000101;
    rom[61721] = 25'b0000000000000011010000011;
    rom[61722] = 25'b0000000000000011010000010;
    rom[61723] = 25'b0000000000000011010000001;
    rom[61724] = 25'b0000000000000011010000000;
    rom[61725] = 25'b0000000000000011001111111;
    rom[61726] = 25'b0000000000000011001111110;
    rom[61727] = 25'b0000000000000011001111100;
    rom[61728] = 25'b0000000000000011001111100;
    rom[61729] = 25'b0000000000000011001111011;
    rom[61730] = 25'b0000000000000011001111001;
    rom[61731] = 25'b0000000000000011001111001;
    rom[61732] = 25'b0000000000000011001110111;
    rom[61733] = 25'b0000000000000011001110110;
    rom[61734] = 25'b0000000000000011001110101;
    rom[61735] = 25'b0000000000000011001110100;
    rom[61736] = 25'b0000000000000011001110011;
    rom[61737] = 25'b0000000000000011001110010;
    rom[61738] = 25'b0000000000000011001110000;
    rom[61739] = 25'b0000000000000011001110000;
    rom[61740] = 25'b0000000000000011001101110;
    rom[61741] = 25'b0000000000000011001101101;
    rom[61742] = 25'b0000000000000011001101100;
    rom[61743] = 25'b0000000000000011001101011;
    rom[61744] = 25'b0000000000000011001101010;
    rom[61745] = 25'b0000000000000011001101001;
    rom[61746] = 25'b0000000000000011001100111;
    rom[61747] = 25'b0000000000000011001100111;
    rom[61748] = 25'b0000000000000011001100101;
    rom[61749] = 25'b0000000000000011001100100;
    rom[61750] = 25'b0000000000000011001100011;
    rom[61751] = 25'b0000000000000011001100010;
    rom[61752] = 25'b0000000000000011001100001;
    rom[61753] = 25'b0000000000000011001100000;
    rom[61754] = 25'b0000000000000011001011110;
    rom[61755] = 25'b0000000000000011001011110;
    rom[61756] = 25'b0000000000000011001011100;
    rom[61757] = 25'b0000000000000011001011011;
    rom[61758] = 25'b0000000000000011001011010;
    rom[61759] = 25'b0000000000000011001011001;
    rom[61760] = 25'b0000000000000011001011000;
    rom[61761] = 25'b0000000000000011001010111;
    rom[61762] = 25'b0000000000000011001010101;
    rom[61763] = 25'b0000000000000011001010101;
    rom[61764] = 25'b0000000000000011001010011;
    rom[61765] = 25'b0000000000000011001010010;
    rom[61766] = 25'b0000000000000011001010001;
    rom[61767] = 25'b0000000000000011001010000;
    rom[61768] = 25'b0000000000000011001001111;
    rom[61769] = 25'b0000000000000011001001101;
    rom[61770] = 25'b0000000000000011001001100;
    rom[61771] = 25'b0000000000000011001001011;
    rom[61772] = 25'b0000000000000011001001010;
    rom[61773] = 25'b0000000000000011001001001;
    rom[61774] = 25'b0000000000000011001001000;
    rom[61775] = 25'b0000000000000011001000111;
    rom[61776] = 25'b0000000000000011001000110;
    rom[61777] = 25'b0000000000000011001000100;
    rom[61778] = 25'b0000000000000011001000100;
    rom[61779] = 25'b0000000000000011001000010;
    rom[61780] = 25'b0000000000000011001000001;
    rom[61781] = 25'b0000000000000011001000000;
    rom[61782] = 25'b0000000000000011000111110;
    rom[61783] = 25'b0000000000000011000111110;
    rom[61784] = 25'b0000000000000011000111100;
    rom[61785] = 25'b0000000000000011000111011;
    rom[61786] = 25'b0000000000000011000111010;
    rom[61787] = 25'b0000000000000011000111000;
    rom[61788] = 25'b0000000000000011000111000;
    rom[61789] = 25'b0000000000000011000110110;
    rom[61790] = 25'b0000000000000011000110101;
    rom[61791] = 25'b0000000000000011000110100;
    rom[61792] = 25'b0000000000000011000110011;
    rom[61793] = 25'b0000000000000011000110010;
    rom[61794] = 25'b0000000000000011000110000;
    rom[61795] = 25'b0000000000000011000101111;
    rom[61796] = 25'b0000000000000011000101110;
    rom[61797] = 25'b0000000000000011000101101;
    rom[61798] = 25'b0000000000000011000101100;
    rom[61799] = 25'b0000000000000011000101010;
    rom[61800] = 25'b0000000000000011000101001;
    rom[61801] = 25'b0000000000000011000101000;
    rom[61802] = 25'b0000000000000011000100111;
    rom[61803] = 25'b0000000000000011000100110;
    rom[61804] = 25'b0000000000000011000100100;
    rom[61805] = 25'b0000000000000011000100011;
    rom[61806] = 25'b0000000000000011000100010;
    rom[61807] = 25'b0000000000000011000100001;
    rom[61808] = 25'b0000000000000011000100000;
    rom[61809] = 25'b0000000000000011000011110;
    rom[61810] = 25'b0000000000000011000011101;
    rom[61811] = 25'b0000000000000011000011100;
    rom[61812] = 25'b0000000000000011000011010;
    rom[61813] = 25'b0000000000000011000011010;
    rom[61814] = 25'b0000000000000011000011000;
    rom[61815] = 25'b0000000000000011000010111;
    rom[61816] = 25'b0000000000000011000010110;
    rom[61817] = 25'b0000000000000011000010100;
    rom[61818] = 25'b0000000000000011000010100;
    rom[61819] = 25'b0000000000000011000010010;
    rom[61820] = 25'b0000000000000011000010001;
    rom[61821] = 25'b0000000000000011000010000;
    rom[61822] = 25'b0000000000000011000001110;
    rom[61823] = 25'b0000000000000011000001110;
    rom[61824] = 25'b0000000000000011000001100;
    rom[61825] = 25'b0000000000000011000001011;
    rom[61826] = 25'b0000000000000011000001010;
    rom[61827] = 25'b0000000000000011000001000;
    rom[61828] = 25'b0000000000000011000000111;
    rom[61829] = 25'b0000000000000011000000110;
    rom[61830] = 25'b0000000000000011000000101;
    rom[61831] = 25'b0000000000000011000000011;
    rom[61832] = 25'b0000000000000011000000011;
    rom[61833] = 25'b0000000000000011000000001;
    rom[61834] = 25'b0000000000000011000000000;
    rom[61835] = 25'b0000000000000010111111111;
    rom[61836] = 25'b0000000000000010111111101;
    rom[61837] = 25'b0000000000000010111111100;
    rom[61838] = 25'b0000000000000010111111011;
    rom[61839] = 25'b0000000000000010111111010;
    rom[61840] = 25'b0000000000000010111111000;
    rom[61841] = 25'b0000000000000010111110111;
    rom[61842] = 25'b0000000000000010111110110;
    rom[61843] = 25'b0000000000000010111110100;
    rom[61844] = 25'b0000000000000010111110100;
    rom[61845] = 25'b0000000000000010111110010;
    rom[61846] = 25'b0000000000000010111110001;
    rom[61847] = 25'b0000000000000010111110000;
    rom[61848] = 25'b0000000000000010111101110;
    rom[61849] = 25'b0000000000000010111101101;
    rom[61850] = 25'b0000000000000010111101100;
    rom[61851] = 25'b0000000000000010111101011;
    rom[61852] = 25'b0000000000000010111101001;
    rom[61853] = 25'b0000000000000010111101000;
    rom[61854] = 25'b0000000000000010111100111;
    rom[61855] = 25'b0000000000000010111100101;
    rom[61856] = 25'b0000000000000010111100100;
    rom[61857] = 25'b0000000000000010111100011;
    rom[61858] = 25'b0000000000000010111100010;
    rom[61859] = 25'b0000000000000010111100000;
    rom[61860] = 25'b0000000000000010111011111;
    rom[61861] = 25'b0000000000000010111011110;
    rom[61862] = 25'b0000000000000010111011100;
    rom[61863] = 25'b0000000000000010111011100;
    rom[61864] = 25'b0000000000000010111011010;
    rom[61865] = 25'b0000000000000010111011001;
    rom[61866] = 25'b0000000000000010111010111;
    rom[61867] = 25'b0000000000000010111010110;
    rom[61868] = 25'b0000000000000010111010101;
    rom[61869] = 25'b0000000000000010111010011;
    rom[61870] = 25'b0000000000000010111010011;
    rom[61871] = 25'b0000000000000010111010001;
    rom[61872] = 25'b0000000000000010111010000;
    rom[61873] = 25'b0000000000000010111001110;
    rom[61874] = 25'b0000000000000010111001101;
    rom[61875] = 25'b0000000000000010111001100;
    rom[61876] = 25'b0000000000000010111001010;
    rom[61877] = 25'b0000000000000010111001010;
    rom[61878] = 25'b0000000000000010111001000;
    rom[61879] = 25'b0000000000000010111000111;
    rom[61880] = 25'b0000000000000010111000101;
    rom[61881] = 25'b0000000000000010111000101;
    rom[61882] = 25'b0000000000000010111000011;
    rom[61883] = 25'b0000000000000010111000010;
    rom[61884] = 25'b0000000000000010111000000;
    rom[61885] = 25'b0000000000000010110111111;
    rom[61886] = 25'b0000000000000010110111110;
    rom[61887] = 25'b0000000000000010110111100;
    rom[61888] = 25'b0000000000000010110111011;
    rom[61889] = 25'b0000000000000010110111010;
    rom[61890] = 25'b0000000000000010110111001;
    rom[61891] = 25'b0000000000000010110110111;
    rom[61892] = 25'b0000000000000010110110110;
    rom[61893] = 25'b0000000000000010110110101;
    rom[61894] = 25'b0000000000000010110110011;
    rom[61895] = 25'b0000000000000010110110010;
    rom[61896] = 25'b0000000000000010110110000;
    rom[61897] = 25'b0000000000000010110110000;
    rom[61898] = 25'b0000000000000010110101110;
    rom[61899] = 25'b0000000000000010110101101;
    rom[61900] = 25'b0000000000000010110101011;
    rom[61901] = 25'b0000000000000010110101010;
    rom[61902] = 25'b0000000000000010110101001;
    rom[61903] = 25'b0000000000000010110100111;
    rom[61904] = 25'b0000000000000010110100110;
    rom[61905] = 25'b0000000000000010110100101;
    rom[61906] = 25'b0000000000000010110100100;
    rom[61907] = 25'b0000000000000010110100010;
    rom[61908] = 25'b0000000000000010110100001;
    rom[61909] = 25'b0000000000000010110011111;
    rom[61910] = 25'b0000000000000010110011110;
    rom[61911] = 25'b0000000000000010110011101;
    rom[61912] = 25'b0000000000000010110011011;
    rom[61913] = 25'b0000000000000010110011010;
    rom[61914] = 25'b0000000000000010110011001;
    rom[61915] = 25'b0000000000000010110011000;
    rom[61916] = 25'b0000000000000010110010110;
    rom[61917] = 25'b0000000000000010110010101;
    rom[61918] = 25'b0000000000000010110010011;
    rom[61919] = 25'b0000000000000010110010010;
    rom[61920] = 25'b0000000000000010110010001;
    rom[61921] = 25'b0000000000000010110001111;
    rom[61922] = 25'b0000000000000010110001110;
    rom[61923] = 25'b0000000000000010110001101;
    rom[61924] = 25'b0000000000000010110001100;
    rom[61925] = 25'b0000000000000010110001010;
    rom[61926] = 25'b0000000000000010110001001;
    rom[61927] = 25'b0000000000000010110000111;
    rom[61928] = 25'b0000000000000010110000111;
    rom[61929] = 25'b0000000000000010110000101;
    rom[61930] = 25'b0000000000000010110000100;
    rom[61931] = 25'b0000000000000010110000010;
    rom[61932] = 25'b0000000000000010110000001;
    rom[61933] = 25'b0000000000000010110000000;
    rom[61934] = 25'b0000000000000010101111110;
    rom[61935] = 25'b0000000000000010101111101;
    rom[61936] = 25'b0000000000000010101111011;
    rom[61937] = 25'b0000000000000010101111010;
    rom[61938] = 25'b0000000000000010101111001;
    rom[61939] = 25'b0000000000000010101111000;
    rom[61940] = 25'b0000000000000010101110110;
    rom[61941] = 25'b0000000000000010101110101;
    rom[61942] = 25'b0000000000000010101110011;
    rom[61943] = 25'b0000000000000010101110010;
    rom[61944] = 25'b0000000000000010101110001;
    rom[61945] = 25'b0000000000000010101101111;
    rom[61946] = 25'b0000000000000010101101110;
    rom[61947] = 25'b0000000000000010101101100;
    rom[61948] = 25'b0000000000000010101101011;
    rom[61949] = 25'b0000000000000010101101010;
    rom[61950] = 25'b0000000000000010101101001;
    rom[61951] = 25'b0000000000000010101100111;
    rom[61952] = 25'b0000000000000010101100110;
    rom[61953] = 25'b0000000000000010101100100;
    rom[61954] = 25'b0000000000000010101100011;
    rom[61955] = 25'b0000000000000010101100010;
    rom[61956] = 25'b0000000000000010101100000;
    rom[61957] = 25'b0000000000000010101011111;
    rom[61958] = 25'b0000000000000010101011101;
    rom[61959] = 25'b0000000000000010101011100;
    rom[61960] = 25'b0000000000000010101011010;
    rom[61961] = 25'b0000000000000010101011010;
    rom[61962] = 25'b0000000000000010101011000;
    rom[61963] = 25'b0000000000000010101010111;
    rom[61964] = 25'b0000000000000010101010101;
    rom[61965] = 25'b0000000000000010101010100;
    rom[61966] = 25'b0000000000000010101010010;
    rom[61967] = 25'b0000000000000010101010001;
    rom[61968] = 25'b0000000000000010101010000;
    rom[61969] = 25'b0000000000000010101001110;
    rom[61970] = 25'b0000000000000010101001101;
    rom[61971] = 25'b0000000000000010101001011;
    rom[61972] = 25'b0000000000000010101001010;
    rom[61973] = 25'b0000000000000010101001000;
    rom[61974] = 25'b0000000000000010101001000;
    rom[61975] = 25'b0000000000000010101000110;
    rom[61976] = 25'b0000000000000010101000101;
    rom[61977] = 25'b0000000000000010101000011;
    rom[61978] = 25'b0000000000000010101000010;
    rom[61979] = 25'b0000000000000010101000000;
    rom[61980] = 25'b0000000000000010100111111;
    rom[61981] = 25'b0000000000000010100111110;
    rom[61982] = 25'b0000000000000010100111101;
    rom[61983] = 25'b0000000000000010100111011;
    rom[61984] = 25'b0000000000000010100111010;
    rom[61985] = 25'b0000000000000010100111000;
    rom[61986] = 25'b0000000000000010100110111;
    rom[61987] = 25'b0000000000000010100110101;
    rom[61988] = 25'b0000000000000010100110100;
    rom[61989] = 25'b0000000000000010100110011;
    rom[61990] = 25'b0000000000000010100110001;
    rom[61991] = 25'b0000000000000010100110000;
    rom[61992] = 25'b0000000000000010100101110;
    rom[61993] = 25'b0000000000000010100101101;
    rom[61994] = 25'b0000000000000010100101011;
    rom[61995] = 25'b0000000000000010100101010;
    rom[61996] = 25'b0000000000000010100101000;
    rom[61997] = 25'b0000000000000010100101000;
    rom[61998] = 25'b0000000000000010100100110;
    rom[61999] = 25'b0000000000000010100100101;
    rom[62000] = 25'b0000000000000010100100011;
    rom[62001] = 25'b0000000000000010100100010;
    rom[62002] = 25'b0000000000000010100100000;
    rom[62003] = 25'b0000000000000010100011111;
    rom[62004] = 25'b0000000000000010100011101;
    rom[62005] = 25'b0000000000000010100011100;
    rom[62006] = 25'b0000000000000010100011011;
    rom[62007] = 25'b0000000000000010100011001;
    rom[62008] = 25'b0000000000000010100011000;
    rom[62009] = 25'b0000000000000010100010110;
    rom[62010] = 25'b0000000000000010100010101;
    rom[62011] = 25'b0000000000000010100010011;
    rom[62012] = 25'b0000000000000010100010010;
    rom[62013] = 25'b0000000000000010100010000;
    rom[62014] = 25'b0000000000000010100010000;
    rom[62015] = 25'b0000000000000010100001110;
    rom[62016] = 25'b0000000000000010100001101;
    rom[62017] = 25'b0000000000000010100001011;
    rom[62018] = 25'b0000000000000010100001010;
    rom[62019] = 25'b0000000000000010100001000;
    rom[62020] = 25'b0000000000000010100000111;
    rom[62021] = 25'b0000000000000010100000101;
    rom[62022] = 25'b0000000000000010100000100;
    rom[62023] = 25'b0000000000000010100000010;
    rom[62024] = 25'b0000000000000010100000010;
    rom[62025] = 25'b0000000000000010100000000;
    rom[62026] = 25'b0000000000000010011111111;
    rom[62027] = 25'b0000000000000010011111101;
    rom[62028] = 25'b0000000000000010011111100;
    rom[62029] = 25'b0000000000000010011111010;
    rom[62030] = 25'b0000000000000010011111001;
    rom[62031] = 25'b0000000000000010011110111;
    rom[62032] = 25'b0000000000000010011110110;
    rom[62033] = 25'b0000000000000010011110100;
    rom[62034] = 25'b0000000000000010011110011;
    rom[62035] = 25'b0000000000000010011110010;
    rom[62036] = 25'b0000000000000010011110000;
    rom[62037] = 25'b0000000000000010011101111;
    rom[62038] = 25'b0000000000000010011101101;
    rom[62039] = 25'b0000000000000010011101100;
    rom[62040] = 25'b0000000000000010011101010;
    rom[62041] = 25'b0000000000000010011101001;
    rom[62042] = 25'b0000000000000010011100111;
    rom[62043] = 25'b0000000000000010011100110;
    rom[62044] = 25'b0000000000000010011100100;
    rom[62045] = 25'b0000000000000010011100011;
    rom[62046] = 25'b0000000000000010011100001;
    rom[62047] = 25'b0000000000000010011100000;
    rom[62048] = 25'b0000000000000010011011111;
    rom[62049] = 25'b0000000000000010011011110;
    rom[62050] = 25'b0000000000000010011011100;
    rom[62051] = 25'b0000000000000010011011011;
    rom[62052] = 25'b0000000000000010011011001;
    rom[62053] = 25'b0000000000000010011011000;
    rom[62054] = 25'b0000000000000010011010110;
    rom[62055] = 25'b0000000000000010011010101;
    rom[62056] = 25'b0000000000000010011010011;
    rom[62057] = 25'b0000000000000010011010010;
    rom[62058] = 25'b0000000000000010011010000;
    rom[62059] = 25'b0000000000000010011001111;
    rom[62060] = 25'b0000000000000010011001101;
    rom[62061] = 25'b0000000000000010011001100;
    rom[62062] = 25'b0000000000000010011001011;
    rom[62063] = 25'b0000000000000010011001001;
    rom[62064] = 25'b0000000000000010011001000;
    rom[62065] = 25'b0000000000000010011000110;
    rom[62066] = 25'b0000000000000010011000101;
    rom[62067] = 25'b0000000000000010011000100;
    rom[62068] = 25'b0000000000000010011000010;
    rom[62069] = 25'b0000000000000010011000001;
    rom[62070] = 25'b0000000000000010010111111;
    rom[62071] = 25'b0000000000000010010111110;
    rom[62072] = 25'b0000000000000010010111100;
    rom[62073] = 25'b0000000000000010010111011;
    rom[62074] = 25'b0000000000000010010111001;
    rom[62075] = 25'b0000000000000010010111000;
    rom[62076] = 25'b0000000000000010010110110;
    rom[62077] = 25'b0000000000000010010110101;
    rom[62078] = 25'b0000000000000010010110011;
    rom[62079] = 25'b0000000000000010010110010;
    rom[62080] = 25'b0000000000000010010110001;
    rom[62081] = 25'b0000000000000010010101111;
    rom[62082] = 25'b0000000000000010010101110;
    rom[62083] = 25'b0000000000000010010101100;
    rom[62084] = 25'b0000000000000010010101011;
    rom[62085] = 25'b0000000000000010010101001;
    rom[62086] = 25'b0000000000000010010101000;
    rom[62087] = 25'b0000000000000010010100110;
    rom[62088] = 25'b0000000000000010010100101;
    rom[62089] = 25'b0000000000000010010100011;
    rom[62090] = 25'b0000000000000010010100010;
    rom[62091] = 25'b0000000000000010010100000;
    rom[62092] = 25'b0000000000000010010011111;
    rom[62093] = 25'b0000000000000010010011101;
    rom[62094] = 25'b0000000000000010010011100;
    rom[62095] = 25'b0000000000000010010011010;
    rom[62096] = 25'b0000000000000010010011001;
    rom[62097] = 25'b0000000000000010010010111;
    rom[62098] = 25'b0000000000000010010010110;
    rom[62099] = 25'b0000000000000010010010100;
    rom[62100] = 25'b0000000000000010010010011;
    rom[62101] = 25'b0000000000000010010010001;
    rom[62102] = 25'b0000000000000010010010000;
    rom[62103] = 25'b0000000000000010010001111;
    rom[62104] = 25'b0000000000000010010001110;
    rom[62105] = 25'b0000000000000010010001100;
    rom[62106] = 25'b0000000000000010010001011;
    rom[62107] = 25'b0000000000000010010001001;
    rom[62108] = 25'b0000000000000010010001000;
    rom[62109] = 25'b0000000000000010010000110;
    rom[62110] = 25'b0000000000000010010000101;
    rom[62111] = 25'b0000000000000010010000011;
    rom[62112] = 25'b0000000000000010010000010;
    rom[62113] = 25'b0000000000000010010000000;
    rom[62114] = 25'b0000000000000010001111111;
    rom[62115] = 25'b0000000000000010001111101;
    rom[62116] = 25'b0000000000000010001111100;
    rom[62117] = 25'b0000000000000010001111010;
    rom[62118] = 25'b0000000000000010001111001;
    rom[62119] = 25'b0000000000000010001110111;
    rom[62120] = 25'b0000000000000010001110110;
    rom[62121] = 25'b0000000000000010001110100;
    rom[62122] = 25'b0000000000000010001110011;
    rom[62123] = 25'b0000000000000010001110001;
    rom[62124] = 25'b0000000000000010001110000;
    rom[62125] = 25'b0000000000000010001101110;
    rom[62126] = 25'b0000000000000010001101101;
    rom[62127] = 25'b0000000000000010001101011;
    rom[62128] = 25'b0000000000000010001101010;
    rom[62129] = 25'b0000000000000010001101000;
    rom[62130] = 25'b0000000000000010001100111;
    rom[62131] = 25'b0000000000000010001100101;
    rom[62132] = 25'b0000000000000010001100100;
    rom[62133] = 25'b0000000000000010001100010;
    rom[62134] = 25'b0000000000000010001100001;
    rom[62135] = 25'b0000000000000010001011111;
    rom[62136] = 25'b0000000000000010001011110;
    rom[62137] = 25'b0000000000000010001011100;
    rom[62138] = 25'b0000000000000010001011011;
    rom[62139] = 25'b0000000000000010001011001;
    rom[62140] = 25'b0000000000000010001011000;
    rom[62141] = 25'b0000000000000010001010110;
    rom[62142] = 25'b0000000000000010001010101;
    rom[62143] = 25'b0000000000000010001010011;
    rom[62144] = 25'b0000000000000010001010010;
    rom[62145] = 25'b0000000000000010001010000;
    rom[62146] = 25'b0000000000000010001010000;
    rom[62147] = 25'b0000000000000010001001110;
    rom[62148] = 25'b0000000000000010001001101;
    rom[62149] = 25'b0000000000000010001001011;
    rom[62150] = 25'b0000000000000010001001010;
    rom[62151] = 25'b0000000000000010001001000;
    rom[62152] = 25'b0000000000000010001000111;
    rom[62153] = 25'b0000000000000010001000101;
    rom[62154] = 25'b0000000000000010001000100;
    rom[62155] = 25'b0000000000000010001000010;
    rom[62156] = 25'b0000000000000010001000001;
    rom[62157] = 25'b0000000000000010000111111;
    rom[62158] = 25'b0000000000000010000111110;
    rom[62159] = 25'b0000000000000010000111100;
    rom[62160] = 25'b0000000000000010000111011;
    rom[62161] = 25'b0000000000000010000111001;
    rom[62162] = 25'b0000000000000010000111000;
    rom[62163] = 25'b0000000000000010000110110;
    rom[62164] = 25'b0000000000000010000110101;
    rom[62165] = 25'b0000000000000010000110011;
    rom[62166] = 25'b0000000000000010000110010;
    rom[62167] = 25'b0000000000000010000110000;
    rom[62168] = 25'b0000000000000010000101111;
    rom[62169] = 25'b0000000000000010000101101;
    rom[62170] = 25'b0000000000000010000101100;
    rom[62171] = 25'b0000000000000010000101010;
    rom[62172] = 25'b0000000000000010000101001;
    rom[62173] = 25'b0000000000000010000100111;
    rom[62174] = 25'b0000000000000010000100110;
    rom[62175] = 25'b0000000000000010000100100;
    rom[62176] = 25'b0000000000000010000100011;
    rom[62177] = 25'b0000000000000010000100001;
    rom[62178] = 25'b0000000000000010000100000;
    rom[62179] = 25'b0000000000000010000011110;
    rom[62180] = 25'b0000000000000010000011101;
    rom[62181] = 25'b0000000000000010000011011;
    rom[62182] = 25'b0000000000000010000011010;
    rom[62183] = 25'b0000000000000010000011000;
    rom[62184] = 25'b0000000000000010000010111;
    rom[62185] = 25'b0000000000000010000010101;
    rom[62186] = 25'b0000000000000010000010100;
    rom[62187] = 25'b0000000000000010000010010;
    rom[62188] = 25'b0000000000000010000010001;
    rom[62189] = 25'b0000000000000010000001111;
    rom[62190] = 25'b0000000000000010000001110;
    rom[62191] = 25'b0000000000000010000001100;
    rom[62192] = 25'b0000000000000010000001011;
    rom[62193] = 25'b0000000000000010000001001;
    rom[62194] = 25'b0000000000000010000001000;
    rom[62195] = 25'b0000000000000010000000110;
    rom[62196] = 25'b0000000000000010000000101;
    rom[62197] = 25'b0000000000000010000000100;
    rom[62198] = 25'b0000000000000010000000010;
    rom[62199] = 25'b0000000000000010000000001;
    rom[62200] = 25'b0000000000000001111111111;
    rom[62201] = 25'b0000000000000001111111110;
    rom[62202] = 25'b0000000000000001111111100;
    rom[62203] = 25'b0000000000000001111111011;
    rom[62204] = 25'b0000000000000001111111001;
    rom[62205] = 25'b0000000000000001111111000;
    rom[62206] = 25'b0000000000000001111110110;
    rom[62207] = 25'b0000000000000001111110101;
    rom[62208] = 25'b0000000000000001111110011;
    rom[62209] = 25'b0000000000000001111110001;
    rom[62210] = 25'b0000000000000001111101111;
    rom[62211] = 25'b0000000000000001111101110;
    rom[62212] = 25'b0000000000000001111101100;
    rom[62213] = 25'b0000000000000001111101011;
    rom[62214] = 25'b0000000000000001111101001;
    rom[62215] = 25'b0000000000000001111101000;
    rom[62216] = 25'b0000000000000001111100110;
    rom[62217] = 25'b0000000000000001111100101;
    rom[62218] = 25'b0000000000000001111100011;
    rom[62219] = 25'b0000000000000001111100010;
    rom[62220] = 25'b0000000000000001111100000;
    rom[62221] = 25'b0000000000000001111011111;
    rom[62222] = 25'b0000000000000001111011101;
    rom[62223] = 25'b0000000000000001111011100;
    rom[62224] = 25'b0000000000000001111011010;
    rom[62225] = 25'b0000000000000001111011001;
    rom[62226] = 25'b0000000000000001111010111;
    rom[62227] = 25'b0000000000000001111010110;
    rom[62228] = 25'b0000000000000001111010100;
    rom[62229] = 25'b0000000000000001111010011;
    rom[62230] = 25'b0000000000000001111010001;
    rom[62231] = 25'b0000000000000001111010000;
    rom[62232] = 25'b0000000000000001111001110;
    rom[62233] = 25'b0000000000000001111001101;
    rom[62234] = 25'b0000000000000001111001011;
    rom[62235] = 25'b0000000000000001111001010;
    rom[62236] = 25'b0000000000000001111001000;
    rom[62237] = 25'b0000000000000001111000111;
    rom[62238] = 25'b0000000000000001111000101;
    rom[62239] = 25'b0000000000000001111000100;
    rom[62240] = 25'b0000000000000001111000011;
    rom[62241] = 25'b0000000000000001111000001;
    rom[62242] = 25'b0000000000000001111000000;
    rom[62243] = 25'b0000000000000001110111110;
    rom[62244] = 25'b0000000000000001110111101;
    rom[62245] = 25'b0000000000000001110111011;
    rom[62246] = 25'b0000000000000001110111010;
    rom[62247] = 25'b0000000000000001110111000;
    rom[62248] = 25'b0000000000000001110110111;
    rom[62249] = 25'b0000000000000001110110101;
    rom[62250] = 25'b0000000000000001110110100;
    rom[62251] = 25'b0000000000000001110110010;
    rom[62252] = 25'b0000000000000001110110001;
    rom[62253] = 25'b0000000000000001110101111;
    rom[62254] = 25'b0000000000000001110101110;
    rom[62255] = 25'b0000000000000001110101100;
    rom[62256] = 25'b0000000000000001110101011;
    rom[62257] = 25'b0000000000000001110101001;
    rom[62258] = 25'b0000000000000001110101000;
    rom[62259] = 25'b0000000000000001110100110;
    rom[62260] = 25'b0000000000000001110100101;
    rom[62261] = 25'b0000000000000001110100011;
    rom[62262] = 25'b0000000000000001110100010;
    rom[62263] = 25'b0000000000000001110100000;
    rom[62264] = 25'b0000000000000001110011111;
    rom[62265] = 25'b0000000000000001110011101;
    rom[62266] = 25'b0000000000000001110011100;
    rom[62267] = 25'b0000000000000001110011010;
    rom[62268] = 25'b0000000000000001110011001;
    rom[62269] = 25'b0000000000000001110010111;
    rom[62270] = 25'b0000000000000001110010110;
    rom[62271] = 25'b0000000000000001110010100;
    rom[62272] = 25'b0000000000000001110010011;
    rom[62273] = 25'b0000000000000001110010001;
    rom[62274] = 25'b0000000000000001110010000;
    rom[62275] = 25'b0000000000000001110001110;
    rom[62276] = 25'b0000000000000001110001100;
    rom[62277] = 25'b0000000000000001110001010;
    rom[62278] = 25'b0000000000000001110001001;
    rom[62279] = 25'b0000000000000001110000111;
    rom[62280] = 25'b0000000000000001110000110;
    rom[62281] = 25'b0000000000000001110000100;
    rom[62282] = 25'b0000000000000001110000011;
    rom[62283] = 25'b0000000000000001110000010;
    rom[62284] = 25'b0000000000000001110000000;
    rom[62285] = 25'b0000000000000001101111111;
    rom[62286] = 25'b0000000000000001101111101;
    rom[62287] = 25'b0000000000000001101111100;
    rom[62288] = 25'b0000000000000001101111010;
    rom[62289] = 25'b0000000000000001101111001;
    rom[62290] = 25'b0000000000000001101110111;
    rom[62291] = 25'b0000000000000001101110110;
    rom[62292] = 25'b0000000000000001101110100;
    rom[62293] = 25'b0000000000000001101110011;
    rom[62294] = 25'b0000000000000001101110001;
    rom[62295] = 25'b0000000000000001101110000;
    rom[62296] = 25'b0000000000000001101101110;
    rom[62297] = 25'b0000000000000001101101101;
    rom[62298] = 25'b0000000000000001101101011;
    rom[62299] = 25'b0000000000000001101101010;
    rom[62300] = 25'b0000000000000001101101000;
    rom[62301] = 25'b0000000000000001101100111;
    rom[62302] = 25'b0000000000000001101100101;
    rom[62303] = 25'b0000000000000001101100100;
    rom[62304] = 25'b0000000000000001101100010;
    rom[62305] = 25'b0000000000000001101100001;
    rom[62306] = 25'b0000000000000001101011111;
    rom[62307] = 25'b0000000000000001101011110;
    rom[62308] = 25'b0000000000000001101011100;
    rom[62309] = 25'b0000000000000001101011011;
    rom[62310] = 25'b0000000000000001101011001;
    rom[62311] = 25'b0000000000000001101011000;
    rom[62312] = 25'b0000000000000001101010110;
    rom[62313] = 25'b0000000000000001101010101;
    rom[62314] = 25'b0000000000000001101010011;
    rom[62315] = 25'b0000000000000001101010010;
    rom[62316] = 25'b0000000000000001101010000;
    rom[62317] = 25'b0000000000000001101001111;
    rom[62318] = 25'b0000000000000001101001101;
    rom[62319] = 25'b0000000000000001101001100;
    rom[62320] = 25'b0000000000000001101001010;
    rom[62321] = 25'b0000000000000001101001001;
    rom[62322] = 25'b0000000000000001101000111;
    rom[62323] = 25'b0000000000000001101000110;
    rom[62324] = 25'b0000000000000001101000100;
    rom[62325] = 25'b0000000000000001101000011;
    rom[62326] = 25'b0000000000000001101000001;
    rom[62327] = 25'b0000000000000001101000000;
    rom[62328] = 25'b0000000000000001100111110;
    rom[62329] = 25'b0000000000000001100111101;
    rom[62330] = 25'b0000000000000001100111011;
    rom[62331] = 25'b0000000000000001100111010;
    rom[62332] = 25'b0000000000000001100111000;
    rom[62333] = 25'b0000000000000001100110111;
    rom[62334] = 25'b0000000000000001100110101;
    rom[62335] = 25'b0000000000000001100110100;
    rom[62336] = 25'b0000000000000001100110010;
    rom[62337] = 25'b0000000000000001100110001;
    rom[62338] = 25'b0000000000000001100101111;
    rom[62339] = 25'b0000000000000001100101101;
    rom[62340] = 25'b0000000000000001100101100;
    rom[62341] = 25'b0000000000000001100101010;
    rom[62342] = 25'b0000000000000001100101001;
    rom[62343] = 25'b0000000000000001100100111;
    rom[62344] = 25'b0000000000000001100100110;
    rom[62345] = 25'b0000000000000001100100100;
    rom[62346] = 25'b0000000000000001100100011;
    rom[62347] = 25'b0000000000000001100100001;
    rom[62348] = 25'b0000000000000001100100000;
    rom[62349] = 25'b0000000000000001100011110;
    rom[62350] = 25'b0000000000000001100011101;
    rom[62351] = 25'b0000000000000001100011011;
    rom[62352] = 25'b0000000000000001100011010;
    rom[62353] = 25'b0000000000000001100011000;
    rom[62354] = 25'b0000000000000001100010111;
    rom[62355] = 25'b0000000000000001100010101;
    rom[62356] = 25'b0000000000000001100010100;
    rom[62357] = 25'b0000000000000001100010010;
    rom[62358] = 25'b0000000000000001100010001;
    rom[62359] = 25'b0000000000000001100001111;
    rom[62360] = 25'b0000000000000001100001110;
    rom[62361] = 25'b0000000000000001100001100;
    rom[62362] = 25'b0000000000000001100001011;
    rom[62363] = 25'b0000000000000001100001001;
    rom[62364] = 25'b0000000000000001100001000;
    rom[62365] = 25'b0000000000000001100000110;
    rom[62366] = 25'b0000000000000001100000101;
    rom[62367] = 25'b0000000000000001100000011;
    rom[62368] = 25'b0000000000000001100000010;
    rom[62369] = 25'b0000000000000001100000000;
    rom[62370] = 25'b0000000000000001011111111;
    rom[62371] = 25'b0000000000000001011111101;
    rom[62372] = 25'b0000000000000001011111100;
    rom[62373] = 25'b0000000000000001011111010;
    rom[62374] = 25'b0000000000000001011111001;
    rom[62375] = 25'b0000000000000001011110111;
    rom[62376] = 25'b0000000000000001011110110;
    rom[62377] = 25'b0000000000000001011110100;
    rom[62378] = 25'b0000000000000001011110011;
    rom[62379] = 25'b0000000000000001011110001;
    rom[62380] = 25'b0000000000000001011110000;
    rom[62381] = 25'b0000000000000001011101110;
    rom[62382] = 25'b0000000000000001011101101;
    rom[62383] = 25'b0000000000000001011101011;
    rom[62384] = 25'b0000000000000001011101010;
    rom[62385] = 25'b0000000000000001011101000;
    rom[62386] = 25'b0000000000000001011100111;
    rom[62387] = 25'b0000000000000001011100101;
    rom[62388] = 25'b0000000000000001011100100;
    rom[62389] = 25'b0000000000000001011100010;
    rom[62390] = 25'b0000000000000001011100001;
    rom[62391] = 25'b0000000000000001011011111;
    rom[62392] = 25'b0000000000000001011011110;
    rom[62393] = 25'b0000000000000001011011100;
    rom[62394] = 25'b0000000000000001011011011;
    rom[62395] = 25'b0000000000000001011011001;
    rom[62396] = 25'b0000000000000001011011000;
    rom[62397] = 25'b0000000000000001011010110;
    rom[62398] = 25'b0000000000000001011010101;
    rom[62399] = 25'b0000000000000001011010011;
    rom[62400] = 25'b0000000000000001011010010;
    rom[62401] = 25'b0000000000000001011010000;
    rom[62402] = 25'b0000000000000001011001111;
    rom[62403] = 25'b0000000000000001011001101;
    rom[62404] = 25'b0000000000000001011001100;
    rom[62405] = 25'b0000000000000001011001010;
    rom[62406] = 25'b0000000000000001011001001;
    rom[62407] = 25'b0000000000000001011000111;
    rom[62408] = 25'b0000000000000001011000110;
    rom[62409] = 25'b0000000000000001011000100;
    rom[62410] = 25'b0000000000000001011000011;
    rom[62411] = 25'b0000000000000001011000010;
    rom[62412] = 25'b0000000000000001011000000;
    rom[62413] = 25'b0000000000000001010111111;
    rom[62414] = 25'b0000000000000001010111101;
    rom[62415] = 25'b0000000000000001010111100;
    rom[62416] = 25'b0000000000000001010111010;
    rom[62417] = 25'b0000000000000001010111001;
    rom[62418] = 25'b0000000000000001010110111;
    rom[62419] = 25'b0000000000000001010110110;
    rom[62420] = 25'b0000000000000001010110100;
    rom[62421] = 25'b0000000000000001010110011;
    rom[62422] = 25'b0000000000000001010110001;
    rom[62423] = 25'b0000000000000001010110000;
    rom[62424] = 25'b0000000000000001010101111;
    rom[62425] = 25'b0000000000000001010101101;
    rom[62426] = 25'b0000000000000001010101100;
    rom[62427] = 25'b0000000000000001010101010;
    rom[62428] = 25'b0000000000000001010101001;
    rom[62429] = 25'b0000000000000001010100111;
    rom[62430] = 25'b0000000000000001010100110;
    rom[62431] = 25'b0000000000000001010100100;
    rom[62432] = 25'b0000000000000001010100011;
    rom[62433] = 25'b0000000000000001010100001;
    rom[62434] = 25'b0000000000000001010100000;
    rom[62435] = 25'b0000000000000001010011110;
    rom[62436] = 25'b0000000000000001010011101;
    rom[62437] = 25'b0000000000000001010011011;
    rom[62438] = 25'b0000000000000001010011010;
    rom[62439] = 25'b0000000000000001010011000;
    rom[62440] = 25'b0000000000000001010010111;
    rom[62441] = 25'b0000000000000001010010101;
    rom[62442] = 25'b0000000000000001010010100;
    rom[62443] = 25'b0000000000000001010010010;
    rom[62444] = 25'b0000000000000001010010001;
    rom[62445] = 25'b0000000000000001010001111;
    rom[62446] = 25'b0000000000000001010001110;
    rom[62447] = 25'b0000000000000001010001100;
    rom[62448] = 25'b0000000000000001010001011;
    rom[62449] = 25'b0000000000000001010001001;
    rom[62450] = 25'b0000000000000001010001000;
    rom[62451] = 25'b0000000000000001010000110;
    rom[62452] = 25'b0000000000000001010000101;
    rom[62453] = 25'b0000000000000001010000011;
    rom[62454] = 25'b0000000000000001010000010;
    rom[62455] = 25'b0000000000000001010000001;
    rom[62456] = 25'b0000000000000001001111111;
    rom[62457] = 25'b0000000000000001001111110;
    rom[62458] = 25'b0000000000000001001111100;
    rom[62459] = 25'b0000000000000001001111011;
    rom[62460] = 25'b0000000000000001001111001;
    rom[62461] = 25'b0000000000000001001111000;
    rom[62462] = 25'b0000000000000001001110110;
    rom[62463] = 25'b0000000000000001001110101;
    rom[62464] = 25'b0000000000000001001110100;
    rom[62465] = 25'b0000000000000001001110010;
    rom[62466] = 25'b0000000000000001001110001;
    rom[62467] = 25'b0000000000000001001101111;
    rom[62468] = 25'b0000000000000001001101110;
    rom[62469] = 25'b0000000000000001001101100;
    rom[62470] = 25'b0000000000000001001101011;
    rom[62471] = 25'b0000000000000001001101001;
    rom[62472] = 25'b0000000000000001001101000;
    rom[62473] = 25'b0000000000000001001100110;
    rom[62474] = 25'b0000000000000001001100101;
    rom[62475] = 25'b0000000000000001001100011;
    rom[62476] = 25'b0000000000000001001100010;
    rom[62477] = 25'b0000000000000001001100000;
    rom[62478] = 25'b0000000000000001001011111;
    rom[62479] = 25'b0000000000000001001011101;
    rom[62480] = 25'b0000000000000001001011100;
    rom[62481] = 25'b0000000000000001001011010;
    rom[62482] = 25'b0000000000000001001011001;
    rom[62483] = 25'b0000000000000001001010111;
    rom[62484] = 25'b0000000000000001001010110;
    rom[62485] = 25'b0000000000000001001010100;
    rom[62486] = 25'b0000000000000001001010011;
    rom[62487] = 25'b0000000000000001001010010;
    rom[62488] = 25'b0000000000000001001010001;
    rom[62489] = 25'b0000000000000001001001111;
    rom[62490] = 25'b0000000000000001001001110;
    rom[62491] = 25'b0000000000000001001001100;
    rom[62492] = 25'b0000000000000001001001011;
    rom[62493] = 25'b0000000000000001001001001;
    rom[62494] = 25'b0000000000000001001001000;
    rom[62495] = 25'b0000000000000001001000110;
    rom[62496] = 25'b0000000000000001001000101;
    rom[62497] = 25'b0000000000000001001000011;
    rom[62498] = 25'b0000000000000001001000010;
    rom[62499] = 25'b0000000000000001001000000;
    rom[62500] = 25'b0000000000000001000111111;
    rom[62501] = 25'b0000000000000001000111101;
    rom[62502] = 25'b0000000000000001000111100;
    rom[62503] = 25'b0000000000000001000111010;
    rom[62504] = 25'b0000000000000001000111001;
    rom[62505] = 25'b0000000000000001000111000;
    rom[62506] = 25'b0000000000000001000110111;
    rom[62507] = 25'b0000000000000001000110101;
    rom[62508] = 25'b0000000000000001000110100;
    rom[62509] = 25'b0000000000000001000110010;
    rom[62510] = 25'b0000000000000001000110001;
    rom[62511] = 25'b0000000000000001000101111;
    rom[62512] = 25'b0000000000000001000101110;
    rom[62513] = 25'b0000000000000001000101100;
    rom[62514] = 25'b0000000000000001000101011;
    rom[62515] = 25'b0000000000000001000101001;
    rom[62516] = 25'b0000000000000001000101000;
    rom[62517] = 25'b0000000000000001000100110;
    rom[62518] = 25'b0000000000000001000100101;
    rom[62519] = 25'b0000000000000001000100011;
    rom[62520] = 25'b0000000000000001000100010;
    rom[62521] = 25'b0000000000000001000100001;
    rom[62522] = 25'b0000000000000001000011111;
    rom[62523] = 25'b0000000000000001000011110;
    rom[62524] = 25'b0000000000000001000011100;
    rom[62525] = 25'b0000000000000001000011011;
    rom[62526] = 25'b0000000000000001000011001;
    rom[62527] = 25'b0000000000000001000011000;
    rom[62528] = 25'b0000000000000001000010110;
    rom[62529] = 25'b0000000000000001000010101;
    rom[62530] = 25'b0000000000000001000010011;
    rom[62531] = 25'b0000000000000001000010010;
    rom[62532] = 25'b0000000000000001000010000;
    rom[62533] = 25'b0000000000000001000010000;
    rom[62534] = 25'b0000000000000001000001110;
    rom[62535] = 25'b0000000000000001000001101;
    rom[62536] = 25'b0000000000000001000001011;
    rom[62537] = 25'b0000000000000001000001010;
    rom[62538] = 25'b0000000000000001000001000;
    rom[62539] = 25'b0000000000000001000000111;
    rom[62540] = 25'b0000000000000001000000101;
    rom[62541] = 25'b0000000000000001000000100;
    rom[62542] = 25'b0000000000000001000000010;
    rom[62543] = 25'b0000000000000001000000001;
    rom[62544] = 25'b0000000000000000111111111;
    rom[62545] = 25'b0000000000000000111111111;
    rom[62546] = 25'b0000000000000000111111101;
    rom[62547] = 25'b0000000000000000111111100;
    rom[62548] = 25'b0000000000000000111111010;
    rom[62549] = 25'b0000000000000000111111001;
    rom[62550] = 25'b0000000000000000111110111;
    rom[62551] = 25'b0000000000000000111110110;
    rom[62552] = 25'b0000000000000000111110100;
    rom[62553] = 25'b0000000000000000111110011;
    rom[62554] = 25'b0000000000000000111110001;
    rom[62555] = 25'b0000000000000000111110000;
    rom[62556] = 25'b0000000000000000111101111;
    rom[62557] = 25'b0000000000000000111101101;
    rom[62558] = 25'b0000000000000000111101100;
    rom[62559] = 25'b0000000000000000111101010;
    rom[62560] = 25'b0000000000000000111101001;
    rom[62561] = 25'b0000000000000000111100111;
    rom[62562] = 25'b0000000000000000111100110;
    rom[62563] = 25'b0000000000000000111100100;
    rom[62564] = 25'b0000000000000000111100011;
    rom[62565] = 25'b0000000000000000111100010;
    rom[62566] = 25'b0000000000000000111100001;
    rom[62567] = 25'b0000000000000000111011111;
    rom[62568] = 25'b0000000000000000111011110;
    rom[62569] = 25'b0000000000000000111011100;
    rom[62570] = 25'b0000000000000000111011011;
    rom[62571] = 25'b0000000000000000111011001;
    rom[62572] = 25'b0000000000000000111011000;
    rom[62573] = 25'b0000000000000000111010110;
    rom[62574] = 25'b0000000000000000111010101;
    rom[62575] = 25'b0000000000000000111010100;
    rom[62576] = 25'b0000000000000000111010010;
    rom[62577] = 25'b0000000000000000111010001;
    rom[62578] = 25'b0000000000000000111001111;
    rom[62579] = 25'b0000000000000000111001110;
    rom[62580] = 25'b0000000000000000111001100;
    rom[62581] = 25'b0000000000000000111001011;
    rom[62582] = 25'b0000000000000000111001010;
    rom[62583] = 25'b0000000000000000111001001;
    rom[62584] = 25'b0000000000000000111000111;
    rom[62585] = 25'b0000000000000000111000110;
    rom[62586] = 25'b0000000000000000111000100;
    rom[62587] = 25'b0000000000000000111000011;
    rom[62588] = 25'b0000000000000000111000001;
    rom[62589] = 25'b0000000000000000111000000;
    rom[62590] = 25'b0000000000000000110111111;
    rom[62591] = 25'b0000000000000000110111110;
    rom[62592] = 25'b0000000000000000110111100;
    rom[62593] = 25'b0000000000000000110111011;
    rom[62594] = 25'b0000000000000000110111001;
    rom[62595] = 25'b0000000000000000110111000;
    rom[62596] = 25'b0000000000000000110110110;
    rom[62597] = 25'b0000000000000000110110101;
    rom[62598] = 25'b0000000000000000110110100;
    rom[62599] = 25'b0000000000000000110110010;
    rom[62600] = 25'b0000000000000000110110001;
    rom[62601] = 25'b0000000000000000110101111;
    rom[62602] = 25'b0000000000000000110101110;
    rom[62603] = 25'b0000000000000000110101100;
    rom[62604] = 25'b0000000000000000110101011;
    rom[62605] = 25'b0000000000000000110101010;
    rom[62606] = 25'b0000000000000000110101001;
    rom[62607] = 25'b0000000000000000110100111;
    rom[62608] = 25'b0000000000000000110100110;
    rom[62609] = 25'b0000000000000000110100100;
    rom[62610] = 25'b0000000000000000110100011;
    rom[62611] = 25'b0000000000000000110100001;
    rom[62612] = 25'b0000000000000000110100000;
    rom[62613] = 25'b0000000000000000110011111;
    rom[62614] = 25'b0000000000000000110011101;
    rom[62615] = 25'b0000000000000000110011100;
    rom[62616] = 25'b0000000000000000110011010;
    rom[62617] = 25'b0000000000000000110011001;
    rom[62618] = 25'b0000000000000000110010111;
    rom[62619] = 25'b0000000000000000110010111;
    rom[62620] = 25'b0000000000000000110010101;
    rom[62621] = 25'b0000000000000000110010100;
    rom[62622] = 25'b0000000000000000110010010;
    rom[62623] = 25'b0000000000000000110010001;
    rom[62624] = 25'b0000000000000000110001111;
    rom[62625] = 25'b0000000000000000110001110;
    rom[62626] = 25'b0000000000000000110001101;
    rom[62627] = 25'b0000000000000000110001011;
    rom[62628] = 25'b0000000000000000110001010;
    rom[62629] = 25'b0000000000000000110001000;
    rom[62630] = 25'b0000000000000000110000111;
    rom[62631] = 25'b0000000000000000110000110;
    rom[62632] = 25'b0000000000000000110000101;
    rom[62633] = 25'b0000000000000000110000011;
    rom[62634] = 25'b0000000000000000110000010;
    rom[62635] = 25'b0000000000000000110000000;
    rom[62636] = 25'b0000000000000000101111111;
    rom[62637] = 25'b0000000000000000101111110;
    rom[62638] = 25'b0000000000000000101111101;
    rom[62639] = 25'b0000000000000000101111011;
    rom[62640] = 25'b0000000000000000101111010;
    rom[62641] = 25'b0000000000000000101111000;
    rom[62642] = 25'b0000000000000000101110111;
    rom[62643] = 25'b0000000000000000101110110;
    rom[62644] = 25'b0000000000000000101110100;
    rom[62645] = 25'b0000000000000000101110011;
    rom[62646] = 25'b0000000000000000101110001;
    rom[62647] = 25'b0000000000000000101110000;
    rom[62648] = 25'b0000000000000000101101111;
    rom[62649] = 25'b0000000000000000101101110;
    rom[62650] = 25'b0000000000000000101101100;
    rom[62651] = 25'b0000000000000000101101011;
    rom[62652] = 25'b0000000000000000101101001;
    rom[62653] = 25'b0000000000000000101101000;
    rom[62654] = 25'b0000000000000000101100111;
    rom[62655] = 25'b0000000000000000101100101;
    rom[62656] = 25'b0000000000000000101100100;
    rom[62657] = 25'b0000000000000000101100010;
    rom[62658] = 25'b0000000000000000101100001;
    rom[62659] = 25'b0000000000000000101100000;
    rom[62660] = 25'b0000000000000000101011111;
    rom[62661] = 25'b0000000000000000101011101;
    rom[62662] = 25'b0000000000000000101011100;
    rom[62663] = 25'b0000000000000000101011010;
    rom[62664] = 25'b0000000000000000101011001;
    rom[62665] = 25'b0000000000000000101011000;
    rom[62666] = 25'b0000000000000000101010110;
    rom[62667] = 25'b0000000000000000101010101;
    rom[62668] = 25'b0000000000000000101010011;
    rom[62669] = 25'b0000000000000000101010011;
    rom[62670] = 25'b0000000000000000101010001;
    rom[62671] = 25'b0000000000000000101010000;
    rom[62672] = 25'b0000000000000000101001110;
    rom[62673] = 25'b0000000000000000101001101;
    rom[62674] = 25'b0000000000000000101001100;
    rom[62675] = 25'b0000000000000000101001010;
    rom[62676] = 25'b0000000000000000101001001;
    rom[62677] = 25'b0000000000000000101000111;
    rom[62678] = 25'b0000000000000000101000111;
    rom[62679] = 25'b0000000000000000101000101;
    rom[62680] = 25'b0000000000000000101000100;
    rom[62681] = 25'b0000000000000000101000010;
    rom[62682] = 25'b0000000000000000101000001;
    rom[62683] = 25'b0000000000000000101000000;
    rom[62684] = 25'b0000000000000000100111111;
    rom[62685] = 25'b0000000000000000100111101;
    rom[62686] = 25'b0000000000000000100111100;
    rom[62687] = 25'b0000000000000000100111011;
    rom[62688] = 25'b0000000000000000100111001;
    rom[62689] = 25'b0000000000000000100111000;
    rom[62690] = 25'b0000000000000000100110110;
    rom[62691] = 25'b0000000000000000100110101;
    rom[62692] = 25'b0000000000000000100110100;
    rom[62693] = 25'b0000000000000000100110011;
    rom[62694] = 25'b0000000000000000100110001;
    rom[62695] = 25'b0000000000000000100110000;
    rom[62696] = 25'b0000000000000000100101111;
    rom[62697] = 25'b0000000000000000100101101;
    rom[62698] = 25'b0000000000000000100101100;
    rom[62699] = 25'b0000000000000000100101010;
    rom[62700] = 25'b0000000000000000100101010;
    rom[62701] = 25'b0000000000000000100101000;
    rom[62702] = 25'b0000000000000000100100111;
    rom[62703] = 25'b0000000000000000100100101;
    rom[62704] = 25'b0000000000000000100100100;
    rom[62705] = 25'b0000000000000000100100011;
    rom[62706] = 25'b0000000000000000100100001;
    rom[62707] = 25'b0000000000000000100100000;
    rom[62708] = 25'b0000000000000000100011110;
    rom[62709] = 25'b0000000000000000100011110;
    rom[62710] = 25'b0000000000000000100011100;
    rom[62711] = 25'b0000000000000000100011011;
    rom[62712] = 25'b0000000000000000100011001;
    rom[62713] = 25'b0000000000000000100011000;
    rom[62714] = 25'b0000000000000000100010111;
    rom[62715] = 25'b0000000000000000100010101;
    rom[62716] = 25'b0000000000000000100010101;
    rom[62717] = 25'b0000000000000000100010011;
    rom[62718] = 25'b0000000000000000100010010;
    rom[62719] = 25'b0000000000000000100010000;
    rom[62720] = 25'b0000000000000000100001111;
    rom[62721] = 25'b0000000000000000100001110;
    rom[62722] = 25'b0000000000000000100001100;
    rom[62723] = 25'b0000000000000000100001011;
    rom[62724] = 25'b0000000000000000100001010;
    rom[62725] = 25'b0000000000000000100001001;
    rom[62726] = 25'b0000000000000000100000111;
    rom[62727] = 25'b0000000000000000100000110;
    rom[62728] = 25'b0000000000000000100000101;
    rom[62729] = 25'b0000000000000000100000011;
    rom[62730] = 25'b0000000000000000100000010;
    rom[62731] = 25'b0000000000000000100000001;
    rom[62732] = 25'b0000000000000000100000000;
    rom[62733] = 25'b0000000000000000011111110;
    rom[62734] = 25'b0000000000000000011111101;
    rom[62735] = 25'b0000000000000000011111100;
    rom[62736] = 25'b0000000000000000011111011;
    rom[62737] = 25'b0000000000000000011111001;
    rom[62738] = 25'b0000000000000000011111000;
    rom[62739] = 25'b0000000000000000011110111;
    rom[62740] = 25'b0000000000000000011110101;
    rom[62741] = 25'b0000000000000000011110100;
    rom[62742] = 25'b0000000000000000011110011;
    rom[62743] = 25'b0000000000000000011110010;
    rom[62744] = 25'b0000000000000000011110000;
    rom[62745] = 25'b0000000000000000011101111;
    rom[62746] = 25'b0000000000000000011101110;
    rom[62747] = 25'b0000000000000000011101100;
    rom[62748] = 25'b0000000000000000011101011;
    rom[62749] = 25'b0000000000000000011101010;
    rom[62750] = 25'b0000000000000000011101001;
    rom[62751] = 25'b0000000000000000011100111;
    rom[62752] = 25'b0000000000000000011100110;
    rom[62753] = 25'b0000000000000000011100101;
    rom[62754] = 25'b0000000000000000011100011;
    rom[62755] = 25'b0000000000000000011100010;
    rom[62756] = 25'b0000000000000000011100001;
    rom[62757] = 25'b0000000000000000011100000;
    rom[62758] = 25'b0000000000000000011011110;
    rom[62759] = 25'b0000000000000000011011101;
    rom[62760] = 25'b0000000000000000011011100;
    rom[62761] = 25'b0000000000000000011011010;
    rom[62762] = 25'b0000000000000000011011010;
    rom[62763] = 25'b0000000000000000011011000;
    rom[62764] = 25'b0000000000000000011010111;
    rom[62765] = 25'b0000000000000000011010110;
    rom[62766] = 25'b0000000000000000011010100;
    rom[62767] = 25'b0000000000000000011010011;
    rom[62768] = 25'b0000000000000000011010010;
    rom[62769] = 25'b0000000000000000011010001;
    rom[62770] = 25'b0000000000000000011001111;
    rom[62771] = 25'b0000000000000000011001110;
    rom[62772] = 25'b0000000000000000011001101;
    rom[62773] = 25'b0000000000000000011001011;
    rom[62774] = 25'b0000000000000000011001010;
    rom[62775] = 25'b0000000000000000011001001;
    rom[62776] = 25'b0000000000000000011001000;
    rom[62777] = 25'b0000000000000000011000110;
    rom[62778] = 25'b0000000000000000011000101;
    rom[62779] = 25'b0000000000000000011000100;
    rom[62780] = 25'b0000000000000000011000010;
    rom[62781] = 25'b0000000000000000011000010;
    rom[62782] = 25'b0000000000000000011000000;
    rom[62783] = 25'b0000000000000000010111111;
    rom[62784] = 25'b0000000000000000010111110;
    rom[62785] = 25'b0000000000000000010111101;
    rom[62786] = 25'b0000000000000000010111100;
    rom[62787] = 25'b0000000000000000010111010;
    rom[62788] = 25'b0000000000000000010111001;
    rom[62789] = 25'b0000000000000000010111000;
    rom[62790] = 25'b0000000000000000010110111;
    rom[62791] = 25'b0000000000000000010110101;
    rom[62792] = 25'b0000000000000000010110100;
    rom[62793] = 25'b0000000000000000010110011;
    rom[62794] = 25'b0000000000000000010110001;
    rom[62795] = 25'b0000000000000000010110001;
    rom[62796] = 25'b0000000000000000010101111;
    rom[62797] = 25'b0000000000000000010101110;
    rom[62798] = 25'b0000000000000000010101101;
    rom[62799] = 25'b0000000000000000010101011;
    rom[62800] = 25'b0000000000000000010101010;
    rom[62801] = 25'b0000000000000000010101001;
    rom[62802] = 25'b0000000000000000010101000;
    rom[62803] = 25'b0000000000000000010100111;
    rom[62804] = 25'b0000000000000000010100101;
    rom[62805] = 25'b0000000000000000010100100;
    rom[62806] = 25'b0000000000000000010100011;
    rom[62807] = 25'b0000000000000000010100010;
    rom[62808] = 25'b0000000000000000010100000;
    rom[62809] = 25'b0000000000000000010011111;
    rom[62810] = 25'b0000000000000000010011110;
    rom[62811] = 25'b0000000000000000010011100;
    rom[62812] = 25'b0000000000000000010011100;
    rom[62813] = 25'b0000000000000000010011010;
    rom[62814] = 25'b0000000000000000010011001;
    rom[62815] = 25'b0000000000000000010011000;
    rom[62816] = 25'b0000000000000000010010110;
    rom[62817] = 25'b0000000000000000010010110;
    rom[62818] = 25'b0000000000000000010010100;
    rom[62819] = 25'b0000000000000000010010011;
    rom[62820] = 25'b0000000000000000010010010;
    rom[62821] = 25'b0000000000000000010010000;
    rom[62822] = 25'b0000000000000000010010000;
    rom[62823] = 25'b0000000000000000010001110;
    rom[62824] = 25'b0000000000000000010001101;
    rom[62825] = 25'b0000000000000000010001100;
    rom[62826] = 25'b0000000000000000010001010;
    rom[62827] = 25'b0000000000000000010001010;
    rom[62828] = 25'b0000000000000000010001000;
    rom[62829] = 25'b0000000000000000010000111;
    rom[62830] = 25'b0000000000000000010000110;
    rom[62831] = 25'b0000000000000000010000100;
    rom[62832] = 25'b0000000000000000010000100;
    rom[62833] = 25'b0000000000000000010000010;
    rom[62834] = 25'b0000000000000000010000001;
    rom[62835] = 25'b0000000000000000010000000;
    rom[62836] = 25'b0000000000000000001111111;
    rom[62837] = 25'b0000000000000000001111110;
    rom[62838] = 25'b0000000000000000001111100;
    rom[62839] = 25'b0000000000000000001111100;
    rom[62840] = 25'b0000000000000000001111010;
    rom[62841] = 25'b0000000000000000001111001;
    rom[62842] = 25'b0000000000000000001111000;
    rom[62843] = 25'b0000000000000000001110110;
    rom[62844] = 25'b0000000000000000001110110;
    rom[62845] = 25'b0000000000000000001110100;
    rom[62846] = 25'b0000000000000000001110011;
    rom[62847] = 25'b0000000000000000001110010;
    rom[62848] = 25'b0000000000000000001110000;
    rom[62849] = 25'b0000000000000000001110000;
    rom[62850] = 25'b0000000000000000001101110;
    rom[62851] = 25'b0000000000000000001101101;
    rom[62852] = 25'b0000000000000000001101100;
    rom[62853] = 25'b0000000000000000001101010;
    rom[62854] = 25'b0000000000000000001101010;
    rom[62855] = 25'b0000000000000000001101000;
    rom[62856] = 25'b0000000000000000001100111;
    rom[62857] = 25'b0000000000000000001100110;
    rom[62858] = 25'b0000000000000000001100101;
    rom[62859] = 25'b0000000000000000001100100;
    rom[62860] = 25'b0000000000000000001100011;
    rom[62861] = 25'b0000000000000000001100001;
    rom[62862] = 25'b0000000000000000001100000;
    rom[62863] = 25'b0000000000000000001011111;
    rom[62864] = 25'b0000000000000000001011110;
    rom[62865] = 25'b0000000000000000001011101;
    rom[62866] = 25'b0000000000000000001011011;
    rom[62867] = 25'b0000000000000000001011011;
    rom[62868] = 25'b0000000000000000001011001;
    rom[62869] = 25'b0000000000000000001011000;
    rom[62870] = 25'b0000000000000000001010111;
    rom[62871] = 25'b0000000000000000001010101;
    rom[62872] = 25'b0000000000000000001010101;
    rom[62873] = 25'b0000000000000000001010011;
    rom[62874] = 25'b0000000000000000001010010;
    rom[62875] = 25'b0000000000000000001010001;
    rom[62876] = 25'b0000000000000000001010000;
    rom[62877] = 25'b0000000000000000001001111;
    rom[62878] = 25'b0000000000000000001001110;
    rom[62879] = 25'b0000000000000000001001100;
    rom[62880] = 25'b0000000000000000001001100;
    rom[62881] = 25'b0000000000000000001001010;
    rom[62882] = 25'b0000000000000000001001001;
    rom[62883] = 25'b0000000000000000001001000;
    rom[62884] = 25'b0000000000000000001000111;
    rom[62885] = 25'b0000000000000000001000110;
    rom[62886] = 25'b0000000000000000001000101;
    rom[62887] = 25'b0000000000000000001000011;
    rom[62888] = 25'b0000000000000000001000010;
    rom[62889] = 25'b0000000000000000001000001;
    rom[62890] = 25'b0000000000000000001000000;
    rom[62891] = 25'b0000000000000000000111111;
    rom[62892] = 25'b0000000000000000000111110;
    rom[62893] = 25'b0000000000000000000111101;
    rom[62894] = 25'b0000000000000000000111011;
    rom[62895] = 25'b0000000000000000000111011;
    rom[62896] = 25'b0000000000000000000111001;
    rom[62897] = 25'b0000000000000000000111000;
    rom[62898] = 25'b0000000000000000000110111;
    rom[62899] = 25'b0000000000000000000110110;
    rom[62900] = 25'b0000000000000000000110101;
    rom[62901] = 25'b0000000000000000000110100;
    rom[62902] = 25'b0000000000000000000110010;
    rom[62903] = 25'b0000000000000000000110010;
    rom[62904] = 25'b0000000000000000000110000;
    rom[62905] = 25'b0000000000000000000101111;
    rom[62906] = 25'b0000000000000000000101110;
    rom[62907] = 25'b0000000000000000000101101;
    rom[62908] = 25'b0000000000000000000101100;
    rom[62909] = 25'b0000000000000000000101011;
    rom[62910] = 25'b0000000000000000000101001;
    rom[62911] = 25'b0000000000000000000101001;
    rom[62912] = 25'b0000000000000000000100111;
    rom[62913] = 25'b0000000000000000000100110;
    rom[62914] = 25'b0000000000000000000100101;
    rom[62915] = 25'b0000000000000000000100100;
    rom[62916] = 25'b0000000000000000000100011;
    rom[62917] = 25'b0000000000000000000100010;
    rom[62918] = 25'b0000000000000000000100001;
    rom[62919] = 25'b0000000000000000000100000;
    rom[62920] = 25'b0000000000000000000011111;
    rom[62921] = 25'b0000000000000000000011101;
    rom[62922] = 25'b0000000000000000000011101;
    rom[62923] = 25'b0000000000000000000011011;
    rom[62924] = 25'b0000000000000000000011010;
    rom[62925] = 25'b0000000000000000000011001;
    rom[62926] = 25'b0000000000000000000011000;
    rom[62927] = 25'b0000000000000000000010111;
    rom[62928] = 25'b0000000000000000000010110;
    rom[62929] = 25'b0000000000000000000010100;
    rom[62930] = 25'b0000000000000000000010100;
    rom[62931] = 25'b0000000000000000000010011;
    rom[62932] = 25'b0000000000000000000010001;
    rom[62933] = 25'b0000000000000000000010001;
    rom[62934] = 25'b0000000000000000000001111;
    rom[62935] = 25'b0000000000000000000001110;
    rom[62936] = 25'b0000000000000000000001101;
    rom[62937] = 25'b0000000000000000000001100;
    rom[62938] = 25'b0000000000000000000001011;
    rom[62939] = 25'b0000000000000000000001010;
    rom[62940] = 25'b0000000000000000000001000;
    rom[62941] = 25'b0000000000000000000001000;
    rom[62942] = 25'b0000000000000000000000111;
    rom[62943] = 25'b0000000000000000000000101;
    rom[62944] = 25'b0000000000000000000000101;
    rom[62945] = 25'b0000000000000000000000011;
    rom[62946] = 25'b0000000000000000000000010;
    rom[62947] = 25'b0000000000000000000000001;
    rom[62948] = 25'b0000000000000000000000000;
    rom[62949] = 25'b0000000000000000000000000;
    rom[62950] = 25'b1111111111111111111111111;
    rom[62951] = 25'b1111111111111111111111110;
    rom[62952] = 25'b1111111111111111111111101;
    rom[62953] = 25'b1111111111111111111111100;
    rom[62954] = 25'b1111111111111111111111010;
    rom[62955] = 25'b1111111111111111111111010;
    rom[62956] = 25'b1111111111111111111111001;
    rom[62957] = 25'b1111111111111111111110111;
    rom[62958] = 25'b1111111111111111111110111;
    rom[62959] = 25'b1111111111111111111110101;
    rom[62960] = 25'b1111111111111111111110100;
    rom[62961] = 25'b1111111111111111111110100;
    rom[62962] = 25'b1111111111111111111110010;
    rom[62963] = 25'b1111111111111111111110001;
    rom[62964] = 25'b1111111111111111111110000;
    rom[62965] = 25'b1111111111111111111101111;
    rom[62966] = 25'b1111111111111111111101110;
    rom[62967] = 25'b1111111111111111111101101;
    rom[62968] = 25'b1111111111111111111101100;
    rom[62969] = 25'b1111111111111111111101011;
    rom[62970] = 25'b1111111111111111111101010;
    rom[62971] = 25'b1111111111111111111101001;
    rom[62972] = 25'b1111111111111111111101000;
    rom[62973] = 25'b1111111111111111111100111;
    rom[62974] = 25'b1111111111111111111100101;
    rom[62975] = 25'b1111111111111111111100101;
    rom[62976] = 25'b1111111111111111111100100;
    rom[62977] = 25'b1111111111111111111100010;
    rom[62978] = 25'b1111111111111111111100010;
    rom[62979] = 25'b1111111111111111111100000;
    rom[62980] = 25'b1111111111111111111011111;
    rom[62981] = 25'b1111111111111111111011111;
    rom[62982] = 25'b1111111111111111111011101;
    rom[62983] = 25'b1111111111111111111011100;
    rom[62984] = 25'b1111111111111111111011100;
    rom[62985] = 25'b1111111111111111111011010;
    rom[62986] = 25'b1111111111111111111011001;
    rom[62987] = 25'b1111111111111111111011000;
    rom[62988] = 25'b1111111111111111111010111;
    rom[62989] = 25'b1111111111111111111010110;
    rom[62990] = 25'b1111111111111111111010101;
    rom[62991] = 25'b1111111111111111111010100;
    rom[62992] = 25'b1111111111111111111010011;
    rom[62993] = 25'b1111111111111111111010010;
    rom[62994] = 25'b1111111111111111111010001;
    rom[62995] = 25'b1111111111111111111010000;
    rom[62996] = 25'b1111111111111111111001111;
    rom[62997] = 25'b1111111111111111111001110;
    rom[62998] = 25'b1111111111111111111001101;
    rom[62999] = 25'b1111111111111111111001100;
    rom[63000] = 25'b1111111111111111111001011;
    rom[63001] = 25'b1111111111111111111001010;
    rom[63002] = 25'b1111111111111111111001001;
    rom[63003] = 25'b1111111111111111111001000;
    rom[63004] = 25'b1111111111111111111000111;
    rom[63005] = 25'b1111111111111111111000110;
    rom[63006] = 25'b1111111111111111111000101;
    rom[63007] = 25'b1111111111111111111000100;
    rom[63008] = 25'b1111111111111111111000011;
    rom[63009] = 25'b1111111111111111111000010;
    rom[63010] = 25'b1111111111111111111000001;
    rom[63011] = 25'b1111111111111111111000000;
    rom[63012] = 25'b1111111111111111110111111;
    rom[63013] = 25'b1111111111111111110111110;
    rom[63014] = 25'b1111111111111111110111101;
    rom[63015] = 25'b1111111111111111110111100;
    rom[63016] = 25'b1111111111111111110111011;
    rom[63017] = 25'b1111111111111111110111010;
    rom[63018] = 25'b1111111111111111110111001;
    rom[63019] = 25'b1111111111111111110111000;
    rom[63020] = 25'b1111111111111111110110111;
    rom[63021] = 25'b1111111111111111110110110;
    rom[63022] = 25'b1111111111111111110110101;
    rom[63023] = 25'b1111111111111111110110100;
    rom[63024] = 25'b1111111111111111110110011;
    rom[63025] = 25'b1111111111111111110110010;
    rom[63026] = 25'b1111111111111111110110001;
    rom[63027] = 25'b1111111111111111110110000;
    rom[63028] = 25'b1111111111111111110110000;
    rom[63029] = 25'b1111111111111111110101110;
    rom[63030] = 25'b1111111111111111110101101;
    rom[63031] = 25'b1111111111111111110101101;
    rom[63032] = 25'b1111111111111111110101011;
    rom[63033] = 25'b1111111111111111110101010;
    rom[63034] = 25'b1111111111111111110101010;
    rom[63035] = 25'b1111111111111111110101000;
    rom[63036] = 25'b1111111111111111110100111;
    rom[63037] = 25'b1111111111111111110100111;
    rom[63038] = 25'b1111111111111111110100110;
    rom[63039] = 25'b1111111111111111110100100;
    rom[63040] = 25'b1111111111111111110100100;
    rom[63041] = 25'b1111111111111111110100011;
    rom[63042] = 25'b1111111111111111110100001;
    rom[63043] = 25'b1111111111111111110100001;
    rom[63044] = 25'b1111111111111111110100000;
    rom[63045] = 25'b1111111111111111110011111;
    rom[63046] = 25'b1111111111111111110011110;
    rom[63047] = 25'b1111111111111111110011101;
    rom[63048] = 25'b1111111111111111110011100;
    rom[63049] = 25'b1111111111111111110011011;
    rom[63050] = 25'b1111111111111111110011010;
    rom[63051] = 25'b1111111111111111110011001;
    rom[63052] = 25'b1111111111111111110011000;
    rom[63053] = 25'b1111111111111111110010111;
    rom[63054] = 25'b1111111111111111110010110;
    rom[63055] = 25'b1111111111111111110010101;
    rom[63056] = 25'b1111111111111111110010101;
    rom[63057] = 25'b1111111111111111110010011;
    rom[63058] = 25'b1111111111111111110010010;
    rom[63059] = 25'b1111111111111111110010010;
    rom[63060] = 25'b1111111111111111110010001;
    rom[63061] = 25'b1111111111111111110001111;
    rom[63062] = 25'b1111111111111111110001111;
    rom[63063] = 25'b1111111111111111110001110;
    rom[63064] = 25'b1111111111111111110001101;
    rom[63065] = 25'b1111111111111111110001100;
    rom[63066] = 25'b1111111111111111110001011;
    rom[63067] = 25'b1111111111111111110001010;
    rom[63068] = 25'b1111111111111111110001001;
    rom[63069] = 25'b1111111111111111110001000;
    rom[63070] = 25'b1111111111111111110000111;
    rom[63071] = 25'b1111111111111111110000110;
    rom[63072] = 25'b1111111111111111110000110;
    rom[63073] = 25'b1111111111111111110000100;
    rom[63074] = 25'b1111111111111111110000011;
    rom[63075] = 25'b1111111111111111110000011;
    rom[63076] = 25'b1111111111111111110000010;
    rom[63077] = 25'b1111111111111111110000000;
    rom[63078] = 25'b1111111111111111110000000;
    rom[63079] = 25'b1111111111111111101111111;
    rom[63080] = 25'b1111111111111111101111110;
    rom[63081] = 25'b1111111111111111101111110;
    rom[63082] = 25'b1111111111111111101111100;
    rom[63083] = 25'b1111111111111111101111011;
    rom[63084] = 25'b1111111111111111101111011;
    rom[63085] = 25'b1111111111111111101111010;
    rom[63086] = 25'b1111111111111111101111000;
    rom[63087] = 25'b1111111111111111101111000;
    rom[63088] = 25'b1111111111111111101110111;
    rom[63089] = 25'b1111111111111111101110110;
    rom[63090] = 25'b1111111111111111101110101;
    rom[63091] = 25'b1111111111111111101110100;
    rom[63092] = 25'b1111111111111111101110011;
    rom[63093] = 25'b1111111111111111101110010;
    rom[63094] = 25'b1111111111111111101110010;
    rom[63095] = 25'b1111111111111111101110001;
    rom[63096] = 25'b1111111111111111101101111;
    rom[63097] = 25'b1111111111111111101101111;
    rom[63098] = 25'b1111111111111111101101110;
    rom[63099] = 25'b1111111111111111101101101;
    rom[63100] = 25'b1111111111111111101101100;
    rom[63101] = 25'b1111111111111111101101011;
    rom[63102] = 25'b1111111111111111101101010;
    rom[63103] = 25'b1111111111111111101101001;
    rom[63104] = 25'b1111111111111111101101001;
    rom[63105] = 25'b1111111111111111101101000;
    rom[63106] = 25'b1111111111111111101100110;
    rom[63107] = 25'b1111111111111111101100110;
    rom[63108] = 25'b1111111111111111101100101;
    rom[63109] = 25'b1111111111111111101100100;
    rom[63110] = 25'b1111111111111111101100011;
    rom[63111] = 25'b1111111111111111101100011;
    rom[63112] = 25'b1111111111111111101100001;
    rom[63113] = 25'b1111111111111111101100000;
    rom[63114] = 25'b1111111111111111101100000;
    rom[63115] = 25'b1111111111111111101011111;
    rom[63116] = 25'b1111111111111111101011110;
    rom[63117] = 25'b1111111111111111101011101;
    rom[63118] = 25'b1111111111111111101011100;
    rom[63119] = 25'b1111111111111111101011011;
    rom[63120] = 25'b1111111111111111101011010;
    rom[63121] = 25'b1111111111111111101011010;
    rom[63122] = 25'b1111111111111111101011001;
    rom[63123] = 25'b1111111111111111101011000;
    rom[63124] = 25'b1111111111111111101010111;
    rom[63125] = 25'b1111111111111111101010110;
    rom[63126] = 25'b1111111111111111101010101;
    rom[63127] = 25'b1111111111111111101010100;
    rom[63128] = 25'b1111111111111111101010100;
    rom[63129] = 25'b1111111111111111101010011;
    rom[63130] = 25'b1111111111111111101010010;
    rom[63131] = 25'b1111111111111111101010001;
    rom[63132] = 25'b1111111111111111101010000;
    rom[63133] = 25'b1111111111111111101001111;
    rom[63134] = 25'b1111111111111111101001110;
    rom[63135] = 25'b1111111111111111101001110;
    rom[63136] = 25'b1111111111111111101001101;
    rom[63137] = 25'b1111111111111111101001100;
    rom[63138] = 25'b1111111111111111101001011;
    rom[63139] = 25'b1111111111111111101001010;
    rom[63140] = 25'b1111111111111111101001001;
    rom[63141] = 25'b1111111111111111101001000;
    rom[63142] = 25'b1111111111111111101001000;
    rom[63143] = 25'b1111111111111111101000111;
    rom[63144] = 25'b1111111111111111101000110;
    rom[63145] = 25'b1111111111111111101000101;
    rom[63146] = 25'b1111111111111111101000101;
    rom[63147] = 25'b1111111111111111101000011;
    rom[63148] = 25'b1111111111111111101000010;
    rom[63149] = 25'b1111111111111111101000010;
    rom[63150] = 25'b1111111111111111101000001;
    rom[63151] = 25'b1111111111111111101000000;
    rom[63152] = 25'b1111111111111111100111111;
    rom[63153] = 25'b1111111111111111100111111;
    rom[63154] = 25'b1111111111111111100111110;
    rom[63155] = 25'b1111111111111111100111101;
    rom[63156] = 25'b1111111111111111100111100;
    rom[63157] = 25'b1111111111111111100111011;
    rom[63158] = 25'b1111111111111111100111010;
    rom[63159] = 25'b1111111111111111100111010;
    rom[63160] = 25'b1111111111111111100111001;
    rom[63161] = 25'b1111111111111111100111000;
    rom[63162] = 25'b1111111111111111100110111;
    rom[63163] = 25'b1111111111111111100110111;
    rom[63164] = 25'b1111111111111111100110110;
    rom[63165] = 25'b1111111111111111100110101;
    rom[63166] = 25'b1111111111111111100110100;
    rom[63167] = 25'b1111111111111111100110011;
    rom[63168] = 25'b1111111111111111100110010;
    rom[63169] = 25'b1111111111111111100110001;
    rom[63170] = 25'b1111111111111111100110001;
    rom[63171] = 25'b1111111111111111100110000;
    rom[63172] = 25'b1111111111111111100101111;
    rom[63173] = 25'b1111111111111111100101110;
    rom[63174] = 25'b1111111111111111100101110;
    rom[63175] = 25'b1111111111111111100101101;
    rom[63176] = 25'b1111111111111111100101100;
    rom[63177] = 25'b1111111111111111100101011;
    rom[63178] = 25'b1111111111111111100101011;
    rom[63179] = 25'b1111111111111111100101010;
    rom[63180] = 25'b1111111111111111100101001;
    rom[63181] = 25'b1111111111111111100101000;
    rom[63182] = 25'b1111111111111111100100111;
    rom[63183] = 25'b1111111111111111100100110;
    rom[63184] = 25'b1111111111111111100100101;
    rom[63185] = 25'b1111111111111111100100101;
    rom[63186] = 25'b1111111111111111100100100;
    rom[63187] = 25'b1111111111111111100100011;
    rom[63188] = 25'b1111111111111111100100010;
    rom[63189] = 25'b1111111111111111100100010;
    rom[63190] = 25'b1111111111111111100100001;
    rom[63191] = 25'b1111111111111111100100000;
    rom[63192] = 25'b1111111111111111100011111;
    rom[63193] = 25'b1111111111111111100011111;
    rom[63194] = 25'b1111111111111111100011110;
    rom[63195] = 25'b1111111111111111100011101;
    rom[63196] = 25'b1111111111111111100011100;
    rom[63197] = 25'b1111111111111111100011100;
    rom[63198] = 25'b1111111111111111100011011;
    rom[63199] = 25'b1111111111111111100011010;
    rom[63200] = 25'b1111111111111111100011001;
    rom[63201] = 25'b1111111111111111100011001;
    rom[63202] = 25'b1111111111111111100011000;
    rom[63203] = 25'b1111111111111111100010111;
    rom[63204] = 25'b1111111111111111100010110;
    rom[63205] = 25'b1111111111111111100010110;
    rom[63206] = 25'b1111111111111111100010101;
    rom[63207] = 25'b1111111111111111100010100;
    rom[63208] = 25'b1111111111111111100010011;
    rom[63209] = 25'b1111111111111111100010011;
    rom[63210] = 25'b1111111111111111100010010;
    rom[63211] = 25'b1111111111111111100010001;
    rom[63212] = 25'b1111111111111111100010000;
    rom[63213] = 25'b1111111111111111100001111;
    rom[63214] = 25'b1111111111111111100001110;
    rom[63215] = 25'b1111111111111111100001101;
    rom[63216] = 25'b1111111111111111100001101;
    rom[63217] = 25'b1111111111111111100001100;
    rom[63218] = 25'b1111111111111111100001011;
    rom[63219] = 25'b1111111111111111100001011;
    rom[63220] = 25'b1111111111111111100001010;
    rom[63221] = 25'b1111111111111111100001010;
    rom[63222] = 25'b1111111111111111100001001;
    rom[63223] = 25'b1111111111111111100001000;
    rom[63224] = 25'b1111111111111111100000111;
    rom[63225] = 25'b1111111111111111100000111;
    rom[63226] = 25'b1111111111111111100000110;
    rom[63227] = 25'b1111111111111111100000101;
    rom[63228] = 25'b1111111111111111100000100;
    rom[63229] = 25'b1111111111111111100000100;
    rom[63230] = 25'b1111111111111111100000011;
    rom[63231] = 25'b1111111111111111100000010;
    rom[63232] = 25'b1111111111111111100000001;
    rom[63233] = 25'b1111111111111111100000001;
    rom[63234] = 25'b1111111111111111100000000;
    rom[63235] = 25'b1111111111111111011111111;
    rom[63236] = 25'b1111111111111111011111110;
    rom[63237] = 25'b1111111111111111011111110;
    rom[63238] = 25'b1111111111111111011111101;
    rom[63239] = 25'b1111111111111111011111100;
    rom[63240] = 25'b1111111111111111011111100;
    rom[63241] = 25'b1111111111111111011111011;
    rom[63242] = 25'b1111111111111111011111010;
    rom[63243] = 25'b1111111111111111011111001;
    rom[63244] = 25'b1111111111111111011111001;
    rom[63245] = 25'b1111111111111111011111000;
    rom[63246] = 25'b1111111111111111011110111;
    rom[63247] = 25'b1111111111111111011110110;
    rom[63248] = 25'b1111111111111111011110110;
    rom[63249] = 25'b1111111111111111011110101;
    rom[63250] = 25'b1111111111111111011110100;
    rom[63251] = 25'b1111111111111111011110100;
    rom[63252] = 25'b1111111111111111011110011;
    rom[63253] = 25'b1111111111111111011110011;
    rom[63254] = 25'b1111111111111111011110010;
    rom[63255] = 25'b1111111111111111011110001;
    rom[63256] = 25'b1111111111111111011110000;
    rom[63257] = 25'b1111111111111111011110000;
    rom[63258] = 25'b1111111111111111011101111;
    rom[63259] = 25'b1111111111111111011101110;
    rom[63260] = 25'b1111111111111111011101101;
    rom[63261] = 25'b1111111111111111011101101;
    rom[63262] = 25'b1111111111111111011101100;
    rom[63263] = 25'b1111111111111111011101011;
    rom[63264] = 25'b1111111111111111011101010;
    rom[63265] = 25'b1111111111111111011101010;
    rom[63266] = 25'b1111111111111111011101010;
    rom[63267] = 25'b1111111111111111011101001;
    rom[63268] = 25'b1111111111111111011101000;
    rom[63269] = 25'b1111111111111111011100111;
    rom[63270] = 25'b1111111111111111011100111;
    rom[63271] = 25'b1111111111111111011100110;
    rom[63272] = 25'b1111111111111111011100101;
    rom[63273] = 25'b1111111111111111011100100;
    rom[63274] = 25'b1111111111111111011100100;
    rom[63275] = 25'b1111111111111111011100011;
    rom[63276] = 25'b1111111111111111011100011;
    rom[63277] = 25'b1111111111111111011100010;
    rom[63278] = 25'b1111111111111111011100001;
    rom[63279] = 25'b1111111111111111011100001;
    rom[63280] = 25'b1111111111111111011100000;
    rom[63281] = 25'b1111111111111111011011111;
    rom[63282] = 25'b1111111111111111011011110;
    rom[63283] = 25'b1111111111111111011011110;
    rom[63284] = 25'b1111111111111111011011101;
    rom[63285] = 25'b1111111111111111011011101;
    rom[63286] = 25'b1111111111111111011011100;
    rom[63287] = 25'b1111111111111111011011011;
    rom[63288] = 25'b1111111111111111011011011;
    rom[63289] = 25'b1111111111111111011011010;
    rom[63290] = 25'b1111111111111111011011001;
    rom[63291] = 25'b1111111111111111011011000;
    rom[63292] = 25'b1111111111111111011011000;
    rom[63293] = 25'b1111111111111111011010111;
    rom[63294] = 25'b1111111111111111011010111;
    rom[63295] = 25'b1111111111111111011010110;
    rom[63296] = 25'b1111111111111111011010101;
    rom[63297] = 25'b1111111111111111011010101;
    rom[63298] = 25'b1111111111111111011010100;
    rom[63299] = 25'b1111111111111111011010011;
    rom[63300] = 25'b1111111111111111011010010;
    rom[63301] = 25'b1111111111111111011010010;
    rom[63302] = 25'b1111111111111111011010010;
    rom[63303] = 25'b1111111111111111011010001;
    rom[63304] = 25'b1111111111111111011010000;
    rom[63305] = 25'b1111111111111111011001111;
    rom[63306] = 25'b1111111111111111011001111;
    rom[63307] = 25'b1111111111111111011001110;
    rom[63308] = 25'b1111111111111111011001110;
    rom[63309] = 25'b1111111111111111011001101;
    rom[63310] = 25'b1111111111111111011001100;
    rom[63311] = 25'b1111111111111111011001100;
    rom[63312] = 25'b1111111111111111011001011;
    rom[63313] = 25'b1111111111111111011001010;
    rom[63314] = 25'b1111111111111111011001010;
    rom[63315] = 25'b1111111111111111011001001;
    rom[63316] = 25'b1111111111111111011001001;
    rom[63317] = 25'b1111111111111111011001000;
    rom[63318] = 25'b1111111111111111011000111;
    rom[63319] = 25'b1111111111111111011000110;
    rom[63320] = 25'b1111111111111111011000110;
    rom[63321] = 25'b1111111111111111011000110;
    rom[63322] = 25'b1111111111111111011000101;
    rom[63323] = 25'b1111111111111111011000100;
    rom[63324] = 25'b1111111111111111011000011;
    rom[63325] = 25'b1111111111111111011000011;
    rom[63326] = 25'b1111111111111111011000011;
    rom[63327] = 25'b1111111111111111011000010;
    rom[63328] = 25'b1111111111111111011000001;
    rom[63329] = 25'b1111111111111111011000000;
    rom[63330] = 25'b1111111111111111011000000;
    rom[63331] = 25'b1111111111111111011000000;
    rom[63332] = 25'b1111111111111111010111111;
    rom[63333] = 25'b1111111111111111010111110;
    rom[63334] = 25'b1111111111111111010111110;
    rom[63335] = 25'b1111111111111111010111101;
    rom[63336] = 25'b1111111111111111010111101;
    rom[63337] = 25'b1111111111111111010111100;
    rom[63338] = 25'b1111111111111111010111011;
    rom[63339] = 25'b1111111111111111010111011;
    rom[63340] = 25'b1111111111111111010111010;
    rom[63341] = 25'b1111111111111111010111010;
    rom[63342] = 25'b1111111111111111010111001;
    rom[63343] = 25'b1111111111111111010111000;
    rom[63344] = 25'b1111111111111111010111000;
    rom[63345] = 25'b1111111111111111010110111;
    rom[63346] = 25'b1111111111111111010110111;
    rom[63347] = 25'b1111111111111111010110110;
    rom[63348] = 25'b1111111111111111010110101;
    rom[63349] = 25'b1111111111111111010110101;
    rom[63350] = 25'b1111111111111111010110101;
    rom[63351] = 25'b1111111111111111010110100;
    rom[63352] = 25'b1111111111111111010110011;
    rom[63353] = 25'b1111111111111111010110010;
    rom[63354] = 25'b1111111111111111010110010;
    rom[63355] = 25'b1111111111111111010110010;
    rom[63356] = 25'b1111111111111111010110001;
    rom[63357] = 25'b1111111111111111010110000;
    rom[63358] = 25'b1111111111111111010101111;
    rom[63359] = 25'b1111111111111111010101111;
    rom[63360] = 25'b1111111111111111010101111;
    rom[63361] = 25'b1111111111111111010101110;
    rom[63362] = 25'b1111111111111111010101101;
    rom[63363] = 25'b1111111111111111010101101;
    rom[63364] = 25'b1111111111111111010101100;
    rom[63365] = 25'b1111111111111111010101100;
    rom[63366] = 25'b1111111111111111010101011;
    rom[63367] = 25'b1111111111111111010101011;
    rom[63368] = 25'b1111111111111111010101010;
    rom[63369] = 25'b1111111111111111010101001;
    rom[63370] = 25'b1111111111111111010101001;
    rom[63371] = 25'b1111111111111111010101001;
    rom[63372] = 25'b1111111111111111010101000;
    rom[63373] = 25'b1111111111111111010100111;
    rom[63374] = 25'b1111111111111111010100110;
    rom[63375] = 25'b1111111111111111010100110;
    rom[63376] = 25'b1111111111111111010100110;
    rom[63377] = 25'b1111111111111111010100101;
    rom[63378] = 25'b1111111111111111010100101;
    rom[63379] = 25'b1111111111111111010100100;
    rom[63380] = 25'b1111111111111111010100011;
    rom[63381] = 25'b1111111111111111010100011;
    rom[63382] = 25'b1111111111111111010100011;
    rom[63383] = 25'b1111111111111111010100010;
    rom[63384] = 25'b1111111111111111010100001;
    rom[63385] = 25'b1111111111111111010100000;
    rom[63386] = 25'b1111111111111111010100000;
    rom[63387] = 25'b1111111111111111010100000;
    rom[63388] = 25'b1111111111111111010011111;
    rom[63389] = 25'b1111111111111111010011111;
    rom[63390] = 25'b1111111111111111010011110;
    rom[63391] = 25'b1111111111111111010011101;
    rom[63392] = 25'b1111111111111111010011101;
    rom[63393] = 25'b1111111111111111010011101;
    rom[63394] = 25'b1111111111111111010011100;
    rom[63395] = 25'b1111111111111111010011011;
    rom[63396] = 25'b1111111111111111010011011;
    rom[63397] = 25'b1111111111111111010011010;
    rom[63398] = 25'b1111111111111111010011010;
    rom[63399] = 25'b1111111111111111010011010;
    rom[63400] = 25'b1111111111111111010011001;
    rom[63401] = 25'b1111111111111111010011000;
    rom[63402] = 25'b1111111111111111010011000;
    rom[63403] = 25'b1111111111111111010010111;
    rom[63404] = 25'b1111111111111111010010111;
    rom[63405] = 25'b1111111111111111010010110;
    rom[63406] = 25'b1111111111111111010010110;
    rom[63407] = 25'b1111111111111111010010101;
    rom[63408] = 25'b1111111111111111010010100;
    rom[63409] = 25'b1111111111111111010010100;
    rom[63410] = 25'b1111111111111111010010100;
    rom[63411] = 25'b1111111111111111010010011;
    rom[63412] = 25'b1111111111111111010010011;
    rom[63413] = 25'b1111111111111111010010010;
    rom[63414] = 25'b1111111111111111010010001;
    rom[63415] = 25'b1111111111111111010010001;
    rom[63416] = 25'b1111111111111111010010001;
    rom[63417] = 25'b1111111111111111010010000;
    rom[63418] = 25'b1111111111111111010010000;
    rom[63419] = 25'b1111111111111111010001111;
    rom[63420] = 25'b1111111111111111010001110;
    rom[63421] = 25'b1111111111111111010001110;
    rom[63422] = 25'b1111111111111111010001110;
    rom[63423] = 25'b1111111111111111010001101;
    rom[63424] = 25'b1111111111111111010001101;
    rom[63425] = 25'b1111111111111111010001100;
    rom[63426] = 25'b1111111111111111010001011;
    rom[63427] = 25'b1111111111111111010001011;
    rom[63428] = 25'b1111111111111111010001011;
    rom[63429] = 25'b1111111111111111010001011;
    rom[63430] = 25'b1111111111111111010001010;
    rom[63431] = 25'b1111111111111111010001001;
    rom[63432] = 25'b1111111111111111010001001;
    rom[63433] = 25'b1111111111111111010001000;
    rom[63434] = 25'b1111111111111111010001000;
    rom[63435] = 25'b1111111111111111010001000;
    rom[63436] = 25'b1111111111111111010000111;
    rom[63437] = 25'b1111111111111111010000110;
    rom[63438] = 25'b1111111111111111010000110;
    rom[63439] = 25'b1111111111111111010000101;
    rom[63440] = 25'b1111111111111111010000101;
    rom[63441] = 25'b1111111111111111010000101;
    rom[63442] = 25'b1111111111111111010000100;
    rom[63443] = 25'b1111111111111111010000100;
    rom[63444] = 25'b1111111111111111010000011;
    rom[63445] = 25'b1111111111111111010000010;
    rom[63446] = 25'b1111111111111111010000010;
    rom[63447] = 25'b1111111111111111010000010;
    rom[63448] = 25'b1111111111111111010000010;
    rom[63449] = 25'b1111111111111111010000001;
    rom[63450] = 25'b1111111111111111010000000;
    rom[63451] = 25'b1111111111111111010000000;
    rom[63452] = 25'b1111111111111111001111111;
    rom[63453] = 25'b1111111111111111001111111;
    rom[63454] = 25'b1111111111111111001111111;
    rom[63455] = 25'b1111111111111111001111110;
    rom[63456] = 25'b1111111111111111001111110;
    rom[63457] = 25'b1111111111111111001111101;
    rom[63458] = 25'b1111111111111111001111101;
    rom[63459] = 25'b1111111111111111001111101;
    rom[63460] = 25'b1111111111111111001111100;
    rom[63461] = 25'b1111111111111111001111100;
    rom[63462] = 25'b1111111111111111001111011;
    rom[63463] = 25'b1111111111111111001111011;
    rom[63464] = 25'b1111111111111111001111010;
    rom[63465] = 25'b1111111111111111001111010;
    rom[63466] = 25'b1111111111111111001111010;
    rom[63467] = 25'b1111111111111111001111001;
    rom[63468] = 25'b1111111111111111001111001;
    rom[63469] = 25'b1111111111111111001111000;
    rom[63470] = 25'b1111111111111111001110111;
    rom[63471] = 25'b1111111111111111001110111;
    rom[63472] = 25'b1111111111111111001110111;
    rom[63473] = 25'b1111111111111111001110111;
    rom[63474] = 25'b1111111111111111001110110;
    rom[63475] = 25'b1111111111111111001110110;
    rom[63476] = 25'b1111111111111111001110101;
    rom[63477] = 25'b1111111111111111001110100;
    rom[63478] = 25'b1111111111111111001110100;
    rom[63479] = 25'b1111111111111111001110100;
    rom[63480] = 25'b1111111111111111001110100;
    rom[63481] = 25'b1111111111111111001110011;
    rom[63482] = 25'b1111111111111111001110011;
    rom[63483] = 25'b1111111111111111001110010;
    rom[63484] = 25'b1111111111111111001110010;
    rom[63485] = 25'b1111111111111111001110001;
    rom[63486] = 25'b1111111111111111001110001;
    rom[63487] = 25'b1111111111111111001110001;
    rom[63488] = 25'b1111111111111111001110000;
    rom[63489] = 25'b1111111111111111001110000;
    rom[63490] = 25'b1111111111111111001101111;
    rom[63491] = 25'b1111111111111111001101111;
    rom[63492] = 25'b1111111111111111001101110;
    rom[63493] = 25'b1111111111111111001101110;
    rom[63494] = 25'b1111111111111111001101110;
    rom[63495] = 25'b1111111111111111001101110;
    rom[63496] = 25'b1111111111111111001101101;
    rom[63497] = 25'b1111111111111111001101100;
    rom[63498] = 25'b1111111111111111001101100;
    rom[63499] = 25'b1111111111111111001101011;
    rom[63500] = 25'b1111111111111111001101011;
    rom[63501] = 25'b1111111111111111001101011;
    rom[63502] = 25'b1111111111111111001101011;
    rom[63503] = 25'b1111111111111111001101010;
    rom[63504] = 25'b1111111111111111001101010;
    rom[63505] = 25'b1111111111111111001101001;
    rom[63506] = 25'b1111111111111111001101001;
    rom[63507] = 25'b1111111111111111001101000;
    rom[63508] = 25'b1111111111111111001101000;
    rom[63509] = 25'b1111111111111111001101000;
    rom[63510] = 25'b1111111111111111001101000;
    rom[63511] = 25'b1111111111111111001100111;
    rom[63512] = 25'b1111111111111111001100111;
    rom[63513] = 25'b1111111111111111001100110;
    rom[63514] = 25'b1111111111111111001100110;
    rom[63515] = 25'b1111111111111111001100101;
    rom[63516] = 25'b1111111111111111001100101;
    rom[63517] = 25'b1111111111111111001100101;
    rom[63518] = 25'b1111111111111111001100101;
    rom[63519] = 25'b1111111111111111001100100;
    rom[63520] = 25'b1111111111111111001100100;
    rom[63521] = 25'b1111111111111111001100011;
    rom[63522] = 25'b1111111111111111001100011;
    rom[63523] = 25'b1111111111111111001100010;
    rom[63524] = 25'b1111111111111111001100010;
    rom[63525] = 25'b1111111111111111001100010;
    rom[63526] = 25'b1111111111111111001100010;
    rom[63527] = 25'b1111111111111111001100001;
    rom[63528] = 25'b1111111111111111001100001;
    rom[63529] = 25'b1111111111111111001100000;
    rom[63530] = 25'b1111111111111111001100000;
    rom[63531] = 25'b1111111111111111001011111;
    rom[63532] = 25'b1111111111111111001011111;
    rom[63533] = 25'b1111111111111111001011111;
    rom[63534] = 25'b1111111111111111001011111;
    rom[63535] = 25'b1111111111111111001011110;
    rom[63536] = 25'b1111111111111111001011110;
    rom[63537] = 25'b1111111111111111001011101;
    rom[63538] = 25'b1111111111111111001011101;
    rom[63539] = 25'b1111111111111111001011100;
    rom[63540] = 25'b1111111111111111001011100;
    rom[63541] = 25'b1111111111111111001011100;
    rom[63542] = 25'b1111111111111111001011100;
    rom[63543] = 25'b1111111111111111001011100;
    rom[63544] = 25'b1111111111111111001011011;
    rom[63545] = 25'b1111111111111111001011011;
    rom[63546] = 25'b1111111111111111001011010;
    rom[63547] = 25'b1111111111111111001011010;
    rom[63548] = 25'b1111111111111111001011001;
    rom[63549] = 25'b1111111111111111001011001;
    rom[63550] = 25'b1111111111111111001011001;
    rom[63551] = 25'b1111111111111111001011001;
    rom[63552] = 25'b1111111111111111001011000;
    rom[63553] = 25'b1111111111111111001011000;
    rom[63554] = 25'b1111111111111111001011000;
    rom[63555] = 25'b1111111111111111001010111;
    rom[63556] = 25'b1111111111111111001010111;
    rom[63557] = 25'b1111111111111111001010110;
    rom[63558] = 25'b1111111111111111001010110;
    rom[63559] = 25'b1111111111111111001010110;
    rom[63560] = 25'b1111111111111111001010110;
    rom[63561] = 25'b1111111111111111001010101;
    rom[63562] = 25'b1111111111111111001010101;
    rom[63563] = 25'b1111111111111111001010101;
    rom[63564] = 25'b1111111111111111001010100;
    rom[63565] = 25'b1111111111111111001010100;
    rom[63566] = 25'b1111111111111111001010011;
    rom[63567] = 25'b1111111111111111001010011;
    rom[63568] = 25'b1111111111111111001010011;
    rom[63569] = 25'b1111111111111111001010011;
    rom[63570] = 25'b1111111111111111001010011;
    rom[63571] = 25'b1111111111111111001010010;
    rom[63572] = 25'b1111111111111111001010010;
    rom[63573] = 25'b1111111111111111001010001;
    rom[63574] = 25'b1111111111111111001010001;
    rom[63575] = 25'b1111111111111111001010001;
    rom[63576] = 25'b1111111111111111001010000;
    rom[63577] = 25'b1111111111111111001010000;
    rom[63578] = 25'b1111111111111111001010000;
    rom[63579] = 25'b1111111111111111001010000;
    rom[63580] = 25'b1111111111111111001010000;
    rom[63581] = 25'b1111111111111111001001111;
    rom[63582] = 25'b1111111111111111001001111;
    rom[63583] = 25'b1111111111111111001001110;
    rom[63584] = 25'b1111111111111111001001110;
    rom[63585] = 25'b1111111111111111001001110;
    rom[63586] = 25'b1111111111111111001001101;
    rom[63587] = 25'b1111111111111111001001101;
    rom[63588] = 25'b1111111111111111001001101;
    rom[63589] = 25'b1111111111111111001001101;
    rom[63590] = 25'b1111111111111111001001101;
    rom[63591] = 25'b1111111111111111001001100;
    rom[63592] = 25'b1111111111111111001001100;
    rom[63593] = 25'b1111111111111111001001011;
    rom[63594] = 25'b1111111111111111001001011;
    rom[63595] = 25'b1111111111111111001001011;
    rom[63596] = 25'b1111111111111111001001010;
    rom[63597] = 25'b1111111111111111001001010;
    rom[63598] = 25'b1111111111111111001001010;
    rom[63599] = 25'b1111111111111111001001010;
    rom[63600] = 25'b1111111111111111001001010;
    rom[63601] = 25'b1111111111111111001001001;
    rom[63602] = 25'b1111111111111111001001001;
    rom[63603] = 25'b1111111111111111001001001;
    rom[63604] = 25'b1111111111111111001001000;
    rom[63605] = 25'b1111111111111111001001000;
    rom[63606] = 25'b1111111111111111001001000;
    rom[63607] = 25'b1111111111111111001000111;
    rom[63608] = 25'b1111111111111111001000111;
    rom[63609] = 25'b1111111111111111001000111;
    rom[63610] = 25'b1111111111111111001000111;
    rom[63611] = 25'b1111111111111111001000111;
    rom[63612] = 25'b1111111111111111001000110;
    rom[63613] = 25'b1111111111111111001000110;
    rom[63614] = 25'b1111111111111111001000110;
    rom[63615] = 25'b1111111111111111001000101;
    rom[63616] = 25'b1111111111111111001000101;
    rom[63617] = 25'b1111111111111111001000101;
    rom[63618] = 25'b1111111111111111001000100;
    rom[63619] = 25'b1111111111111111001000100;
    rom[63620] = 25'b1111111111111111001000100;
    rom[63621] = 25'b1111111111111111001000100;
    rom[63622] = 25'b1111111111111111001000100;
    rom[63623] = 25'b1111111111111111001000100;
    rom[63624] = 25'b1111111111111111001000011;
    rom[63625] = 25'b1111111111111111001000011;
    rom[63626] = 25'b1111111111111111001000011;
    rom[63627] = 25'b1111111111111111001000010;
    rom[63628] = 25'b1111111111111111001000010;
    rom[63629] = 25'b1111111111111111001000010;
    rom[63630] = 25'b1111111111111111001000001;
    rom[63631] = 25'b1111111111111111001000001;
    rom[63632] = 25'b1111111111111111001000001;
    rom[63633] = 25'b1111111111111111001000001;
    rom[63634] = 25'b1111111111111111001000001;
    rom[63635] = 25'b1111111111111111001000001;
    rom[63636] = 25'b1111111111111111001000000;
    rom[63637] = 25'b1111111111111111001000000;
    rom[63638] = 25'b1111111111111111001000000;
    rom[63639] = 25'b1111111111111111000111111;
    rom[63640] = 25'b1111111111111111000111111;
    rom[63641] = 25'b1111111111111111000111111;
    rom[63642] = 25'b1111111111111111000111110;
    rom[63643] = 25'b1111111111111111000111110;
    rom[63644] = 25'b1111111111111111000111110;
    rom[63645] = 25'b1111111111111111000111110;
    rom[63646] = 25'b1111111111111111000111110;
    rom[63647] = 25'b1111111111111111000111110;
    rom[63648] = 25'b1111111111111111000111110;
    rom[63649] = 25'b1111111111111111000111101;
    rom[63650] = 25'b1111111111111111000111101;
    rom[63651] = 25'b1111111111111111000111101;
    rom[63652] = 25'b1111111111111111000111100;
    rom[63653] = 25'b1111111111111111000111100;
    rom[63654] = 25'b1111111111111111000111100;
    rom[63655] = 25'b1111111111111111000111100;
    rom[63656] = 25'b1111111111111111000111100;
    rom[63657] = 25'b1111111111111111000111100;
    rom[63658] = 25'b1111111111111111000111100;
    rom[63659] = 25'b1111111111111111000111011;
    rom[63660] = 25'b1111111111111111000111011;
    rom[63661] = 25'b1111111111111111000111011;
    rom[63662] = 25'b1111111111111111000111011;
    rom[63663] = 25'b1111111111111111000111010;
    rom[63664] = 25'b1111111111111111000111010;
    rom[63665] = 25'b1111111111111111000111010;
    rom[63666] = 25'b1111111111111111000111001;
    rom[63667] = 25'b1111111111111111000111001;
    rom[63668] = 25'b1111111111111111000111001;
    rom[63669] = 25'b1111111111111111000111001;
    rom[63670] = 25'b1111111111111111000111001;
    rom[63671] = 25'b1111111111111111000111001;
    rom[63672] = 25'b1111111111111111000111001;
    rom[63673] = 25'b1111111111111111000111001;
    rom[63674] = 25'b1111111111111111000111000;
    rom[63675] = 25'b1111111111111111000111000;
    rom[63676] = 25'b1111111111111111000111000;
    rom[63677] = 25'b1111111111111111000110111;
    rom[63678] = 25'b1111111111111111000110111;
    rom[63679] = 25'b1111111111111111000110111;
    rom[63680] = 25'b1111111111111111000110111;
    rom[63681] = 25'b1111111111111111000110110;
    rom[63682] = 25'b1111111111111111000110110;
    rom[63683] = 25'b1111111111111111000110110;
    rom[63684] = 25'b1111111111111111000110110;
    rom[63685] = 25'b1111111111111111000110110;
    rom[63686] = 25'b1111111111111111000110110;
    rom[63687] = 25'b1111111111111111000110110;
    rom[63688] = 25'b1111111111111111000110110;
    rom[63689] = 25'b1111111111111111000110101;
    rom[63690] = 25'b1111111111111111000110101;
    rom[63691] = 25'b1111111111111111000110101;
    rom[63692] = 25'b1111111111111111000110101;
    rom[63693] = 25'b1111111111111111000110101;
    rom[63694] = 25'b1111111111111111000110100;
    rom[63695] = 25'b1111111111111111000110100;
    rom[63696] = 25'b1111111111111111000110100;
    rom[63697] = 25'b1111111111111111000110100;
    rom[63698] = 25'b1111111111111111000110011;
    rom[63699] = 25'b1111111111111111000110011;
    rom[63700] = 25'b1111111111111111000110011;
    rom[63701] = 25'b1111111111111111000110011;
    rom[63702] = 25'b1111111111111111000110011;
    rom[63703] = 25'b1111111111111111000110011;
    rom[63704] = 25'b1111111111111111000110011;
    rom[63705] = 25'b1111111111111111000110011;
    rom[63706] = 25'b1111111111111111000110011;
    rom[63707] = 25'b1111111111111111000110010;
    rom[63708] = 25'b1111111111111111000110010;
    rom[63709] = 25'b1111111111111111000110010;
    rom[63710] = 25'b1111111111111111000110010;
    rom[63711] = 25'b1111111111111111000110001;
    rom[63712] = 25'b1111111111111111000110001;
    rom[63713] = 25'b1111111111111111000110001;
    rom[63714] = 25'b1111111111111111000110001;
    rom[63715] = 25'b1111111111111111000110001;
    rom[63716] = 25'b1111111111111111000110000;
    rom[63717] = 25'b1111111111111111000110000;
    rom[63718] = 25'b1111111111111111000110000;
    rom[63719] = 25'b1111111111111111000110000;
    rom[63720] = 25'b1111111111111111000110000;
    rom[63721] = 25'b1111111111111111000110000;
    rom[63722] = 25'b1111111111111111000110000;
    rom[63723] = 25'b1111111111111111000110000;
    rom[63724] = 25'b1111111111111111000110000;
    rom[63725] = 25'b1111111111111111000110000;
    rom[63726] = 25'b1111111111111111000101111;
    rom[63727] = 25'b1111111111111111000101111;
    rom[63728] = 25'b1111111111111111000101111;
    rom[63729] = 25'b1111111111111111000101111;
    rom[63730] = 25'b1111111111111111000101111;
    rom[63731] = 25'b1111111111111111000101111;
    rom[63732] = 25'b1111111111111111000101110;
    rom[63733] = 25'b1111111111111111000101110;
    rom[63734] = 25'b1111111111111111000101110;
    rom[63735] = 25'b1111111111111111000101110;
    rom[63736] = 25'b1111111111111111000101110;
    rom[63737] = 25'b1111111111111111000101110;
    rom[63738] = 25'b1111111111111111000101101;
    rom[63739] = 25'b1111111111111111000101101;
    rom[63740] = 25'b1111111111111111000101101;
    rom[63741] = 25'b1111111111111111000101101;
    rom[63742] = 25'b1111111111111111000101101;
    rom[63743] = 25'b1111111111111111000101101;
    rom[63744] = 25'b1111111111111111000101101;
    rom[63745] = 25'b1111111111111111000101101;
    rom[63746] = 25'b1111111111111111000101101;
    rom[63747] = 25'b1111111111111111000101101;
    rom[63748] = 25'b1111111111111111000101101;
    rom[63749] = 25'b1111111111111111000101101;
    rom[63750] = 25'b1111111111111111000101100;
    rom[63751] = 25'b1111111111111111000101100;
    rom[63752] = 25'b1111111111111111000101100;
    rom[63753] = 25'b1111111111111111000101100;
    rom[63754] = 25'b1111111111111111000101100;
    rom[63755] = 25'b1111111111111111000101100;
    rom[63756] = 25'b1111111111111111000101011;
    rom[63757] = 25'b1111111111111111000101011;
    rom[63758] = 25'b1111111111111111000101011;
    rom[63759] = 25'b1111111111111111000101011;
    rom[63760] = 25'b1111111111111111000101011;
    rom[63761] = 25'b1111111111111111000101011;
    rom[63762] = 25'b1111111111111111000101011;
    rom[63763] = 25'b1111111111111111000101010;
    rom[63764] = 25'b1111111111111111000101010;
    rom[63765] = 25'b1111111111111111000101010;
    rom[63766] = 25'b1111111111111111000101010;
    rom[63767] = 25'b1111111111111111000101010;
    rom[63768] = 25'b1111111111111111000101010;
    rom[63769] = 25'b1111111111111111000101010;
    rom[63770] = 25'b1111111111111111000101010;
    rom[63771] = 25'b1111111111111111000101010;
    rom[63772] = 25'b1111111111111111000101010;
    rom[63773] = 25'b1111111111111111000101010;
    rom[63774] = 25'b1111111111111111000101010;
    rom[63775] = 25'b1111111111111111000101010;
    rom[63776] = 25'b1111111111111111000101010;
    rom[63777] = 25'b1111111111111111000101010;
    rom[63778] = 25'b1111111111111111000101010;
    rom[63779] = 25'b1111111111111111000101001;
    rom[63780] = 25'b1111111111111111000101001;
    rom[63781] = 25'b1111111111111111000101001;
    rom[63782] = 25'b1111111111111111000101001;
    rom[63783] = 25'b1111111111111111000101001;
    rom[63784] = 25'b1111111111111111000101001;
    rom[63785] = 25'b1111111111111111000101001;
    rom[63786] = 25'b1111111111111111000101001;
    rom[63787] = 25'b1111111111111111000101001;
    rom[63788] = 25'b1111111111111111000101000;
    rom[63789] = 25'b1111111111111111000101000;
    rom[63790] = 25'b1111111111111111000101000;
    rom[63791] = 25'b1111111111111111000101000;
    rom[63792] = 25'b1111111111111111000101000;
    rom[63793] = 25'b1111111111111111000101000;
    rom[63794] = 25'b1111111111111111000101000;
    rom[63795] = 25'b1111111111111111000101000;
    rom[63796] = 25'b1111111111111111000101000;
    rom[63797] = 25'b1111111111111111000101000;
    rom[63798] = 25'b1111111111111111000100111;
    rom[63799] = 25'b1111111111111111000100111;
    rom[63800] = 25'b1111111111111111000100111;
    rom[63801] = 25'b1111111111111111000100111;
    rom[63802] = 25'b1111111111111111000100111;
    rom[63803] = 25'b1111111111111111000100111;
    rom[63804] = 25'b1111111111111111000100111;
    rom[63805] = 25'b1111111111111111000100111;
    rom[63806] = 25'b1111111111111111000100111;
    rom[63807] = 25'b1111111111111111000100111;
    rom[63808] = 25'b1111111111111111000100111;
    rom[63809] = 25'b1111111111111111000100111;
    rom[63810] = 25'b1111111111111111000100111;
    rom[63811] = 25'b1111111111111111000100111;
    rom[63812] = 25'b1111111111111111000100111;
    rom[63813] = 25'b1111111111111111000100111;
    rom[63814] = 25'b1111111111111111000100111;
    rom[63815] = 25'b1111111111111111000100111;
    rom[63816] = 25'b1111111111111111000100111;
    rom[63817] = 25'b1111111111111111000100111;
    rom[63818] = 25'b1111111111111111000100111;
    rom[63819] = 25'b1111111111111111000100111;
    rom[63820] = 25'b1111111111111111000100111;
    rom[63821] = 25'b1111111111111111000100111;
    rom[63822] = 25'b1111111111111111000100111;
    rom[63823] = 25'b1111111111111111000100111;
    rom[63824] = 25'b1111111111111111000100110;
    rom[63825] = 25'b1111111111111111000100110;
    rom[63826] = 25'b1111111111111111000100110;
    rom[63827] = 25'b1111111111111111000100110;
    rom[63828] = 25'b1111111111111111000100110;
    rom[63829] = 25'b1111111111111111000100110;
    rom[63830] = 25'b1111111111111111000100110;
    rom[63831] = 25'b1111111111111111000100110;
    rom[63832] = 25'b1111111111111111000100110;
    rom[63833] = 25'b1111111111111111000100110;
    rom[63834] = 25'b1111111111111111000100110;
    rom[63835] = 25'b1111111111111111000100110;
    rom[63836] = 25'b1111111111111111000100110;
    rom[63837] = 25'b1111111111111111000100110;
    rom[63838] = 25'b1111111111111111000100110;
    rom[63839] = 25'b1111111111111111000100110;
    rom[63840] = 25'b1111111111111111000100110;
    rom[63841] = 25'b1111111111111111000100110;
    rom[63842] = 25'b1111111111111111000100110;
    rom[63843] = 25'b1111111111111111000100110;
    rom[63844] = 25'b1111111111111111000100110;
    rom[63845] = 25'b1111111111111111000100110;
    rom[63846] = 25'b1111111111111111000100110;
    rom[63847] = 25'b1111111111111111000100101;
    rom[63848] = 25'b1111111111111111000100101;
    rom[63849] = 25'b1111111111111111000100101;
    rom[63850] = 25'b1111111111111111000100101;
    rom[63851] = 25'b1111111111111111000100101;
    rom[63852] = 25'b1111111111111111000100101;
    rom[63853] = 25'b1111111111111111000100101;
    rom[63854] = 25'b1111111111111111000100101;
    rom[63855] = 25'b1111111111111111000100101;
    rom[63856] = 25'b1111111111111111000100101;
    rom[63857] = 25'b1111111111111111000100101;
    rom[63858] = 25'b1111111111111111000100101;
    rom[63859] = 25'b1111111111111111000100101;
    rom[63860] = 25'b1111111111111111000100101;
    rom[63861] = 25'b1111111111111111000100101;
    rom[63862] = 25'b1111111111111111000100101;
    rom[63863] = 25'b1111111111111111000100101;
    rom[63864] = 25'b1111111111111111000100101;
    rom[63865] = 25'b1111111111111111000100101;
    rom[63866] = 25'b1111111111111111000100101;
    rom[63867] = 25'b1111111111111111000100101;
    rom[63868] = 25'b1111111111111111000100101;
    rom[63869] = 25'b1111111111111111000100101;
    rom[63870] = 25'b1111111111111111000100101;
    rom[63871] = 25'b1111111111111111000100101;
    rom[63872] = 25'b1111111111111111000100101;
    rom[63873] = 25'b1111111111111111000100101;
    rom[63874] = 25'b1111111111111111000100101;
    rom[63875] = 25'b1111111111111111000100101;
    rom[63876] = 25'b1111111111111111000100101;
    rom[63877] = 25'b1111111111111111000100101;
    rom[63878] = 25'b1111111111111111000100101;
    rom[63879] = 25'b1111111111111111000100101;
    rom[63880] = 25'b1111111111111111000100101;
    rom[63881] = 25'b1111111111111111000100101;
    rom[63882] = 25'b1111111111111111000100101;
    rom[63883] = 25'b1111111111111111000100101;
    rom[63884] = 25'b1111111111111111000100101;
    rom[63885] = 25'b1111111111111111000100101;
    rom[63886] = 25'b1111111111111111000100101;
    rom[63887] = 25'b1111111111111111000100101;
    rom[63888] = 25'b1111111111111111000100101;
    rom[63889] = 25'b1111111111111111000100101;
    rom[63890] = 25'b1111111111111111000100101;
    rom[63891] = 25'b1111111111111111000100101;
    rom[63892] = 25'b1111111111111111000100101;
    rom[63893] = 25'b1111111111111111000100101;
    rom[63894] = 25'b1111111111111111000100101;
    rom[63895] = 25'b1111111111111111000100101;
    rom[63896] = 25'b1111111111111111000100110;
    rom[63897] = 25'b1111111111111111000100110;
    rom[63898] = 25'b1111111111111111000100110;
    rom[63899] = 25'b1111111111111111000100110;
    rom[63900] = 25'b1111111111111111000100110;
    rom[63901] = 25'b1111111111111111000100110;
    rom[63902] = 25'b1111111111111111000100110;
    rom[63903] = 25'b1111111111111111000100110;
    rom[63904] = 25'b1111111111111111000100110;
    rom[63905] = 25'b1111111111111111000100110;
    rom[63906] = 25'b1111111111111111000100110;
    rom[63907] = 25'b1111111111111111000100110;
    rom[63908] = 25'b1111111111111111000100110;
    rom[63909] = 25'b1111111111111111000100110;
    rom[63910] = 25'b1111111111111111000100110;
    rom[63911] = 25'b1111111111111111000100110;
    rom[63912] = 25'b1111111111111111000100110;
    rom[63913] = 25'b1111111111111111000100110;
    rom[63914] = 25'b1111111111111111000100110;
    rom[63915] = 25'b1111111111111111000100110;
    rom[63916] = 25'b1111111111111111000100110;
    rom[63917] = 25'b1111111111111111000100110;
    rom[63918] = 25'b1111111111111111000100110;
    rom[63919] = 25'b1111111111111111000100111;
    rom[63920] = 25'b1111111111111111000100111;
    rom[63921] = 25'b1111111111111111000100111;
    rom[63922] = 25'b1111111111111111000100111;
    rom[63923] = 25'b1111111111111111000100111;
    rom[63924] = 25'b1111111111111111000100111;
    rom[63925] = 25'b1111111111111111000100111;
    rom[63926] = 25'b1111111111111111000100111;
    rom[63927] = 25'b1111111111111111000100111;
    rom[63928] = 25'b1111111111111111000100111;
    rom[63929] = 25'b1111111111111111000100111;
    rom[63930] = 25'b1111111111111111000100111;
    rom[63931] = 25'b1111111111111111000100111;
    rom[63932] = 25'b1111111111111111000100111;
    rom[63933] = 25'b1111111111111111000100111;
    rom[63934] = 25'b1111111111111111000100111;
    rom[63935] = 25'b1111111111111111000100111;
    rom[63936] = 25'b1111111111111111000100111;
    rom[63937] = 25'b1111111111111111000100111;
    rom[63938] = 25'b1111111111111111000100111;
    rom[63939] = 25'b1111111111111111000100111;
    rom[63940] = 25'b1111111111111111000100111;
    rom[63941] = 25'b1111111111111111000100111;
    rom[63942] = 25'b1111111111111111000100111;
    rom[63943] = 25'b1111111111111111000100111;
    rom[63944] = 25'b1111111111111111000100111;
    rom[63945] = 25'b1111111111111111000100111;
    rom[63946] = 25'b1111111111111111000100111;
    rom[63947] = 25'b1111111111111111000101000;
    rom[63948] = 25'b1111111111111111000101000;
    rom[63949] = 25'b1111111111111111000101000;
    rom[63950] = 25'b1111111111111111000101000;
    rom[63951] = 25'b1111111111111111000101000;
    rom[63952] = 25'b1111111111111111000101000;
    rom[63953] = 25'b1111111111111111000101000;
    rom[63954] = 25'b1111111111111111000101000;
    rom[63955] = 25'b1111111111111111000101000;
    rom[63956] = 25'b1111111111111111000101000;
    rom[63957] = 25'b1111111111111111000101001;
    rom[63958] = 25'b1111111111111111000101001;
    rom[63959] = 25'b1111111111111111000101001;
    rom[63960] = 25'b1111111111111111000101001;
    rom[63961] = 25'b1111111111111111000101001;
    rom[63962] = 25'b1111111111111111000101001;
    rom[63963] = 25'b1111111111111111000101001;
    rom[63964] = 25'b1111111111111111000101001;
    rom[63965] = 25'b1111111111111111000101001;
    rom[63966] = 25'b1111111111111111000101001;
    rom[63967] = 25'b1111111111111111000101010;
    rom[63968] = 25'b1111111111111111000101010;
    rom[63969] = 25'b1111111111111111000101010;
    rom[63970] = 25'b1111111111111111000101010;
    rom[63971] = 25'b1111111111111111000101010;
    rom[63972] = 25'b1111111111111111000101010;
    rom[63973] = 25'b1111111111111111000101010;
    rom[63974] = 25'b1111111111111111000101010;
    rom[63975] = 25'b1111111111111111000101010;
    rom[63976] = 25'b1111111111111111000101010;
    rom[63977] = 25'b1111111111111111000101010;
    rom[63978] = 25'b1111111111111111000101010;
    rom[63979] = 25'b1111111111111111000101010;
    rom[63980] = 25'b1111111111111111000101010;
    rom[63981] = 25'b1111111111111111000101010;
    rom[63982] = 25'b1111111111111111000101010;
    rom[63983] = 25'b1111111111111111000101010;
    rom[63984] = 25'b1111111111111111000101011;
    rom[63985] = 25'b1111111111111111000101011;
    rom[63986] = 25'b1111111111111111000101011;
    rom[63987] = 25'b1111111111111111000101011;
    rom[63988] = 25'b1111111111111111000101011;
    rom[63989] = 25'b1111111111111111000101011;
    rom[63990] = 25'b1111111111111111000101011;
    rom[63991] = 25'b1111111111111111000101100;
    rom[63992] = 25'b1111111111111111000101100;
    rom[63993] = 25'b1111111111111111000101100;
    rom[63994] = 25'b1111111111111111000101100;
    rom[63995] = 25'b1111111111111111000101100;
    rom[63996] = 25'b1111111111111111000101100;
    rom[63997] = 25'b1111111111111111000101100;
    rom[63998] = 25'b1111111111111111000101100;
    rom[63999] = 25'b1111111111111111000101101;
    rom[64000] = 25'b1111111111111111000101101;
    rom[64001] = 25'b1111111111111111000101101;
    rom[64002] = 25'b1111111111111111000101101;
    rom[64003] = 25'b1111111111111111000101101;
    rom[64004] = 25'b1111111111111111000101101;
    rom[64005] = 25'b1111111111111111000101101;
    rom[64006] = 25'b1111111111111111000101101;
    rom[64007] = 25'b1111111111111111000101101;
    rom[64008] = 25'b1111111111111111000101101;
    rom[64009] = 25'b1111111111111111000101101;
    rom[64010] = 25'b1111111111111111000101101;
    rom[64011] = 25'b1111111111111111000101101;
    rom[64012] = 25'b1111111111111111000101110;
    rom[64013] = 25'b1111111111111111000101110;
    rom[64014] = 25'b1111111111111111000101110;
    rom[64015] = 25'b1111111111111111000101110;
    rom[64016] = 25'b1111111111111111000101110;
    rom[64017] = 25'b1111111111111111000101110;
    rom[64018] = 25'b1111111111111111000101111;
    rom[64019] = 25'b1111111111111111000101111;
    rom[64020] = 25'b1111111111111111000101111;
    rom[64021] = 25'b1111111111111111000101111;
    rom[64022] = 25'b1111111111111111000101111;
    rom[64023] = 25'b1111111111111111000101111;
    rom[64024] = 25'b1111111111111111000110000;
    rom[64025] = 25'b1111111111111111000110000;
    rom[64026] = 25'b1111111111111111000110000;
    rom[64027] = 25'b1111111111111111000110000;
    rom[64028] = 25'b1111111111111111000110000;
    rom[64029] = 25'b1111111111111111000110000;
    rom[64030] = 25'b1111111111111111000110000;
    rom[64031] = 25'b1111111111111111000110000;
    rom[64032] = 25'b1111111111111111000110000;
    rom[64033] = 25'b1111111111111111000110000;
    rom[64034] = 25'b1111111111111111000110000;
    rom[64035] = 25'b1111111111111111000110000;
    rom[64036] = 25'b1111111111111111000110001;
    rom[64037] = 25'b1111111111111111000110001;
    rom[64038] = 25'b1111111111111111000110001;
    rom[64039] = 25'b1111111111111111000110001;
    rom[64040] = 25'b1111111111111111000110001;
    rom[64041] = 25'b1111111111111111000110010;
    rom[64042] = 25'b1111111111111111000110010;
    rom[64043] = 25'b1111111111111111000110010;
    rom[64044] = 25'b1111111111111111000110010;
    rom[64045] = 25'b1111111111111111000110010;
    rom[64046] = 25'b1111111111111111000110010;
    rom[64047] = 25'b1111111111111111000110011;
    rom[64048] = 25'b1111111111111111000110011;
    rom[64049] = 25'b1111111111111111000110011;
    rom[64050] = 25'b1111111111111111000110011;
    rom[64051] = 25'b1111111111111111000110011;
    rom[64052] = 25'b1111111111111111000110011;
    rom[64053] = 25'b1111111111111111000110011;
    rom[64054] = 25'b1111111111111111000110011;
    rom[64055] = 25'b1111111111111111000110011;
    rom[64056] = 25'b1111111111111111000110011;
    rom[64057] = 25'b1111111111111111000110100;
    rom[64058] = 25'b1111111111111111000110100;
    rom[64059] = 25'b1111111111111111000110100;
    rom[64060] = 25'b1111111111111111000110100;
    rom[64061] = 25'b1111111111111111000110100;
    rom[64062] = 25'b1111111111111111000110101;
    rom[64063] = 25'b1111111111111111000110101;
    rom[64064] = 25'b1111111111111111000110101;
    rom[64065] = 25'b1111111111111111000110101;
    rom[64066] = 25'b1111111111111111000110101;
    rom[64067] = 25'b1111111111111111000110110;
    rom[64068] = 25'b1111111111111111000110110;
    rom[64069] = 25'b1111111111111111000110110;
    rom[64070] = 25'b1111111111111111000110110;
    rom[64071] = 25'b1111111111111111000110110;
    rom[64072] = 25'b1111111111111111000110110;
    rom[64073] = 25'b1111111111111111000110110;
    rom[64074] = 25'b1111111111111111000110110;
    rom[64075] = 25'b1111111111111111000110110;
    rom[64076] = 25'b1111111111111111000110111;
    rom[64077] = 25'b1111111111111111000110111;
    rom[64078] = 25'b1111111111111111000110111;
    rom[64079] = 25'b1111111111111111000110111;
    rom[64080] = 25'b1111111111111111000111000;
    rom[64081] = 25'b1111111111111111000111000;
    rom[64082] = 25'b1111111111111111000111000;
    rom[64083] = 25'b1111111111111111000111000;
    rom[64084] = 25'b1111111111111111000111000;
    rom[64085] = 25'b1111111111111111000111001;
    rom[64086] = 25'b1111111111111111000111001;
    rom[64087] = 25'b1111111111111111000111001;
    rom[64088] = 25'b1111111111111111000111001;
    rom[64089] = 25'b1111111111111111000111001;
    rom[64090] = 25'b1111111111111111000111001;
    rom[64091] = 25'b1111111111111111000111001;
    rom[64092] = 25'b1111111111111111000111001;
    rom[64093] = 25'b1111111111111111000111001;
    rom[64094] = 25'b1111111111111111000111010;
    rom[64095] = 25'b1111111111111111000111010;
    rom[64096] = 25'b1111111111111111000111010;
    rom[64097] = 25'b1111111111111111000111010;
    rom[64098] = 25'b1111111111111111000111011;
    rom[64099] = 25'b1111111111111111000111011;
    rom[64100] = 25'b1111111111111111000111011;
    rom[64101] = 25'b1111111111111111000111011;
    rom[64102] = 25'b1111111111111111000111100;
    rom[64103] = 25'b1111111111111111000111100;
    rom[64104] = 25'b1111111111111111000111100;
    rom[64105] = 25'b1111111111111111000111100;
    rom[64106] = 25'b1111111111111111000111100;
    rom[64107] = 25'b1111111111111111000111100;
    rom[64108] = 25'b1111111111111111000111100;
    rom[64109] = 25'b1111111111111111000111100;
    rom[64110] = 25'b1111111111111111000111101;
    rom[64111] = 25'b1111111111111111000111101;
    rom[64112] = 25'b1111111111111111000111101;
    rom[64113] = 25'b1111111111111111000111101;
    rom[64114] = 25'b1111111111111111000111110;
    rom[64115] = 25'b1111111111111111000111110;
    rom[64116] = 25'b1111111111111111000111110;
    rom[64117] = 25'b1111111111111111000111110;
    rom[64118] = 25'b1111111111111111000111110;
    rom[64119] = 25'b1111111111111111000111110;
    rom[64120] = 25'b1111111111111111000111110;
    rom[64121] = 25'b1111111111111111000111110;
    rom[64122] = 25'b1111111111111111000111111;
    rom[64123] = 25'b1111111111111111000111111;
    rom[64124] = 25'b1111111111111111000111111;
    rom[64125] = 25'b1111111111111111000111111;
    rom[64126] = 25'b1111111111111111001000000;
    rom[64127] = 25'b1111111111111111001000000;
    rom[64128] = 25'b1111111111111111001000000;
    rom[64129] = 25'b1111111111111111001000000;
    rom[64130] = 25'b1111111111111111001000001;
    rom[64131] = 25'b1111111111111111001000001;
    rom[64132] = 25'b1111111111111111001000001;
    rom[64133] = 25'b1111111111111111001000001;
    rom[64134] = 25'b1111111111111111001000001;
    rom[64135] = 25'b1111111111111111001000001;
    rom[64136] = 25'b1111111111111111001000001;
    rom[64137] = 25'b1111111111111111001000010;
    rom[64138] = 25'b1111111111111111001000010;
    rom[64139] = 25'b1111111111111111001000010;
    rom[64140] = 25'b1111111111111111001000010;
    rom[64141] = 25'b1111111111111111001000011;
    rom[64142] = 25'b1111111111111111001000011;
    rom[64143] = 25'b1111111111111111001000011;
    rom[64144] = 25'b1111111111111111001000011;
    rom[64145] = 25'b1111111111111111001000100;
    rom[64146] = 25'b1111111111111111001000100;
    rom[64147] = 25'b1111111111111111001000100;
    rom[64148] = 25'b1111111111111111001000100;
    rom[64149] = 25'b1111111111111111001000100;
    rom[64150] = 25'b1111111111111111001000100;
    rom[64151] = 25'b1111111111111111001000100;
    rom[64152] = 25'b1111111111111111001000101;
    rom[64153] = 25'b1111111111111111001000101;
    rom[64154] = 25'b1111111111111111001000101;
    rom[64155] = 25'b1111111111111111001000110;
    rom[64156] = 25'b1111111111111111001000110;
    rom[64157] = 25'b1111111111111111001000110;
    rom[64158] = 25'b1111111111111111001000110;
    rom[64159] = 25'b1111111111111111001000111;
    rom[64160] = 25'b1111111111111111001000111;
    rom[64161] = 25'b1111111111111111001000111;
    rom[64162] = 25'b1111111111111111001000111;
    rom[64163] = 25'b1111111111111111001000111;
    rom[64164] = 25'b1111111111111111001000111;
    rom[64165] = 25'b1111111111111111001000111;
    rom[64166] = 25'b1111111111111111001001000;
    rom[64167] = 25'b1111111111111111001001000;
    rom[64168] = 25'b1111111111111111001001000;
    rom[64169] = 25'b1111111111111111001001001;
    rom[64170] = 25'b1111111111111111001001001;
    rom[64171] = 25'b1111111111111111001001001;
    rom[64172] = 25'b1111111111111111001001010;
    rom[64173] = 25'b1111111111111111001001010;
    rom[64174] = 25'b1111111111111111001001010;
    rom[64175] = 25'b1111111111111111001001010;
    rom[64176] = 25'b1111111111111111001001010;
    rom[64177] = 25'b1111111111111111001001010;
    rom[64178] = 25'b1111111111111111001001010;
    rom[64179] = 25'b1111111111111111001001011;
    rom[64180] = 25'b1111111111111111001001011;
    rom[64181] = 25'b1111111111111111001001011;
    rom[64182] = 25'b1111111111111111001001100;
    rom[64183] = 25'b1111111111111111001001100;
    rom[64184] = 25'b1111111111111111001001100;
    rom[64185] = 25'b1111111111111111001001100;
    rom[64186] = 25'b1111111111111111001001101;
    rom[64187] = 25'b1111111111111111001001101;
    rom[64188] = 25'b1111111111111111001001101;
    rom[64189] = 25'b1111111111111111001001101;
    rom[64190] = 25'b1111111111111111001001101;
    rom[64191] = 25'b1111111111111111001001101;
    rom[64192] = 25'b1111111111111111001001110;
    rom[64193] = 25'b1111111111111111001001110;
    rom[64194] = 25'b1111111111111111001001110;
    rom[64195] = 25'b1111111111111111001001111;
    rom[64196] = 25'b1111111111111111001001111;
    rom[64197] = 25'b1111111111111111001001111;
    rom[64198] = 25'b1111111111111111001010000;
    rom[64199] = 25'b1111111111111111001010000;
    rom[64200] = 25'b1111111111111111001010000;
    rom[64201] = 25'b1111111111111111001010000;
    rom[64202] = 25'b1111111111111111001010000;
    rom[64203] = 25'b1111111111111111001010000;
    rom[64204] = 25'b1111111111111111001010000;
    rom[64205] = 25'b1111111111111111001010001;
    rom[64206] = 25'b1111111111111111001010001;
    rom[64207] = 25'b1111111111111111001010001;
    rom[64208] = 25'b1111111111111111001010010;
    rom[64209] = 25'b1111111111111111001010010;
    rom[64210] = 25'b1111111111111111001010010;
    rom[64211] = 25'b1111111111111111001010011;
    rom[64212] = 25'b1111111111111111001010011;
    rom[64213] = 25'b1111111111111111001010011;
    rom[64214] = 25'b1111111111111111001010011;
    rom[64215] = 25'b1111111111111111001010011;
    rom[64216] = 25'b1111111111111111001010011;
    rom[64217] = 25'b1111111111111111001010100;
    rom[64218] = 25'b1111111111111111001010100;
    rom[64219] = 25'b1111111111111111001010100;
    rom[64220] = 25'b1111111111111111001010101;
    rom[64221] = 25'b1111111111111111001010101;
    rom[64222] = 25'b1111111111111111001010101;
    rom[64223] = 25'b1111111111111111001010110;
    rom[64224] = 25'b1111111111111111001010110;
    rom[64225] = 25'b1111111111111111001010110;
    rom[64226] = 25'b1111111111111111001010110;
    rom[64227] = 25'b1111111111111111001010110;
    rom[64228] = 25'b1111111111111111001010110;
    rom[64229] = 25'b1111111111111111001010111;
    rom[64230] = 25'b1111111111111111001010111;
    rom[64231] = 25'b1111111111111111001010111;
    rom[64232] = 25'b1111111111111111001011000;
    rom[64233] = 25'b1111111111111111001011000;
    rom[64234] = 25'b1111111111111111001011000;
    rom[64235] = 25'b1111111111111111001011001;
    rom[64236] = 25'b1111111111111111001011001;
    rom[64237] = 25'b1111111111111111001011001;
    rom[64238] = 25'b1111111111111111001011001;
    rom[64239] = 25'b1111111111111111001011001;
    rom[64240] = 25'b1111111111111111001011001;
    rom[64241] = 25'b1111111111111111001011010;
    rom[64242] = 25'b1111111111111111001011010;
    rom[64243] = 25'b1111111111111111001011010;
    rom[64244] = 25'b1111111111111111001011011;
    rom[64245] = 25'b1111111111111111001011011;
    rom[64246] = 25'b1111111111111111001011011;
    rom[64247] = 25'b1111111111111111001011100;
    rom[64248] = 25'b1111111111111111001011100;
    rom[64249] = 25'b1111111111111111001011100;
    rom[64250] = 25'b1111111111111111001011100;
    rom[64251] = 25'b1111111111111111001011100;
    rom[64252] = 25'b1111111111111111001011101;
    rom[64253] = 25'b1111111111111111001011101;
    rom[64254] = 25'b1111111111111111001011101;
    rom[64255] = 25'b1111111111111111001011110;
    rom[64256] = 25'b1111111111111111001011110;
    rom[64257] = 25'b1111111111111111001011110;
    rom[64258] = 25'b1111111111111111001011111;
    rom[64259] = 25'b1111111111111111001011111;
    rom[64260] = 25'b1111111111111111001011111;
    rom[64261] = 25'b1111111111111111001011111;
    rom[64262] = 25'b1111111111111111001011111;
    rom[64263] = 25'b1111111111111111001100000;
    rom[64264] = 25'b1111111111111111001100000;
    rom[64265] = 25'b1111111111111111001100000;
    rom[64266] = 25'b1111111111111111001100001;
    rom[64267] = 25'b1111111111111111001100001;
    rom[64268] = 25'b1111111111111111001100001;
    rom[64269] = 25'b1111111111111111001100010;
    rom[64270] = 25'b1111111111111111001100010;
    rom[64271] = 25'b1111111111111111001100010;
    rom[64272] = 25'b1111111111111111001100010;
    rom[64273] = 25'b1111111111111111001100010;
    rom[64274] = 25'b1111111111111111001100010;
    rom[64275] = 25'b1111111111111111001100011;
    rom[64276] = 25'b1111111111111111001100011;
    rom[64277] = 25'b1111111111111111001100100;
    rom[64278] = 25'b1111111111111111001100100;
    rom[64279] = 25'b1111111111111111001100100;
    rom[64280] = 25'b1111111111111111001100101;
    rom[64281] = 25'b1111111111111111001100101;
    rom[64282] = 25'b1111111111111111001100101;
    rom[64283] = 25'b1111111111111111001100101;
    rom[64284] = 25'b1111111111111111001100101;
    rom[64285] = 25'b1111111111111111001100110;
    rom[64286] = 25'b1111111111111111001100110;
    rom[64287] = 25'b1111111111111111001100110;
    rom[64288] = 25'b1111111111111111001100111;
    rom[64289] = 25'b1111111111111111001100111;
    rom[64290] = 25'b1111111111111111001100111;
    rom[64291] = 25'b1111111111111111001101000;
    rom[64292] = 25'b1111111111111111001101000;
    rom[64293] = 25'b1111111111111111001101000;
    rom[64294] = 25'b1111111111111111001101000;
    rom[64295] = 25'b1111111111111111001101000;
    rom[64296] = 25'b1111111111111111001101001;
    rom[64297] = 25'b1111111111111111001101001;
    rom[64298] = 25'b1111111111111111001101001;
    rom[64299] = 25'b1111111111111111001101010;
    rom[64300] = 25'b1111111111111111001101010;
    rom[64301] = 25'b1111111111111111001101011;
    rom[64302] = 25'b1111111111111111001101011;
    rom[64303] = 25'b1111111111111111001101011;
    rom[64304] = 25'b1111111111111111001101011;
    rom[64305] = 25'b1111111111111111001101011;
    rom[64306] = 25'b1111111111111111001101011;
    rom[64307] = 25'b1111111111111111001101100;
    rom[64308] = 25'b1111111111111111001101100;
    rom[64309] = 25'b1111111111111111001101101;
    rom[64310] = 25'b1111111111111111001101101;
    rom[64311] = 25'b1111111111111111001101101;
    rom[64312] = 25'b1111111111111111001101110;
    rom[64313] = 25'b1111111111111111001101110;
    rom[64314] = 25'b1111111111111111001101110;
    rom[64315] = 25'b1111111111111111001101110;
    rom[64316] = 25'b1111111111111111001101110;
    rom[64317] = 25'b1111111111111111001101111;
    rom[64318] = 25'b1111111111111111001101111;
    rom[64319] = 25'b1111111111111111001101111;
    rom[64320] = 25'b1111111111111111001110000;
    rom[64321] = 25'b1111111111111111001110000;
    rom[64322] = 25'b1111111111111111001110001;
    rom[64323] = 25'b1111111111111111001110001;
    rom[64324] = 25'b1111111111111111001110001;
    rom[64325] = 25'b1111111111111111001110001;
    rom[64326] = 25'b1111111111111111001110001;
    rom[64327] = 25'b1111111111111111001110010;
    rom[64328] = 25'b1111111111111111001110010;
    rom[64329] = 25'b1111111111111111001110010;
    rom[64330] = 25'b1111111111111111001110011;
    rom[64331] = 25'b1111111111111111001110011;
    rom[64332] = 25'b1111111111111111001110100;
    rom[64333] = 25'b1111111111111111001110100;
    rom[64334] = 25'b1111111111111111001110100;
    rom[64335] = 25'b1111111111111111001110100;
    rom[64336] = 25'b1111111111111111001110100;
    rom[64337] = 25'b1111111111111111001110101;
    rom[64338] = 25'b1111111111111111001110101;
    rom[64339] = 25'b1111111111111111001110101;
    rom[64340] = 25'b1111111111111111001110110;
    rom[64341] = 25'b1111111111111111001110110;
    rom[64342] = 25'b1111111111111111001110111;
    rom[64343] = 25'b1111111111111111001110111;
    rom[64344] = 25'b1111111111111111001110111;
    rom[64345] = 25'b1111111111111111001110111;
    rom[64346] = 25'b1111111111111111001110111;
    rom[64347] = 25'b1111111111111111001111000;
    rom[64348] = 25'b1111111111111111001111000;
    rom[64349] = 25'b1111111111111111001111000;
    rom[64350] = 25'b1111111111111111001111001;
    rom[64351] = 25'b1111111111111111001111001;
    rom[64352] = 25'b1111111111111111001111010;
    rom[64353] = 25'b1111111111111111001111010;
    rom[64354] = 25'b1111111111111111001111010;
    rom[64355] = 25'b1111111111111111001111010;
    rom[64356] = 25'b1111111111111111001111010;
    rom[64357] = 25'b1111111111111111001111011;
    rom[64358] = 25'b1111111111111111001111011;
    rom[64359] = 25'b1111111111111111001111011;
    rom[64360] = 25'b1111111111111111001111100;
    rom[64361] = 25'b1111111111111111001111100;
    rom[64362] = 25'b1111111111111111001111101;
    rom[64363] = 25'b1111111111111111001111101;
    rom[64364] = 25'b1111111111111111001111101;
    rom[64365] = 25'b1111111111111111001111101;
    rom[64366] = 25'b1111111111111111001111101;
    rom[64367] = 25'b1111111111111111001111110;
    rom[64368] = 25'b1111111111111111001111110;
    rom[64369] = 25'b1111111111111111001111111;
    rom[64370] = 25'b1111111111111111001111111;
    rom[64371] = 25'b1111111111111111001111111;
    rom[64372] = 25'b1111111111111111001111111;
    rom[64373] = 25'b1111111111111111001111111;
    rom[64374] = 25'b1111111111111111010000000;
    rom[64375] = 25'b1111111111111111010000000;
    rom[64376] = 25'b1111111111111111010000000;
    rom[64377] = 25'b1111111111111111010000001;
    rom[64378] = 25'b1111111111111111010000001;
    rom[64379] = 25'b1111111111111111010000010;
    rom[64380] = 25'b1111111111111111010000010;
    rom[64381] = 25'b1111111111111111010000010;
    rom[64382] = 25'b1111111111111111010000010;
    rom[64383] = 25'b1111111111111111010000010;
    rom[64384] = 25'b1111111111111111010000011;
    rom[64385] = 25'b1111111111111111010000011;
    rom[64386] = 25'b1111111111111111010000100;
    rom[64387] = 25'b1111111111111111010000100;
    rom[64388] = 25'b1111111111111111010000100;
    rom[64389] = 25'b1111111111111111010000101;
    rom[64390] = 25'b1111111111111111010000101;
    rom[64391] = 25'b1111111111111111010000101;
    rom[64392] = 25'b1111111111111111010000101;
    rom[64393] = 25'b1111111111111111010000110;
    rom[64394] = 25'b1111111111111111010000110;
    rom[64395] = 25'b1111111111111111010000110;
    rom[64396] = 25'b1111111111111111010000111;
    rom[64397] = 25'b1111111111111111010000111;
    rom[64398] = 25'b1111111111111111010001000;
    rom[64399] = 25'b1111111111111111010001000;
    rom[64400] = 25'b1111111111111111010001000;
    rom[64401] = 25'b1111111111111111010001000;
    rom[64402] = 25'b1111111111111111010001000;
    rom[64403] = 25'b1111111111111111010001001;
    rom[64404] = 25'b1111111111111111010001001;
    rom[64405] = 25'b1111111111111111010001010;
    rom[64406] = 25'b1111111111111111010001010;
    rom[64407] = 25'b1111111111111111010001011;
    rom[64408] = 25'b1111111111111111010001011;
    rom[64409] = 25'b1111111111111111010001011;
    rom[64410] = 25'b1111111111111111010001011;
    rom[64411] = 25'b1111111111111111010001011;
    rom[64412] = 25'b1111111111111111010001100;
    rom[64413] = 25'b1111111111111111010001100;
    rom[64414] = 25'b1111111111111111010001101;
    rom[64415] = 25'b1111111111111111010001101;
    rom[64416] = 25'b1111111111111111010001101;
    rom[64417] = 25'b1111111111111111010001110;
    rom[64418] = 25'b1111111111111111010001110;
    rom[64419] = 25'b1111111111111111010001110;
    rom[64420] = 25'b1111111111111111010001110;
    rom[64421] = 25'b1111111111111111010001111;
    rom[64422] = 25'b1111111111111111010001111;
    rom[64423] = 25'b1111111111111111010001111;
    rom[64424] = 25'b1111111111111111010010000;
    rom[64425] = 25'b1111111111111111010010000;
    rom[64426] = 25'b1111111111111111010010001;
    rom[64427] = 25'b1111111111111111010010001;
    rom[64428] = 25'b1111111111111111010010001;
    rom[64429] = 25'b1111111111111111010010001;
    rom[64430] = 25'b1111111111111111010010001;
    rom[64431] = 25'b1111111111111111010010010;
    rom[64432] = 25'b1111111111111111010010010;
    rom[64433] = 25'b1111111111111111010010011;
    rom[64434] = 25'b1111111111111111010010011;
    rom[64435] = 25'b1111111111111111010010100;
    rom[64436] = 25'b1111111111111111010010100;
    rom[64437] = 25'b1111111111111111010010100;
    rom[64438] = 25'b1111111111111111010010100;
    rom[64439] = 25'b1111111111111111010010100;
    rom[64440] = 25'b1111111111111111010010101;
    rom[64441] = 25'b1111111111111111010010101;
    rom[64442] = 25'b1111111111111111010010110;
    rom[64443] = 25'b1111111111111111010010110;
    rom[64444] = 25'b1111111111111111010010111;
    rom[64445] = 25'b1111111111111111010010111;
    rom[64446] = 25'b1111111111111111010010111;
    rom[64447] = 25'b1111111111111111010010111;
    rom[64448] = 25'b1111111111111111010010111;
    rom[64449] = 25'b1111111111111111010011000;
    rom[64450] = 25'b1111111111111111010011000;
    rom[64451] = 25'b1111111111111111010011001;
    rom[64452] = 25'b1111111111111111010011001;
    rom[64453] = 25'b1111111111111111010011010;
    rom[64454] = 25'b1111111111111111010011010;
    rom[64455] = 25'b1111111111111111010011010;
    rom[64456] = 25'b1111111111111111010011010;
    rom[64457] = 25'b1111111111111111010011010;
    rom[64458] = 25'b1111111111111111010011011;
    rom[64459] = 25'b1111111111111111010011011;
    rom[64460] = 25'b1111111111111111010011100;
    rom[64461] = 25'b1111111111111111010011100;
    rom[64462] = 25'b1111111111111111010011101;
    rom[64463] = 25'b1111111111111111010011101;
    rom[64464] = 25'b1111111111111111010011101;
    rom[64465] = 25'b1111111111111111010011101;
    rom[64466] = 25'b1111111111111111010011101;
    rom[64467] = 25'b1111111111111111010011110;
    rom[64468] = 25'b1111111111111111010011110;
    rom[64469] = 25'b1111111111111111010011111;
    rom[64470] = 25'b1111111111111111010011111;
    rom[64471] = 25'b1111111111111111010100000;
    rom[64472] = 25'b1111111111111111010100000;
    rom[64473] = 25'b1111111111111111010100000;
    rom[64474] = 25'b1111111111111111010100000;
    rom[64475] = 25'b1111111111111111010100000;
    rom[64476] = 25'b1111111111111111010100001;
    rom[64477] = 25'b1111111111111111010100001;
    rom[64478] = 25'b1111111111111111010100010;
    rom[64479] = 25'b1111111111111111010100010;
    rom[64480] = 25'b1111111111111111010100011;
    rom[64481] = 25'b1111111111111111010100011;
    rom[64482] = 25'b1111111111111111010100011;
    rom[64483] = 25'b1111111111111111010100011;
    rom[64484] = 25'b1111111111111111010100011;
    rom[64485] = 25'b1111111111111111010100100;
    rom[64486] = 25'b1111111111111111010100100;
    rom[64487] = 25'b1111111111111111010100101;
    rom[64488] = 25'b1111111111111111010100101;
    rom[64489] = 25'b1111111111111111010100110;
    rom[64490] = 25'b1111111111111111010100110;
    rom[64491] = 25'b1111111111111111010100110;
    rom[64492] = 25'b1111111111111111010100110;
    rom[64493] = 25'b1111111111111111010100110;
    rom[64494] = 25'b1111111111111111010100111;
    rom[64495] = 25'b1111111111111111010100111;
    rom[64496] = 25'b1111111111111111010101000;
    rom[64497] = 25'b1111111111111111010101000;
    rom[64498] = 25'b1111111111111111010101001;
    rom[64499] = 25'b1111111111111111010101001;
    rom[64500] = 25'b1111111111111111010101001;
    rom[64501] = 25'b1111111111111111010101001;
    rom[64502] = 25'b1111111111111111010101010;
    rom[64503] = 25'b1111111111111111010101010;
    rom[64504] = 25'b1111111111111111010101010;
    rom[64505] = 25'b1111111111111111010101011;
    rom[64506] = 25'b1111111111111111010101011;
    rom[64507] = 25'b1111111111111111010101100;
    rom[64508] = 25'b1111111111111111010101100;
    rom[64509] = 25'b1111111111111111010101100;
    rom[64510] = 25'b1111111111111111010101100;
    rom[64511] = 25'b1111111111111111010101101;
    rom[64512] = 25'b1111111111111111010101101;
    rom[64513] = 25'b1111111111111111010101110;
    rom[64514] = 25'b1111111111111111010101110;
    rom[64515] = 25'b1111111111111111010101110;
    rom[64516] = 25'b1111111111111111010101111;
    rom[64517] = 25'b1111111111111111010101111;
    rom[64518] = 25'b1111111111111111010101111;
    rom[64519] = 25'b1111111111111111010101111;
    rom[64520] = 25'b1111111111111111010110000;
    rom[64521] = 25'b1111111111111111010110000;
    rom[64522] = 25'b1111111111111111010110001;
    rom[64523] = 25'b1111111111111111010110001;
    rom[64524] = 25'b1111111111111111010110010;
    rom[64525] = 25'b1111111111111111010110010;
    rom[64526] = 25'b1111111111111111010110010;
    rom[64527] = 25'b1111111111111111010110010;
    rom[64528] = 25'b1111111111111111010110010;
    rom[64529] = 25'b1111111111111111010110011;
    rom[64530] = 25'b1111111111111111010110011;
    rom[64531] = 25'b1111111111111111010110100;
    rom[64532] = 25'b1111111111111111010110100;
    rom[64533] = 25'b1111111111111111010110101;
    rom[64534] = 25'b1111111111111111010110101;
    rom[64535] = 25'b1111111111111111010110101;
    rom[64536] = 25'b1111111111111111010110101;
    rom[64537] = 25'b1111111111111111010110110;
    rom[64538] = 25'b1111111111111111010110110;
    rom[64539] = 25'b1111111111111111010110110;
    rom[64540] = 25'b1111111111111111010110111;
    rom[64541] = 25'b1111111111111111010110111;
    rom[64542] = 25'b1111111111111111010111000;
    rom[64543] = 25'b1111111111111111010111000;
    rom[64544] = 25'b1111111111111111010111000;
    rom[64545] = 25'b1111111111111111010111000;
    rom[64546] = 25'b1111111111111111010111001;
    rom[64547] = 25'b1111111111111111010111001;
    rom[64548] = 25'b1111111111111111010111010;
    rom[64549] = 25'b1111111111111111010111010;
    rom[64550] = 25'b1111111111111111010111010;
    rom[64551] = 25'b1111111111111111010111011;
    rom[64552] = 25'b1111111111111111010111011;
    rom[64553] = 25'b1111111111111111010111011;
    rom[64554] = 25'b1111111111111111010111011;
    rom[64555] = 25'b1111111111111111010111100;
    rom[64556] = 25'b1111111111111111010111100;
    rom[64557] = 25'b1111111111111111010111101;
    rom[64558] = 25'b1111111111111111010111101;
    rom[64559] = 25'b1111111111111111010111110;
    rom[64560] = 25'b1111111111111111010111110;
    rom[64561] = 25'b1111111111111111010111110;
    rom[64562] = 25'b1111111111111111010111110;
    rom[64563] = 25'b1111111111111111010111111;
    rom[64564] = 25'b1111111111111111010111111;
    rom[64565] = 25'b1111111111111111010111111;
    rom[64566] = 25'b1111111111111111011000000;
    rom[64567] = 25'b1111111111111111011000000;
    rom[64568] = 25'b1111111111111111011000000;
    rom[64569] = 25'b1111111111111111011000000;
    rom[64570] = 25'b1111111111111111011000001;
    rom[64571] = 25'b1111111111111111011000001;
    rom[64572] = 25'b1111111111111111011000010;
    rom[64573] = 25'b1111111111111111011000010;
    rom[64574] = 25'b1111111111111111011000011;
    rom[64575] = 25'b1111111111111111011000011;
    rom[64576] = 25'b1111111111111111011000011;
    rom[64577] = 25'b1111111111111111011000011;
    rom[64578] = 25'b1111111111111111011000011;
    rom[64579] = 25'b1111111111111111011000100;
    rom[64580] = 25'b1111111111111111011000100;
    rom[64581] = 25'b1111111111111111011000101;
    rom[64582] = 25'b1111111111111111011000101;
    rom[64583] = 25'b1111111111111111011000110;
    rom[64584] = 25'b1111111111111111011000110;
    rom[64585] = 25'b1111111111111111011000110;
    rom[64586] = 25'b1111111111111111011000110;
    rom[64587] = 25'b1111111111111111011000111;
    rom[64588] = 25'b1111111111111111011000111;
    rom[64589] = 25'b1111111111111111011001000;
    rom[64590] = 25'b1111111111111111011001000;
    rom[64591] = 25'b1111111111111111011001000;
    rom[64592] = 25'b1111111111111111011001001;
    rom[64593] = 25'b1111111111111111011001001;
    rom[64594] = 25'b1111111111111111011001001;
    rom[64595] = 25'b1111111111111111011001001;
    rom[64596] = 25'b1111111111111111011001010;
    rom[64597] = 25'b1111111111111111011001010;
    rom[64598] = 25'b1111111111111111011001011;
    rom[64599] = 25'b1111111111111111011001011;
    rom[64600] = 25'b1111111111111111011001100;
    rom[64601] = 25'b1111111111111111011001100;
    rom[64602] = 25'b1111111111111111011001100;
    rom[64603] = 25'b1111111111111111011001100;
    rom[64604] = 25'b1111111111111111011001101;
    rom[64605] = 25'b1111111111111111011001101;
    rom[64606] = 25'b1111111111111111011001101;
    rom[64607] = 25'b1111111111111111011001110;
    rom[64608] = 25'b1111111111111111011001110;
    rom[64609] = 25'b1111111111111111011001111;
    rom[64610] = 25'b1111111111111111011001111;
    rom[64611] = 25'b1111111111111111011001111;
    rom[64612] = 25'b1111111111111111011001111;
    rom[64613] = 25'b1111111111111111011010000;
    rom[64614] = 25'b1111111111111111011010000;
    rom[64615] = 25'b1111111111111111011010001;
    rom[64616] = 25'b1111111111111111011010001;
    rom[64617] = 25'b1111111111111111011010010;
    rom[64618] = 25'b1111111111111111011010010;
    rom[64619] = 25'b1111111111111111011010010;
    rom[64620] = 25'b1111111111111111011010010;
    rom[64621] = 25'b1111111111111111011010010;
    rom[64622] = 25'b1111111111111111011010011;
    rom[64623] = 25'b1111111111111111011010011;
    rom[64624] = 25'b1111111111111111011010100;
    rom[64625] = 25'b1111111111111111011010100;
    rom[64626] = 25'b1111111111111111011010101;
    rom[64627] = 25'b1111111111111111011010101;
    rom[64628] = 25'b1111111111111111011010101;
    rom[64629] = 25'b1111111111111111011010101;
    rom[64630] = 25'b1111111111111111011010110;
    rom[64631] = 25'b1111111111111111011010110;
    rom[64632] = 25'b1111111111111111011010111;
    rom[64633] = 25'b1111111111111111011010111;
    rom[64634] = 25'b1111111111111111011011000;
    rom[64635] = 25'b1111111111111111011011000;
    rom[64636] = 25'b1111111111111111011011000;
    rom[64637] = 25'b1111111111111111011011000;
    rom[64638] = 25'b1111111111111111011011000;
    rom[64639] = 25'b1111111111111111011011001;
    rom[64640] = 25'b1111111111111111011011001;
    rom[64641] = 25'b1111111111111111011011010;
    rom[64642] = 25'b1111111111111111011011010;
    rom[64643] = 25'b1111111111111111011011011;
    rom[64644] = 25'b1111111111111111011011011;
    rom[64645] = 25'b1111111111111111011011011;
    rom[64646] = 25'b1111111111111111011011011;
    rom[64647] = 25'b1111111111111111011011100;
    rom[64648] = 25'b1111111111111111011011100;
    rom[64649] = 25'b1111111111111111011011101;
    rom[64650] = 25'b1111111111111111011011101;
    rom[64651] = 25'b1111111111111111011011101;
    rom[64652] = 25'b1111111111111111011011110;
    rom[64653] = 25'b1111111111111111011011110;
    rom[64654] = 25'b1111111111111111011011110;
    rom[64655] = 25'b1111111111111111011011110;
    rom[64656] = 25'b1111111111111111011011111;
    rom[64657] = 25'b1111111111111111011011111;
    rom[64658] = 25'b1111111111111111011100000;
    rom[64659] = 25'b1111111111111111011100000;
    rom[64660] = 25'b1111111111111111011100001;
    rom[64661] = 25'b1111111111111111011100001;
    rom[64662] = 25'b1111111111111111011100001;
    rom[64663] = 25'b1111111111111111011100001;
    rom[64664] = 25'b1111111111111111011100001;
    rom[64665] = 25'b1111111111111111011100010;
    rom[64666] = 25'b1111111111111111011100010;
    rom[64667] = 25'b1111111111111111011100011;
    rom[64668] = 25'b1111111111111111011100011;
    rom[64669] = 25'b1111111111111111011100100;
    rom[64670] = 25'b1111111111111111011100100;
    rom[64671] = 25'b1111111111111111011100100;
    rom[64672] = 25'b1111111111111111011100100;
    rom[64673] = 25'b1111111111111111011100101;
    rom[64674] = 25'b1111111111111111011100101;
    rom[64675] = 25'b1111111111111111011100110;
    rom[64676] = 25'b1111111111111111011100110;
    rom[64677] = 25'b1111111111111111011100111;
    rom[64678] = 25'b1111111111111111011100111;
    rom[64679] = 25'b1111111111111111011100111;
    rom[64680] = 25'b1111111111111111011100111;
    rom[64681] = 25'b1111111111111111011100111;
    rom[64682] = 25'b1111111111111111011101000;
    rom[64683] = 25'b1111111111111111011101000;
    rom[64684] = 25'b1111111111111111011101001;
    rom[64685] = 25'b1111111111111111011101001;
    rom[64686] = 25'b1111111111111111011101010;
    rom[64687] = 25'b1111111111111111011101010;
    rom[64688] = 25'b1111111111111111011101010;
    rom[64689] = 25'b1111111111111111011101010;
    rom[64690] = 25'b1111111111111111011101011;
    rom[64691] = 25'b1111111111111111011101011;
    rom[64692] = 25'b1111111111111111011101011;
    rom[64693] = 25'b1111111111111111011101100;
    rom[64694] = 25'b1111111111111111011101100;
    rom[64695] = 25'b1111111111111111011101101;
    rom[64696] = 25'b1111111111111111011101101;
    rom[64697] = 25'b1111111111111111011101101;
    rom[64698] = 25'b1111111111111111011101101;
    rom[64699] = 25'b1111111111111111011101110;
    rom[64700] = 25'b1111111111111111011101110;
    rom[64701] = 25'b1111111111111111011101111;
    rom[64702] = 25'b1111111111111111011101111;
    rom[64703] = 25'b1111111111111111011110000;
    rom[64704] = 25'b1111111111111111011110000;
    rom[64705] = 25'b1111111111111111011110000;
    rom[64706] = 25'b1111111111111111011110000;
    rom[64707] = 25'b1111111111111111011110000;
    rom[64708] = 25'b1111111111111111011110001;
    rom[64709] = 25'b1111111111111111011110001;
    rom[64710] = 25'b1111111111111111011110010;
    rom[64711] = 25'b1111111111111111011110010;
    rom[64712] = 25'b1111111111111111011110011;
    rom[64713] = 25'b1111111111111111011110011;
    rom[64714] = 25'b1111111111111111011110011;
    rom[64715] = 25'b1111111111111111011110011;
    rom[64716] = 25'b1111111111111111011110100;
    rom[64717] = 25'b1111111111111111011110100;
    rom[64718] = 25'b1111111111111111011110100;
    rom[64719] = 25'b1111111111111111011110101;
    rom[64720] = 25'b1111111111111111011110101;
    rom[64721] = 25'b1111111111111111011110110;
    rom[64722] = 25'b1111111111111111011110110;
    rom[64723] = 25'b1111111111111111011110110;
    rom[64724] = 25'b1111111111111111011110110;
    rom[64725] = 25'b1111111111111111011110111;
    rom[64726] = 25'b1111111111111111011110111;
    rom[64727] = 25'b1111111111111111011111000;
    rom[64728] = 25'b1111111111111111011111000;
    rom[64729] = 25'b1111111111111111011111001;
    rom[64730] = 25'b1111111111111111011111001;
    rom[64731] = 25'b1111111111111111011111001;
    rom[64732] = 25'b1111111111111111011111001;
    rom[64733] = 25'b1111111111111111011111001;
    rom[64734] = 25'b1111111111111111011111010;
    rom[64735] = 25'b1111111111111111011111010;
    rom[64736] = 25'b1111111111111111011111011;
    rom[64737] = 25'b1111111111111111011111011;
    rom[64738] = 25'b1111111111111111011111100;
    rom[64739] = 25'b1111111111111111011111100;
    rom[64740] = 25'b1111111111111111011111100;
    rom[64741] = 25'b1111111111111111011111100;
    rom[64742] = 25'b1111111111111111011111100;
    rom[64743] = 25'b1111111111111111011111101;
    rom[64744] = 25'b1111111111111111011111101;
    rom[64745] = 25'b1111111111111111011111110;
    rom[64746] = 25'b1111111111111111011111110;
    rom[64747] = 25'b1111111111111111011111110;
    rom[64748] = 25'b1111111111111111011111110;
    rom[64749] = 25'b1111111111111111011111111;
    rom[64750] = 25'b1111111111111111011111111;
    rom[64751] = 25'b1111111111111111100000000;
    rom[64752] = 25'b1111111111111111100000000;
    rom[64753] = 25'b1111111111111111100000000;
    rom[64754] = 25'b1111111111111111100000001;
    rom[64755] = 25'b1111111111111111100000001;
    rom[64756] = 25'b1111111111111111100000001;
    rom[64757] = 25'b1111111111111111100000001;
    rom[64758] = 25'b1111111111111111100000010;
    rom[64759] = 25'b1111111111111111100000010;
    rom[64760] = 25'b1111111111111111100000011;
    rom[64761] = 25'b1111111111111111100000011;
    rom[64762] = 25'b1111111111111111100000100;
    rom[64763] = 25'b1111111111111111100000100;
    rom[64764] = 25'b1111111111111111100000100;
    rom[64765] = 25'b1111111111111111100000100;
    rom[64766] = 25'b1111111111111111100000100;
    rom[64767] = 25'b1111111111111111100000101;
    rom[64768] = 25'b1111111111111111100000101;
    rom[64769] = 25'b1111111111111111100000110;
    rom[64770] = 25'b1111111111111111100000110;
    rom[64771] = 25'b1111111111111111100000111;
    rom[64772] = 25'b1111111111111111100000111;
    rom[64773] = 25'b1111111111111111100000111;
    rom[64774] = 25'b1111111111111111100000111;
    rom[64775] = 25'b1111111111111111100000111;
    rom[64776] = 25'b1111111111111111100001000;
    rom[64777] = 25'b1111111111111111100001000;
    rom[64778] = 25'b1111111111111111100001001;
    rom[64779] = 25'b1111111111111111100001001;
    rom[64780] = 25'b1111111111111111100001010;
    rom[64781] = 25'b1111111111111111100001010;
    rom[64782] = 25'b1111111111111111100001010;
    rom[64783] = 25'b1111111111111111100001010;
    rom[64784] = 25'b1111111111111111100001010;
    rom[64785] = 25'b1111111111111111100001011;
    rom[64786] = 25'b1111111111111111100001011;
    rom[64787] = 25'b1111111111111111100001100;
    rom[64788] = 25'b1111111111111111100001100;
    rom[64789] = 25'b1111111111111111100001101;
    rom[64790] = 25'b1111111111111111100001101;
    rom[64791] = 25'b1111111111111111100001101;
    rom[64792] = 25'b1111111111111111100001101;
    rom[64793] = 25'b1111111111111111100001101;
    rom[64794] = 25'b1111111111111111100001110;
    rom[64795] = 25'b1111111111111111100001110;
    rom[64796] = 25'b1111111111111111100001111;
    rom[64797] = 25'b1111111111111111100001111;
    rom[64798] = 25'b1111111111111111100010000;
    rom[64799] = 25'b1111111111111111100010000;
    rom[64800] = 25'b1111111111111111100010000;
    rom[64801] = 25'b1111111111111111100010000;
    rom[64802] = 25'b1111111111111111100010000;
    rom[64803] = 25'b1111111111111111100010001;
    rom[64804] = 25'b1111111111111111100010001;
    rom[64805] = 25'b1111111111111111100010010;
    rom[64806] = 25'b1111111111111111100010010;
    rom[64807] = 25'b1111111111111111100010011;
    rom[64808] = 25'b1111111111111111100010011;
    rom[64809] = 25'b1111111111111111100010011;
    rom[64810] = 25'b1111111111111111100010011;
    rom[64811] = 25'b1111111111111111100010011;
    rom[64812] = 25'b1111111111111111100010100;
    rom[64813] = 25'b1111111111111111100010100;
    rom[64814] = 25'b1111111111111111100010101;
    rom[64815] = 25'b1111111111111111100010101;
    rom[64816] = 25'b1111111111111111100010110;
    rom[64817] = 25'b1111111111111111100010110;
    rom[64818] = 25'b1111111111111111100010110;
    rom[64819] = 25'b1111111111111111100010110;
    rom[64820] = 25'b1111111111111111100010110;
    rom[64821] = 25'b1111111111111111100010111;
    rom[64822] = 25'b1111111111111111100010111;
    rom[64823] = 25'b1111111111111111100011000;
    rom[64824] = 25'b1111111111111111100011000;
    rom[64825] = 25'b1111111111111111100011001;
    rom[64826] = 25'b1111111111111111100011001;
    rom[64827] = 25'b1111111111111111100011001;
    rom[64828] = 25'b1111111111111111100011001;
    rom[64829] = 25'b1111111111111111100011001;
    rom[64830] = 25'b1111111111111111100011010;
    rom[64831] = 25'b1111111111111111100011010;
    rom[64832] = 25'b1111111111111111100011011;
    rom[64833] = 25'b1111111111111111100011011;
    rom[64834] = 25'b1111111111111111100011011;
    rom[64835] = 25'b1111111111111111100011100;
    rom[64836] = 25'b1111111111111111100011100;
    rom[64837] = 25'b1111111111111111100011100;
    rom[64838] = 25'b1111111111111111100011100;
    rom[64839] = 25'b1111111111111111100011101;
    rom[64840] = 25'b1111111111111111100011101;
    rom[64841] = 25'b1111111111111111100011110;
    rom[64842] = 25'b1111111111111111100011110;
    rom[64843] = 25'b1111111111111111100011110;
    rom[64844] = 25'b1111111111111111100011111;
    rom[64845] = 25'b1111111111111111100011111;
    rom[64846] = 25'b1111111111111111100011111;
    rom[64847] = 25'b1111111111111111100011111;
    rom[64848] = 25'b1111111111111111100100000;
    rom[64849] = 25'b1111111111111111100100000;
    rom[64850] = 25'b1111111111111111100100000;
    rom[64851] = 25'b1111111111111111100100001;
    rom[64852] = 25'b1111111111111111100100001;
    rom[64853] = 25'b1111111111111111100100010;
    rom[64854] = 25'b1111111111111111100100010;
    rom[64855] = 25'b1111111111111111100100010;
    rom[64856] = 25'b1111111111111111100100010;
    rom[64857] = 25'b1111111111111111100100010;
    rom[64858] = 25'b1111111111111111100100011;
    rom[64859] = 25'b1111111111111111100100011;
    rom[64860] = 25'b1111111111111111100100100;
    rom[64861] = 25'b1111111111111111100100100;
    rom[64862] = 25'b1111111111111111100100101;
    rom[64863] = 25'b1111111111111111100100101;
    rom[64864] = 25'b1111111111111111100100101;
    rom[64865] = 25'b1111111111111111100100101;
    rom[64866] = 25'b1111111111111111100100101;
    rom[64867] = 25'b1111111111111111100100110;
    rom[64868] = 25'b1111111111111111100100110;
    rom[64869] = 25'b1111111111111111100100110;
    rom[64870] = 25'b1111111111111111100100111;
    rom[64871] = 25'b1111111111111111100100111;
    rom[64872] = 25'b1111111111111111100101000;
    rom[64873] = 25'b1111111111111111100101000;
    rom[64874] = 25'b1111111111111111100101000;
    rom[64875] = 25'b1111111111111111100101000;
    rom[64876] = 25'b1111111111111111100101000;
    rom[64877] = 25'b1111111111111111100101001;
    rom[64878] = 25'b1111111111111111100101001;
    rom[64879] = 25'b1111111111111111100101010;
    rom[64880] = 25'b1111111111111111100101010;
    rom[64881] = 25'b1111111111111111100101011;
    rom[64882] = 25'b1111111111111111100101011;
    rom[64883] = 25'b1111111111111111100101011;
    rom[64884] = 25'b1111111111111111100101011;
    rom[64885] = 25'b1111111111111111100101011;
    rom[64886] = 25'b1111111111111111100101100;
    rom[64887] = 25'b1111111111111111100101100;
    rom[64888] = 25'b1111111111111111100101100;
    rom[64889] = 25'b1111111111111111100101101;
    rom[64890] = 25'b1111111111111111100101101;
    rom[64891] = 25'b1111111111111111100101110;
    rom[64892] = 25'b1111111111111111100101110;
    rom[64893] = 25'b1111111111111111100101110;
    rom[64894] = 25'b1111111111111111100101110;
    rom[64895] = 25'b1111111111111111100101110;
    rom[64896] = 25'b1111111111111111100101111;
    rom[64897] = 25'b1111111111111111100101111;
    rom[64898] = 25'b1111111111111111100110000;
    rom[64899] = 25'b1111111111111111100110000;
    rom[64900] = 25'b1111111111111111100110000;
    rom[64901] = 25'b1111111111111111100110001;
    rom[64902] = 25'b1111111111111111100110001;
    rom[64903] = 25'b1111111111111111100110001;
    rom[64904] = 25'b1111111111111111100110001;
    rom[64905] = 25'b1111111111111111100110001;
    rom[64906] = 25'b1111111111111111100110010;
    rom[64907] = 25'b1111111111111111100110010;
    rom[64908] = 25'b1111111111111111100110011;
    rom[64909] = 25'b1111111111111111100110011;
    rom[64910] = 25'b1111111111111111100110100;
    rom[64911] = 25'b1111111111111111100110100;
    rom[64912] = 25'b1111111111111111100110100;
    rom[64913] = 25'b1111111111111111100110100;
    rom[64914] = 25'b1111111111111111100110100;
    rom[64915] = 25'b1111111111111111100110101;
    rom[64916] = 25'b1111111111111111100110101;
    rom[64917] = 25'b1111111111111111100110101;
    rom[64918] = 25'b1111111111111111100110110;
    rom[64919] = 25'b1111111111111111100110110;
    rom[64920] = 25'b1111111111111111100110111;
    rom[64921] = 25'b1111111111111111100110111;
    rom[64922] = 25'b1111111111111111100110111;
    rom[64923] = 25'b1111111111111111100110111;
    rom[64924] = 25'b1111111111111111100110111;
    rom[64925] = 25'b1111111111111111100111000;
    rom[64926] = 25'b1111111111111111100111000;
    rom[64927] = 25'b1111111111111111100111000;
    rom[64928] = 25'b1111111111111111100111001;
    rom[64929] = 25'b1111111111111111100111001;
    rom[64930] = 25'b1111111111111111100111010;
    rom[64931] = 25'b1111111111111111100111010;
    rom[64932] = 25'b1111111111111111100111010;
    rom[64933] = 25'b1111111111111111100111010;
    rom[64934] = 25'b1111111111111111100111010;
    rom[64935] = 25'b1111111111111111100111011;
    rom[64936] = 25'b1111111111111111100111011;
    rom[64937] = 25'b1111111111111111100111011;
    rom[64938] = 25'b1111111111111111100111100;
    rom[64939] = 25'b1111111111111111100111100;
    rom[64940] = 25'b1111111111111111100111101;
    rom[64941] = 25'b1111111111111111100111101;
    rom[64942] = 25'b1111111111111111100111101;
    rom[64943] = 25'b1111111111111111100111101;
    rom[64944] = 25'b1111111111111111100111101;
    rom[64945] = 25'b1111111111111111100111110;
    rom[64946] = 25'b1111111111111111100111110;
    rom[64947] = 25'b1111111111111111100111110;
    rom[64948] = 25'b1111111111111111100111111;
    rom[64949] = 25'b1111111111111111100111111;
    rom[64950] = 25'b1111111111111111100111111;
    rom[64951] = 25'b1111111111111111100111111;
    rom[64952] = 25'b1111111111111111100111111;
    rom[64953] = 25'b1111111111111111101000000;
    rom[64954] = 25'b1111111111111111101000000;
    rom[64955] = 25'b1111111111111111101000000;
    rom[64956] = 25'b1111111111111111101000001;
    rom[64957] = 25'b1111111111111111101000001;
    rom[64958] = 25'b1111111111111111101000010;
    rom[64959] = 25'b1111111111111111101000010;
    rom[64960] = 25'b1111111111111111101000010;
    rom[64961] = 25'b1111111111111111101000010;
    rom[64962] = 25'b1111111111111111101000010;
    rom[64963] = 25'b1111111111111111101000011;
    rom[64964] = 25'b1111111111111111101000011;
    rom[64965] = 25'b1111111111111111101000011;
    rom[64966] = 25'b1111111111111111101000100;
    rom[64967] = 25'b1111111111111111101000100;
    rom[64968] = 25'b1111111111111111101000101;
    rom[64969] = 25'b1111111111111111101000101;
    rom[64970] = 25'b1111111111111111101000101;
    rom[64971] = 25'b1111111111111111101000101;
    rom[64972] = 25'b1111111111111111101000101;
    rom[64973] = 25'b1111111111111111101000101;
    rom[64974] = 25'b1111111111111111101000110;
    rom[64975] = 25'b1111111111111111101000110;
    rom[64976] = 25'b1111111111111111101000111;
    rom[64977] = 25'b1111111111111111101000111;
    rom[64978] = 25'b1111111111111111101000111;
    rom[64979] = 25'b1111111111111111101001000;
    rom[64980] = 25'b1111111111111111101001000;
    rom[64981] = 25'b1111111111111111101001000;
    rom[64982] = 25'b1111111111111111101001000;
    rom[64983] = 25'b1111111111111111101001000;
    rom[64984] = 25'b1111111111111111101001001;
    rom[64985] = 25'b1111111111111111101001001;
    rom[64986] = 25'b1111111111111111101001001;
    rom[64987] = 25'b1111111111111111101001010;
    rom[64988] = 25'b1111111111111111101001010;
    rom[64989] = 25'b1111111111111111101001010;
    rom[64990] = 25'b1111111111111111101001011;
    rom[64991] = 25'b1111111111111111101001011;
    rom[64992] = 25'b1111111111111111101001011;
    rom[64993] = 25'b1111111111111111101001011;
    rom[64994] = 25'b1111111111111111101001011;
    rom[64995] = 25'b1111111111111111101001100;
    rom[64996] = 25'b1111111111111111101001100;
    rom[64997] = 25'b1111111111111111101001100;
    rom[64998] = 25'b1111111111111111101001101;
    rom[64999] = 25'b1111111111111111101001101;
    rom[65000] = 25'b1111111111111111101001110;
    rom[65001] = 25'b1111111111111111101001110;
    rom[65002] = 25'b1111111111111111101001110;
    rom[65003] = 25'b1111111111111111101001110;
    rom[65004] = 25'b1111111111111111101001110;
    rom[65005] = 25'b1111111111111111101001110;
    rom[65006] = 25'b1111111111111111101001111;
    rom[65007] = 25'b1111111111111111101001111;
    rom[65008] = 25'b1111111111111111101001111;
    rom[65009] = 25'b1111111111111111101010000;
    rom[65010] = 25'b1111111111111111101010000;
    rom[65011] = 25'b1111111111111111101010001;
    rom[65012] = 25'b1111111111111111101010001;
    rom[65013] = 25'b1111111111111111101010001;
    rom[65014] = 25'b1111111111111111101010001;
    rom[65015] = 25'b1111111111111111101010001;
    rom[65016] = 25'b1111111111111111101010001;
    rom[65017] = 25'b1111111111111111101010010;
    rom[65018] = 25'b1111111111111111101010010;
    rom[65019] = 25'b1111111111111111101010010;
    rom[65020] = 25'b1111111111111111101010011;
    rom[65021] = 25'b1111111111111111101010011;
    rom[65022] = 25'b1111111111111111101010100;
    rom[65023] = 25'b1111111111111111101010100;
    rom[65024] = 25'b1111111111111111101010100;
    rom[65025] = 25'b1111111111111111101010100;
    rom[65026] = 25'b1111111111111111101010100;
    rom[65027] = 25'b1111111111111111101010100;
    rom[65028] = 25'b1111111111111111101010101;
    rom[65029] = 25'b1111111111111111101010101;
    rom[65030] = 25'b1111111111111111101010101;
    rom[65031] = 25'b1111111111111111101010110;
    rom[65032] = 25'b1111111111111111101010110;
    rom[65033] = 25'b1111111111111111101010110;
    rom[65034] = 25'b1111111111111111101010111;
    rom[65035] = 25'b1111111111111111101010111;
    rom[65036] = 25'b1111111111111111101010111;
    rom[65037] = 25'b1111111111111111101010111;
    rom[65038] = 25'b1111111111111111101010111;
    rom[65039] = 25'b1111111111111111101011000;
    rom[65040] = 25'b1111111111111111101011000;
    rom[65041] = 25'b1111111111111111101011000;
    rom[65042] = 25'b1111111111111111101011001;
    rom[65043] = 25'b1111111111111111101011001;
    rom[65044] = 25'b1111111111111111101011001;
    rom[65045] = 25'b1111111111111111101011010;
    rom[65046] = 25'b1111111111111111101011010;
    rom[65047] = 25'b1111111111111111101011010;
    rom[65048] = 25'b1111111111111111101011010;
    rom[65049] = 25'b1111111111111111101011010;
    rom[65050] = 25'b1111111111111111101011010;
    rom[65051] = 25'b1111111111111111101011011;
    rom[65052] = 25'b1111111111111111101011011;
    rom[65053] = 25'b1111111111111111101011011;
    rom[65054] = 25'b1111111111111111101011100;
    rom[65055] = 25'b1111111111111111101011100;
    rom[65056] = 25'b1111111111111111101011100;
    rom[65057] = 25'b1111111111111111101011101;
    rom[65058] = 25'b1111111111111111101011101;
    rom[65059] = 25'b1111111111111111101011101;
    rom[65060] = 25'b1111111111111111101011101;
    rom[65061] = 25'b1111111111111111101011101;
    rom[65062] = 25'b1111111111111111101011101;
    rom[65063] = 25'b1111111111111111101011110;
    rom[65064] = 25'b1111111111111111101011110;
    rom[65065] = 25'b1111111111111111101011110;
    rom[65066] = 25'b1111111111111111101011111;
    rom[65067] = 25'b1111111111111111101011111;
    rom[65068] = 25'b1111111111111111101011111;
    rom[65069] = 25'b1111111111111111101100000;
    rom[65070] = 25'b1111111111111111101100000;
    rom[65071] = 25'b1111111111111111101100000;
    rom[65072] = 25'b1111111111111111101100000;
    rom[65073] = 25'b1111111111111111101100000;
    rom[65074] = 25'b1111111111111111101100000;
    rom[65075] = 25'b1111111111111111101100001;
    rom[65076] = 25'b1111111111111111101100001;
    rom[65077] = 25'b1111111111111111101100001;
    rom[65078] = 25'b1111111111111111101100010;
    rom[65079] = 25'b1111111111111111101100010;
    rom[65080] = 25'b1111111111111111101100010;
    rom[65081] = 25'b1111111111111111101100011;
    rom[65082] = 25'b1111111111111111101100011;
    rom[65083] = 25'b1111111111111111101100011;
    rom[65084] = 25'b1111111111111111101100011;
    rom[65085] = 25'b1111111111111111101100011;
    rom[65086] = 25'b1111111111111111101100011;
    rom[65087] = 25'b1111111111111111101100100;
    rom[65088] = 25'b1111111111111111101100100;
    rom[65089] = 25'b1111111111111111101100100;
    rom[65090] = 25'b1111111111111111101100101;
    rom[65091] = 25'b1111111111111111101100101;
    rom[65092] = 25'b1111111111111111101100101;
    rom[65093] = 25'b1111111111111111101100101;
    rom[65094] = 25'b1111111111111111101100110;
    rom[65095] = 25'b1111111111111111101100110;
    rom[65096] = 25'b1111111111111111101100110;
    rom[65097] = 25'b1111111111111111101100110;
    rom[65098] = 25'b1111111111111111101100110;
    rom[65099] = 25'b1111111111111111101100110;
    rom[65100] = 25'b1111111111111111101100111;
    rom[65101] = 25'b1111111111111111101100111;
    rom[65102] = 25'b1111111111111111101100111;
    rom[65103] = 25'b1111111111111111101101000;
    rom[65104] = 25'b1111111111111111101101000;
    rom[65105] = 25'b1111111111111111101101000;
    rom[65106] = 25'b1111111111111111101101001;
    rom[65107] = 25'b1111111111111111101101001;
    rom[65108] = 25'b1111111111111111101101001;
    rom[65109] = 25'b1111111111111111101101001;
    rom[65110] = 25'b1111111111111111101101001;
    rom[65111] = 25'b1111111111111111101101001;
    rom[65112] = 25'b1111111111111111101101001;
    rom[65113] = 25'b1111111111111111101101010;
    rom[65114] = 25'b1111111111111111101101010;
    rom[65115] = 25'b1111111111111111101101010;
    rom[65116] = 25'b1111111111111111101101011;
    rom[65117] = 25'b1111111111111111101101011;
    rom[65118] = 25'b1111111111111111101101011;
    rom[65119] = 25'b1111111111111111101101100;
    rom[65120] = 25'b1111111111111111101101100;
    rom[65121] = 25'b1111111111111111101101100;
    rom[65122] = 25'b1111111111111111101101100;
    rom[65123] = 25'b1111111111111111101101100;
    rom[65124] = 25'b1111111111111111101101100;
    rom[65125] = 25'b1111111111111111101101100;
    rom[65126] = 25'b1111111111111111101101101;
    rom[65127] = 25'b1111111111111111101101101;
    rom[65128] = 25'b1111111111111111101101101;
    rom[65129] = 25'b1111111111111111101101110;
    rom[65130] = 25'b1111111111111111101101110;
    rom[65131] = 25'b1111111111111111101101110;
    rom[65132] = 25'b1111111111111111101101110;
    rom[65133] = 25'b1111111111111111101101111;
    rom[65134] = 25'b1111111111111111101101111;
    rom[65135] = 25'b1111111111111111101101111;
    rom[65136] = 25'b1111111111111111101101111;
    rom[65137] = 25'b1111111111111111101101111;
    rom[65138] = 25'b1111111111111111101101111;
    rom[65139] = 25'b1111111111111111101101111;
    rom[65140] = 25'b1111111111111111101110000;
    rom[65141] = 25'b1111111111111111101110000;
    rom[65142] = 25'b1111111111111111101110000;
    rom[65143] = 25'b1111111111111111101110001;
    rom[65144] = 25'b1111111111111111101110001;
    rom[65145] = 25'b1111111111111111101110001;
    rom[65146] = 25'b1111111111111111101110010;
    rom[65147] = 25'b1111111111111111101110010;
    rom[65148] = 25'b1111111111111111101110010;
    rom[65149] = 25'b1111111111111111101110010;
    rom[65150] = 25'b1111111111111111101110010;
    rom[65151] = 25'b1111111111111111101110010;
    rom[65152] = 25'b1111111111111111101110010;
    rom[65153] = 25'b1111111111111111101110010;
    rom[65154] = 25'b1111111111111111101110011;
    rom[65155] = 25'b1111111111111111101110011;
    rom[65156] = 25'b1111111111111111101110011;
    rom[65157] = 25'b1111111111111111101110100;
    rom[65158] = 25'b1111111111111111101110100;
    rom[65159] = 25'b1111111111111111101110100;
    rom[65160] = 25'b1111111111111111101110100;
    rom[65161] = 25'b1111111111111111101110101;
    rom[65162] = 25'b1111111111111111101110101;
    rom[65163] = 25'b1111111111111111101110101;
    rom[65164] = 25'b1111111111111111101110101;
    rom[65165] = 25'b1111111111111111101110101;
    rom[65166] = 25'b1111111111111111101110101;
    rom[65167] = 25'b1111111111111111101110101;
    rom[65168] = 25'b1111111111111111101110110;
    rom[65169] = 25'b1111111111111111101110110;
    rom[65170] = 25'b1111111111111111101110110;
    rom[65171] = 25'b1111111111111111101110110;
    rom[65172] = 25'b1111111111111111101110111;
    rom[65173] = 25'b1111111111111111101110111;
    rom[65174] = 25'b1111111111111111101110111;
    rom[65175] = 25'b1111111111111111101111000;
    rom[65176] = 25'b1111111111111111101111000;
    rom[65177] = 25'b1111111111111111101111000;
    rom[65178] = 25'b1111111111111111101111000;
    rom[65179] = 25'b1111111111111111101111000;
    rom[65180] = 25'b1111111111111111101111000;
    rom[65181] = 25'b1111111111111111101111000;
    rom[65182] = 25'b1111111111111111101111000;
    rom[65183] = 25'b1111111111111111101111001;
    rom[65184] = 25'b1111111111111111101111001;
    rom[65185] = 25'b1111111111111111101111001;
    rom[65186] = 25'b1111111111111111101111001;
    rom[65187] = 25'b1111111111111111101111010;
    rom[65188] = 25'b1111111111111111101111010;
    rom[65189] = 25'b1111111111111111101111010;
    rom[65190] = 25'b1111111111111111101111010;
    rom[65191] = 25'b1111111111111111101111011;
    rom[65192] = 25'b1111111111111111101111011;
    rom[65193] = 25'b1111111111111111101111011;
    rom[65194] = 25'b1111111111111111101111011;
    rom[65195] = 25'b1111111111111111101111011;
    rom[65196] = 25'b1111111111111111101111011;
    rom[65197] = 25'b1111111111111111101111011;
    rom[65198] = 25'b1111111111111111101111011;
    rom[65199] = 25'b1111111111111111101111100;
    rom[65200] = 25'b1111111111111111101111100;
    rom[65201] = 25'b1111111111111111101111100;
    rom[65202] = 25'b1111111111111111101111101;
    rom[65203] = 25'b1111111111111111101111101;
    rom[65204] = 25'b1111111111111111101111101;
    rom[65205] = 25'b1111111111111111101111101;
    rom[65206] = 25'b1111111111111111101111101;
    rom[65207] = 25'b1111111111111111101111110;
    rom[65208] = 25'b1111111111111111101111110;
    rom[65209] = 25'b1111111111111111101111110;
    rom[65210] = 25'b1111111111111111101111110;
    rom[65211] = 25'b1111111111111111101111110;
    rom[65212] = 25'b1111111111111111101111110;
    rom[65213] = 25'b1111111111111111101111110;
    rom[65214] = 25'b1111111111111111101111110;
    rom[65215] = 25'b1111111111111111101111111;
    rom[65216] = 25'b1111111111111111101111111;
    rom[65217] = 25'b1111111111111111101111111;
    rom[65218] = 25'b1111111111111111101111111;
    rom[65219] = 25'b1111111111111111110000000;
    rom[65220] = 25'b1111111111111111110000000;
    rom[65221] = 25'b1111111111111111110000000;
    rom[65222] = 25'b1111111111111111110000000;
    rom[65223] = 25'b1111111111111111110000000;
    rom[65224] = 25'b1111111111111111110000000;
    rom[65225] = 25'b1111111111111111110000000;
    rom[65226] = 25'b1111111111111111110000000;
    rom[65227] = 25'b1111111111111111110000001;
    rom[65228] = 25'b1111111111111111110000001;
    rom[65229] = 25'b1111111111111111110000001;
    rom[65230] = 25'b1111111111111111110000001;
    rom[65231] = 25'b1111111111111111110000001;
    rom[65232] = 25'b1111111111111111110000010;
    rom[65233] = 25'b1111111111111111110000010;
    rom[65234] = 25'b1111111111111111110000010;
    rom[65235] = 25'b1111111111111111110000010;
    rom[65236] = 25'b1111111111111111110000011;
    rom[65237] = 25'b1111111111111111110000011;
    rom[65238] = 25'b1111111111111111110000011;
    rom[65239] = 25'b1111111111111111110000011;
    rom[65240] = 25'b1111111111111111110000011;
    rom[65241] = 25'b1111111111111111110000011;
    rom[65242] = 25'b1111111111111111110000011;
    rom[65243] = 25'b1111111111111111110000011;
    rom[65244] = 25'b1111111111111111110000011;
    rom[65245] = 25'b1111111111111111110000100;
    rom[65246] = 25'b1111111111111111110000100;
    rom[65247] = 25'b1111111111111111110000100;
    rom[65248] = 25'b1111111111111111110000100;
    rom[65249] = 25'b1111111111111111110000100;
    rom[65250] = 25'b1111111111111111110000101;
    rom[65251] = 25'b1111111111111111110000101;
    rom[65252] = 25'b1111111111111111110000101;
    rom[65253] = 25'b1111111111111111110000101;
    rom[65254] = 25'b1111111111111111110000110;
    rom[65255] = 25'b1111111111111111110000110;
    rom[65256] = 25'b1111111111111111110000110;
    rom[65257] = 25'b1111111111111111110000110;
    rom[65258] = 25'b1111111111111111110000110;
    rom[65259] = 25'b1111111111111111110000110;
    rom[65260] = 25'b1111111111111111110000110;
    rom[65261] = 25'b1111111111111111110000110;
    rom[65262] = 25'b1111111111111111110000110;
    rom[65263] = 25'b1111111111111111110000110;
    rom[65264] = 25'b1111111111111111110000111;
    rom[65265] = 25'b1111111111111111110000111;
    rom[65266] = 25'b1111111111111111110000111;
    rom[65267] = 25'b1111111111111111110000111;
    rom[65268] = 25'b1111111111111111110000111;
    rom[65269] = 25'b1111111111111111110001000;
    rom[65270] = 25'b1111111111111111110001000;
    rom[65271] = 25'b1111111111111111110001000;
    rom[65272] = 25'b1111111111111111110001000;
    rom[65273] = 25'b1111111111111111110001000;
    rom[65274] = 25'b1111111111111111110001001;
    rom[65275] = 25'b1111111111111111110001001;
    rom[65276] = 25'b1111111111111111110001001;
    rom[65277] = 25'b1111111111111111110001001;
    rom[65278] = 25'b1111111111111111110001001;
    rom[65279] = 25'b1111111111111111110001001;
    rom[65280] = 25'b1111111111111111110001001;
    rom[65281] = 25'b1111111111111111110001001;
    rom[65282] = 25'b1111111111111111110001001;
    rom[65283] = 25'b1111111111111111110001001;
    rom[65284] = 25'b1111111111111111110001010;
    rom[65285] = 25'b1111111111111111110001010;
    rom[65286] = 25'b1111111111111111110001010;
    rom[65287] = 25'b1111111111111111110001010;
    rom[65288] = 25'b1111111111111111110001010;
    rom[65289] = 25'b1111111111111111110001011;
    rom[65290] = 25'b1111111111111111110001011;
    rom[65291] = 25'b1111111111111111110001011;
    rom[65292] = 25'b1111111111111111110001011;
    rom[65293] = 25'b1111111111111111110001011;
    rom[65294] = 25'b1111111111111111110001100;
    rom[65295] = 25'b1111111111111111110001100;
    rom[65296] = 25'b1111111111111111110001100;
    rom[65297] = 25'b1111111111111111110001100;
    rom[65298] = 25'b1111111111111111110001100;
    rom[65299] = 25'b1111111111111111110001100;
    rom[65300] = 25'b1111111111111111110001100;
    rom[65301] = 25'b1111111111111111110001100;
    rom[65302] = 25'b1111111111111111110001100;
    rom[65303] = 25'b1111111111111111110001100;
    rom[65304] = 25'b1111111111111111110001100;
    rom[65305] = 25'b1111111111111111110001101;
    rom[65306] = 25'b1111111111111111110001101;
    rom[65307] = 25'b1111111111111111110001101;
    rom[65308] = 25'b1111111111111111110001101;
    rom[65309] = 25'b1111111111111111110001101;
    rom[65310] = 25'b1111111111111111110001101;
    rom[65311] = 25'b1111111111111111110001110;
    rom[65312] = 25'b1111111111111111110001110;
    rom[65313] = 25'b1111111111111111110001110;
    rom[65314] = 25'b1111111111111111110001110;
    rom[65315] = 25'b1111111111111111110001110;
    rom[65316] = 25'b1111111111111111110001110;
    rom[65317] = 25'b1111111111111111110001111;
    rom[65318] = 25'b1111111111111111110001111;
    rom[65319] = 25'b1111111111111111110001111;
    rom[65320] = 25'b1111111111111111110001111;
    rom[65321] = 25'b1111111111111111110001111;
    rom[65322] = 25'b1111111111111111110001111;
    rom[65323] = 25'b1111111111111111110001111;
    rom[65324] = 25'b1111111111111111110001111;
    rom[65325] = 25'b1111111111111111110001111;
    rom[65326] = 25'b1111111111111111110001111;
    rom[65327] = 25'b1111111111111111110001111;
    rom[65328] = 25'b1111111111111111110001111;
    rom[65329] = 25'b1111111111111111110010000;
    rom[65330] = 25'b1111111111111111110010000;
    rom[65331] = 25'b1111111111111111110010000;
    rom[65332] = 25'b1111111111111111110010000;
    rom[65333] = 25'b1111111111111111110010000;
    rom[65334] = 25'b1111111111111111110010000;
    rom[65335] = 25'b1111111111111111110010001;
    rom[65336] = 25'b1111111111111111110010001;
    rom[65337] = 25'b1111111111111111110010001;
    rom[65338] = 25'b1111111111111111110010001;
    rom[65339] = 25'b1111111111111111110010001;
    rom[65340] = 25'b1111111111111111110010001;
    rom[65341] = 25'b1111111111111111110010001;
    rom[65342] = 25'b1111111111111111110010010;
    rom[65343] = 25'b1111111111111111110010010;
    rom[65344] = 25'b1111111111111111110010010;
    rom[65345] = 25'b1111111111111111110010010;
    rom[65346] = 25'b1111111111111111110010010;
    rom[65347] = 25'b1111111111111111110010010;
    rom[65348] = 25'b1111111111111111110010010;
    rom[65349] = 25'b1111111111111111110010010;
    rom[65350] = 25'b1111111111111111110010010;
    rom[65351] = 25'b1111111111111111110010010;
    rom[65352] = 25'b1111111111111111110010010;
    rom[65353] = 25'b1111111111111111110010010;
    rom[65354] = 25'b1111111111111111110010010;
    rom[65355] = 25'b1111111111111111110010010;
    rom[65356] = 25'b1111111111111111110010011;
    rom[65357] = 25'b1111111111111111110010011;
    rom[65358] = 25'b1111111111111111110010011;
    rom[65359] = 25'b1111111111111111110010011;
    rom[65360] = 25'b1111111111111111110010011;
    rom[65361] = 25'b1111111111111111110010011;
    rom[65362] = 25'b1111111111111111110010011;
    rom[65363] = 25'b1111111111111111110010100;
    rom[65364] = 25'b1111111111111111110010100;
    rom[65365] = 25'b1111111111111111110010100;
    rom[65366] = 25'b1111111111111111110010100;
    rom[65367] = 25'b1111111111111111110010100;
    rom[65368] = 25'b1111111111111111110010100;
    rom[65369] = 25'b1111111111111111110010100;
    rom[65370] = 25'b1111111111111111110010100;
    rom[65371] = 25'b1111111111111111110010101;
    rom[65372] = 25'b1111111111111111110010101;
    rom[65373] = 25'b1111111111111111110010101;
    rom[65374] = 25'b1111111111111111110010101;
    rom[65375] = 25'b1111111111111111110010101;
    rom[65376] = 25'b1111111111111111110010101;
    rom[65377] = 25'b1111111111111111110010101;
    rom[65378] = 25'b1111111111111111110010101;
    rom[65379] = 25'b1111111111111111110010101;
    rom[65380] = 25'b1111111111111111110010101;
    rom[65381] = 25'b1111111111111111110010101;
    rom[65382] = 25'b1111111111111111110010101;
    rom[65383] = 25'b1111111111111111110010101;
    rom[65384] = 25'b1111111111111111110010101;
    rom[65385] = 25'b1111111111111111110010101;
    rom[65386] = 25'b1111111111111111110010101;
    rom[65387] = 25'b1111111111111111110010110;
    rom[65388] = 25'b1111111111111111110010110;
    rom[65389] = 25'b1111111111111111110010110;
    rom[65390] = 25'b1111111111111111110010110;
    rom[65391] = 25'b1111111111111111110010110;
    rom[65392] = 25'b1111111111111111110010110;
    rom[65393] = 25'b1111111111111111110010110;
    rom[65394] = 25'b1111111111111111110010110;
    rom[65395] = 25'b1111111111111111110010110;
    rom[65396] = 25'b1111111111111111110010111;
    rom[65397] = 25'b1111111111111111110010111;
    rom[65398] = 25'b1111111111111111110010111;
    rom[65399] = 25'b1111111111111111110010111;
    rom[65400] = 25'b1111111111111111110010111;
    rom[65401] = 25'b1111111111111111110010111;
    rom[65402] = 25'b1111111111111111110010111;
    rom[65403] = 25'b1111111111111111110010111;
    rom[65404] = 25'b1111111111111111110010111;
    rom[65405] = 25'b1111111111111111110011000;
    rom[65406] = 25'b1111111111111111110011000;
    rom[65407] = 25'b1111111111111111110011000;
    rom[65408] = 25'b1111111111111111110011000;
    rom[65409] = 25'b1111111111111111110011000;
    rom[65410] = 25'b1111111111111111110011000;
    rom[65411] = 25'b1111111111111111110011000;
    rom[65412] = 25'b1111111111111111110011000;
    rom[65413] = 25'b1111111111111111110011000;
    rom[65414] = 25'b1111111111111111110011000;
    rom[65415] = 25'b1111111111111111110011000;
    rom[65416] = 25'b1111111111111111110011000;
    rom[65417] = 25'b1111111111111111110011000;
    rom[65418] = 25'b1111111111111111110011000;
    rom[65419] = 25'b1111111111111111110011000;
    rom[65420] = 25'b1111111111111111110011000;
    rom[65421] = 25'b1111111111111111110011000;
    rom[65422] = 25'b1111111111111111110011000;
    rom[65423] = 25'b1111111111111111110011000;
    rom[65424] = 25'b1111111111111111110011000;
    rom[65425] = 25'b1111111111111111110011000;
    rom[65426] = 25'b1111111111111111110011000;
    rom[65427] = 25'b1111111111111111110011001;
    rom[65428] = 25'b1111111111111111110011001;
    rom[65429] = 25'b1111111111111111110011001;
    rom[65430] = 25'b1111111111111111110011001;
    rom[65431] = 25'b1111111111111111110011001;
    rom[65432] = 25'b1111111111111111110011001;
    rom[65433] = 25'b1111111111111111110011001;
    rom[65434] = 25'b1111111111111111110011001;
    rom[65435] = 25'b1111111111111111110011001;
    rom[65436] = 25'b1111111111111111110011001;
    rom[65437] = 25'b1111111111111111110011001;
    rom[65438] = 25'b1111111111111111110011001;
    rom[65439] = 25'b1111111111111111110011010;
    rom[65440] = 25'b1111111111111111110011010;
    rom[65441] = 25'b1111111111111111110011010;
    rom[65442] = 25'b1111111111111111110011010;
    rom[65443] = 25'b1111111111111111110011010;
    rom[65444] = 25'b1111111111111111110011010;
    rom[65445] = 25'b1111111111111111110011010;
    rom[65446] = 25'b1111111111111111110011010;
    rom[65447] = 25'b1111111111111111110011010;
    rom[65448] = 25'b1111111111111111110011010;
    rom[65449] = 25'b1111111111111111110011010;
    rom[65450] = 25'b1111111111111111110011010;
    rom[65451] = 25'b1111111111111111110011010;
    rom[65452] = 25'b1111111111111111110011010;
    rom[65453] = 25'b1111111111111111110011011;
    rom[65454] = 25'b1111111111111111110011011;
    rom[65455] = 25'b1111111111111111110011011;
    rom[65456] = 25'b1111111111111111110011011;
    rom[65457] = 25'b1111111111111111110011011;
    rom[65458] = 25'b1111111111111111110011011;
    rom[65459] = 25'b1111111111111111110011011;
    rom[65460] = 25'b1111111111111111110011011;
    rom[65461] = 25'b1111111111111111110011011;
    rom[65462] = 25'b1111111111111111110011011;
    rom[65463] = 25'b1111111111111111110011011;
    rom[65464] = 25'b1111111111111111110011011;
    rom[65465] = 25'b1111111111111111110011011;
    rom[65466] = 25'b1111111111111111110011011;
    rom[65467] = 25'b1111111111111111110011011;
    rom[65468] = 25'b1111111111111111110011011;
    rom[65469] = 25'b1111111111111111110011011;
    rom[65470] = 25'b1111111111111111110011011;
    rom[65471] = 25'b1111111111111111110011011;
    rom[65472] = 25'b1111111111111111110011011;
    rom[65473] = 25'b1111111111111111110011011;
    rom[65474] = 25'b1111111111111111110011011;
    rom[65475] = 25'b1111111111111111110011011;
    rom[65476] = 25'b1111111111111111110011011;
    rom[65477] = 25'b1111111111111111110011011;
    rom[65478] = 25'b1111111111111111110011011;
    rom[65479] = 25'b1111111111111111110011011;
    rom[65480] = 25'b1111111111111111110011011;
    rom[65481] = 25'b1111111111111111110011011;
    rom[65482] = 25'b1111111111111111110011011;
    rom[65483] = 25'b1111111111111111110011011;
    rom[65484] = 25'b1111111111111111110011011;
    rom[65485] = 25'b1111111111111111110011011;
    rom[65486] = 25'b1111111111111111110011011;
    rom[65487] = 25'b1111111111111111110011011;
    rom[65488] = 25'b1111111111111111110011011;
    rom[65489] = 25'b1111111111111111110011011;
    rom[65490] = 25'b1111111111111111110011011;
    rom[65491] = 25'b1111111111111111110011011;
    rom[65492] = 25'b1111111111111111110011011;
    rom[65493] = 25'b1111111111111111110011100;
    rom[65494] = 25'b1111111111111111110011100;
    rom[65495] = 25'b1111111111111111110011100;
    rom[65496] = 25'b1111111111111111110011100;
    rom[65497] = 25'b1111111111111111110011100;
    rom[65498] = 25'b1111111111111111110011100;
    rom[65499] = 25'b1111111111111111110011100;
    rom[65500] = 25'b1111111111111111110011100;
    rom[65501] = 25'b1111111111111111110011100;
    rom[65502] = 25'b1111111111111111110011100;
    rom[65503] = 25'b1111111111111111110011100;
    rom[65504] = 25'b1111111111111111110011100;
    rom[65505] = 25'b1111111111111111110011100;
    rom[65506] = 25'b1111111111111111110011100;
    rom[65507] = 25'b1111111111111111110011100;
    rom[65508] = 25'b1111111111111111110011100;
    rom[65509] = 25'b1111111111111111110011100;
    rom[65510] = 25'b1111111111111111110011100;
    rom[65511] = 25'b1111111111111111110011100;
    rom[65512] = 25'b1111111111111111110011100;
    rom[65513] = 25'b1111111111111111110011100;
    rom[65514] = 25'b1111111111111111110011100;
    rom[65515] = 25'b1111111111111111110011100;
    rom[65516] = 25'b1111111111111111110011100;
    rom[65517] = 25'b1111111111111111110011100;
    rom[65518] = 25'b1111111111111111110011100;
    rom[65519] = 25'b1111111111111111110011100;
    rom[65520] = 25'b1111111111111111110011100;
    rom[65521] = 25'b1111111111111111110011100;
    rom[65522] = 25'b1111111111111111110011100;
    rom[65523] = 25'b1111111111111111110011100;
    rom[65524] = 25'b1111111111111111110011100;
    rom[65525] = 25'b1111111111111111110011100;
    rom[65526] = 25'b1111111111111111110011100;
    rom[65527] = 25'b1111111111111111110011100;
    rom[65528] = 25'b1111111111111111110011100;
    rom[65529] = 25'b1111111111111111110011100;
    rom[65530] = 25'b1111111111111111110011100;
    rom[65531] = 25'b1111111111111111110011100;
    rom[65532] = 25'b1111111111111111110011100;
    rom[65533] = 25'b1111111111111111110011100;
    rom[65534] = 25'b1111111111111111110011100;
    rom[65535] = 25'b1111111111111111110011100;
end

// port a
always @(posedge clk)
begin
    if (wea_d == 1'b1) begin
      rom[addra_d] <= dia_d;
    end
    wea_d <= wea;
    dia_d <= dia;
    addra_d <= addra;
end

// port b
always @(posedge clk)
begin
    addrb_d <= addrb;
    rom_pipea <= rom[addrb_d];
    dob_d <= rom_pipea;
end

endmodule
