
/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : cic_M256_N1_R1_iw5_0_offset_sp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data                                                     
//
//
/*****************************************************************************/


module cic_M256_N1_R1_iw5_0_offset_sp_rom
(
  input clk, 

  input [8:0] addra,
  output [0:0] doa
);

(* rom_style = "distributed" *) reg [0:0] rom [511:0];
reg [8:0] addra_d;
reg [0:0] doa_d;
reg [0:0] rom_pipea;

assign doa = doa_d;

initial
begin
    rom[0] = 1'b0;
    rom[1] = 1'b0;
    rom[2] = 1'b0;
    rom[3] = 1'b0;
    rom[4] = 1'b0;
    rom[5] = 1'b0;
    rom[6] = 1'b0;
    rom[7] = 1'b0;
    rom[8] = 1'b0;
    rom[9] = 1'b0;
    rom[10] = 1'b0;
    rom[11] = 1'b0;
    rom[12] = 1'b0;
    rom[13] = 1'b0;
    rom[14] = 1'b0;
    rom[15] = 1'b0;
    rom[16] = 1'b0;
    rom[17] = 1'b0;
    rom[18] = 1'b0;
    rom[19] = 1'b0;
    rom[20] = 1'b0;
    rom[21] = 1'b0;
    rom[22] = 1'b0;
    rom[23] = 1'b0;
    rom[24] = 1'b0;
    rom[25] = 1'b0;
    rom[26] = 1'b0;
    rom[27] = 1'b0;
    rom[28] = 1'b0;
    rom[29] = 1'b0;
    rom[30] = 1'b0;
    rom[31] = 1'b0;
    rom[32] = 1'b0;
    rom[33] = 1'b0;
    rom[34] = 1'b0;
    rom[35] = 1'b0;
    rom[36] = 1'b0;
    rom[37] = 1'b0;
    rom[38] = 1'b0;
    rom[39] = 1'b0;
    rom[40] = 1'b0;
    rom[41] = 1'b0;
    rom[42] = 1'b0;
    rom[43] = 1'b0;
    rom[44] = 1'b0;
    rom[45] = 1'b0;
    rom[46] = 1'b0;
    rom[47] = 1'b0;
    rom[48] = 1'b0;
    rom[49] = 1'b0;
    rom[50] = 1'b0;
    rom[51] = 1'b0;
    rom[52] = 1'b0;
    rom[53] = 1'b0;
    rom[54] = 1'b0;
    rom[55] = 1'b0;
    rom[56] = 1'b0;
    rom[57] = 1'b0;
    rom[58] = 1'b0;
    rom[59] = 1'b0;
    rom[60] = 1'b0;
    rom[61] = 1'b0;
    rom[62] = 1'b0;
    rom[63] = 1'b0;
    rom[64] = 1'b0;
    rom[65] = 1'b0;
    rom[66] = 1'b0;
    rom[67] = 1'b0;
    rom[68] = 1'b0;
    rom[69] = 1'b0;
    rom[70] = 1'b0;
    rom[71] = 1'b0;
    rom[72] = 1'b0;
    rom[73] = 1'b0;
    rom[74] = 1'b0;
    rom[75] = 1'b0;
    rom[76] = 1'b0;
    rom[77] = 1'b0;
    rom[78] = 1'b0;
    rom[79] = 1'b0;
    rom[80] = 1'b0;
    rom[81] = 1'b0;
    rom[82] = 1'b0;
    rom[83] = 1'b0;
    rom[84] = 1'b0;
    rom[85] = 1'b0;
    rom[86] = 1'b0;
    rom[87] = 1'b0;
    rom[88] = 1'b0;
    rom[89] = 1'b0;
    rom[90] = 1'b0;
    rom[91] = 1'b0;
    rom[92] = 1'b0;
    rom[93] = 1'b0;
    rom[94] = 1'b0;
    rom[95] = 1'b0;
    rom[96] = 1'b0;
    rom[97] = 1'b0;
    rom[98] = 1'b0;
    rom[99] = 1'b0;
    rom[100] = 1'b0;
    rom[101] = 1'b0;
    rom[102] = 1'b0;
    rom[103] = 1'b0;
    rom[104] = 1'b0;
    rom[105] = 1'b0;
    rom[106] = 1'b0;
    rom[107] = 1'b0;
    rom[108] = 1'b0;
    rom[109] = 1'b0;
    rom[110] = 1'b0;
    rom[111] = 1'b0;
    rom[112] = 1'b0;
    rom[113] = 1'b0;
    rom[114] = 1'b0;
    rom[115] = 1'b0;
    rom[116] = 1'b0;
    rom[117] = 1'b0;
    rom[118] = 1'b0;
    rom[119] = 1'b0;
    rom[120] = 1'b0;
    rom[121] = 1'b0;
    rom[122] = 1'b0;
    rom[123] = 1'b0;
    rom[124] = 1'b0;
    rom[125] = 1'b0;
    rom[126] = 1'b0;
    rom[127] = 1'b0;
    rom[128] = 1'b0;
    rom[129] = 1'b0;
    rom[130] = 1'b0;
    rom[131] = 1'b0;
    rom[132] = 1'b0;
    rom[133] = 1'b0;
    rom[134] = 1'b0;
    rom[135] = 1'b0;
    rom[136] = 1'b0;
    rom[137] = 1'b0;
    rom[138] = 1'b0;
    rom[139] = 1'b0;
    rom[140] = 1'b0;
    rom[141] = 1'b0;
    rom[142] = 1'b0;
    rom[143] = 1'b0;
    rom[144] = 1'b0;
    rom[145] = 1'b0;
    rom[146] = 1'b0;
    rom[147] = 1'b0;
    rom[148] = 1'b0;
    rom[149] = 1'b0;
    rom[150] = 1'b0;
    rom[151] = 1'b0;
    rom[152] = 1'b0;
    rom[153] = 1'b0;
    rom[154] = 1'b0;
    rom[155] = 1'b0;
    rom[156] = 1'b0;
    rom[157] = 1'b0;
    rom[158] = 1'b0;
    rom[159] = 1'b0;
    rom[160] = 1'b0;
    rom[161] = 1'b0;
    rom[162] = 1'b0;
    rom[163] = 1'b0;
    rom[164] = 1'b0;
    rom[165] = 1'b0;
    rom[166] = 1'b0;
    rom[167] = 1'b0;
    rom[168] = 1'b0;
    rom[169] = 1'b0;
    rom[170] = 1'b0;
    rom[171] = 1'b0;
    rom[172] = 1'b0;
    rom[173] = 1'b0;
    rom[174] = 1'b0;
    rom[175] = 1'b0;
    rom[176] = 1'b0;
    rom[177] = 1'b0;
    rom[178] = 1'b0;
    rom[179] = 1'b0;
    rom[180] = 1'b0;
    rom[181] = 1'b0;
    rom[182] = 1'b0;
    rom[183] = 1'b0;
    rom[184] = 1'b0;
    rom[185] = 1'b0;
    rom[186] = 1'b0;
    rom[187] = 1'b0;
    rom[188] = 1'b0;
    rom[189] = 1'b0;
    rom[190] = 1'b0;
    rom[191] = 1'b0;
    rom[192] = 1'b0;
    rom[193] = 1'b0;
    rom[194] = 1'b0;
    rom[195] = 1'b0;
    rom[196] = 1'b0;
    rom[197] = 1'b0;
    rom[198] = 1'b0;
    rom[199] = 1'b0;
    rom[200] = 1'b0;
    rom[201] = 1'b0;
    rom[202] = 1'b0;
    rom[203] = 1'b0;
    rom[204] = 1'b0;
    rom[205] = 1'b0;
    rom[206] = 1'b0;
    rom[207] = 1'b0;
    rom[208] = 1'b0;
    rom[209] = 1'b0;
    rom[210] = 1'b0;
    rom[211] = 1'b0;
    rom[212] = 1'b0;
    rom[213] = 1'b0;
    rom[214] = 1'b0;
    rom[215] = 1'b0;
    rom[216] = 1'b0;
    rom[217] = 1'b0;
    rom[218] = 1'b0;
    rom[219] = 1'b0;
    rom[220] = 1'b0;
    rom[221] = 1'b0;
    rom[222] = 1'b0;
    rom[223] = 1'b0;
    rom[224] = 1'b0;
    rom[225] = 1'b0;
    rom[226] = 1'b0;
    rom[227] = 1'b0;
    rom[228] = 1'b0;
    rom[229] = 1'b0;
    rom[230] = 1'b0;
    rom[231] = 1'b0;
    rom[232] = 1'b0;
    rom[233] = 1'b0;
    rom[234] = 1'b0;
    rom[235] = 1'b0;
    rom[236] = 1'b0;
    rom[237] = 1'b0;
    rom[238] = 1'b0;
    rom[239] = 1'b0;
    rom[240] = 1'b0;
    rom[241] = 1'b0;
    rom[242] = 1'b0;
    rom[243] = 1'b0;
    rom[244] = 1'b0;
    rom[245] = 1'b0;
    rom[246] = 1'b0;
    rom[247] = 1'b0;
    rom[248] = 1'b0;
    rom[249] = 1'b0;
    rom[250] = 1'b0;
    rom[251] = 1'b0;
    rom[252] = 1'b0;
    rom[253] = 1'b0;
    rom[254] = 1'b0;
    rom[255] = 1'b0;
    rom[256] = 1'b0;
    rom[257] = 1'b0;
    rom[258] = 1'b0;
    rom[259] = 1'b0;
    rom[260] = 1'b0;
    rom[261] = 1'b0;
    rom[262] = 1'b0;
    rom[263] = 1'b0;
    rom[264] = 1'b0;
    rom[265] = 1'b0;
    rom[266] = 1'b0;
    rom[267] = 1'b0;
    rom[268] = 1'b0;
    rom[269] = 1'b0;
    rom[270] = 1'b0;
    rom[271] = 1'b0;
    rom[272] = 1'b0;
    rom[273] = 1'b0;
    rom[274] = 1'b0;
    rom[275] = 1'b0;
    rom[276] = 1'b0;
    rom[277] = 1'b0;
    rom[278] = 1'b0;
    rom[279] = 1'b0;
    rom[280] = 1'b0;
    rom[281] = 1'b0;
    rom[282] = 1'b0;
    rom[283] = 1'b0;
    rom[284] = 1'b0;
    rom[285] = 1'b0;
    rom[286] = 1'b0;
    rom[287] = 1'b0;
    rom[288] = 1'b0;
    rom[289] = 1'b0;
    rom[290] = 1'b0;
    rom[291] = 1'b0;
    rom[292] = 1'b0;
    rom[293] = 1'b0;
    rom[294] = 1'b0;
    rom[295] = 1'b0;
    rom[296] = 1'b0;
    rom[297] = 1'b0;
    rom[298] = 1'b0;
    rom[299] = 1'b0;
    rom[300] = 1'b0;
    rom[301] = 1'b0;
    rom[302] = 1'b0;
    rom[303] = 1'b0;
    rom[304] = 1'b0;
    rom[305] = 1'b0;
    rom[306] = 1'b0;
    rom[307] = 1'b0;
    rom[308] = 1'b0;
    rom[309] = 1'b0;
    rom[310] = 1'b0;
    rom[311] = 1'b0;
    rom[312] = 1'b0;
    rom[313] = 1'b0;
    rom[314] = 1'b0;
    rom[315] = 1'b0;
    rom[316] = 1'b0;
    rom[317] = 1'b0;
    rom[318] = 1'b0;
    rom[319] = 1'b0;
    rom[320] = 1'b0;
    rom[321] = 1'b0;
    rom[322] = 1'b0;
    rom[323] = 1'b0;
    rom[324] = 1'b0;
    rom[325] = 1'b0;
    rom[326] = 1'b0;
    rom[327] = 1'b0;
    rom[328] = 1'b0;
    rom[329] = 1'b0;
    rom[330] = 1'b0;
    rom[331] = 1'b0;
    rom[332] = 1'b0;
    rom[333] = 1'b0;
    rom[334] = 1'b0;
    rom[335] = 1'b0;
    rom[336] = 1'b0;
    rom[337] = 1'b0;
    rom[338] = 1'b0;
    rom[339] = 1'b0;
    rom[340] = 1'b0;
    rom[341] = 1'b0;
    rom[342] = 1'b0;
    rom[343] = 1'b0;
    rom[344] = 1'b0;
    rom[345] = 1'b0;
    rom[346] = 1'b0;
    rom[347] = 1'b0;
    rom[348] = 1'b0;
    rom[349] = 1'b0;
    rom[350] = 1'b0;
    rom[351] = 1'b0;
    rom[352] = 1'b0;
    rom[353] = 1'b0;
    rom[354] = 1'b0;
    rom[355] = 1'b0;
    rom[356] = 1'b0;
    rom[357] = 1'b0;
    rom[358] = 1'b0;
    rom[359] = 1'b0;
    rom[360] = 1'b0;
    rom[361] = 1'b0;
    rom[362] = 1'b0;
    rom[363] = 1'b0;
    rom[364] = 1'b0;
    rom[365] = 1'b0;
    rom[366] = 1'b0;
    rom[367] = 1'b0;
    rom[368] = 1'b0;
    rom[369] = 1'b0;
    rom[370] = 1'b0;
    rom[371] = 1'b0;
    rom[372] = 1'b0;
    rom[373] = 1'b0;
    rom[374] = 1'b0;
    rom[375] = 1'b0;
    rom[376] = 1'b0;
    rom[377] = 1'b0;
    rom[378] = 1'b0;
    rom[379] = 1'b0;
    rom[380] = 1'b0;
    rom[381] = 1'b0;
    rom[382] = 1'b0;
    rom[383] = 1'b0;
    rom[384] = 1'b0;
    rom[385] = 1'b0;
    rom[386] = 1'b0;
    rom[387] = 1'b0;
    rom[388] = 1'b0;
    rom[389] = 1'b0;
    rom[390] = 1'b0;
    rom[391] = 1'b0;
    rom[392] = 1'b0;
    rom[393] = 1'b0;
    rom[394] = 1'b0;
    rom[395] = 1'b0;
    rom[396] = 1'b0;
    rom[397] = 1'b0;
    rom[398] = 1'b0;
    rom[399] = 1'b0;
    rom[400] = 1'b0;
    rom[401] = 1'b0;
    rom[402] = 1'b0;
    rom[403] = 1'b0;
    rom[404] = 1'b0;
    rom[405] = 1'b0;
    rom[406] = 1'b0;
    rom[407] = 1'b0;
    rom[408] = 1'b0;
    rom[409] = 1'b0;
    rom[410] = 1'b0;
    rom[411] = 1'b0;
    rom[412] = 1'b0;
    rom[413] = 1'b0;
    rom[414] = 1'b0;
    rom[415] = 1'b0;
    rom[416] = 1'b0;
    rom[417] = 1'b0;
    rom[418] = 1'b0;
    rom[419] = 1'b0;
    rom[420] = 1'b0;
    rom[421] = 1'b0;
    rom[422] = 1'b0;
    rom[423] = 1'b0;
    rom[424] = 1'b0;
    rom[425] = 1'b0;
    rom[426] = 1'b0;
    rom[427] = 1'b0;
    rom[428] = 1'b0;
    rom[429] = 1'b0;
    rom[430] = 1'b0;
    rom[431] = 1'b0;
    rom[432] = 1'b0;
    rom[433] = 1'b0;
    rom[434] = 1'b0;
    rom[435] = 1'b0;
    rom[436] = 1'b0;
    rom[437] = 1'b0;
    rom[438] = 1'b0;
    rom[439] = 1'b0;
    rom[440] = 1'b0;
    rom[441] = 1'b0;
    rom[442] = 1'b0;
    rom[443] = 1'b0;
    rom[444] = 1'b0;
    rom[445] = 1'b0;
    rom[446] = 1'b0;
    rom[447] = 1'b0;
    rom[448] = 1'b0;
    rom[449] = 1'b0;
    rom[450] = 1'b0;
    rom[451] = 1'b0;
    rom[452] = 1'b0;
    rom[453] = 1'b0;
    rom[454] = 1'b0;
    rom[455] = 1'b0;
    rom[456] = 1'b0;
    rom[457] = 1'b0;
    rom[458] = 1'b0;
    rom[459] = 1'b0;
    rom[460] = 1'b0;
    rom[461] = 1'b0;
    rom[462] = 1'b0;
    rom[463] = 1'b0;
    rom[464] = 1'b0;
    rom[465] = 1'b0;
    rom[466] = 1'b0;
    rom[467] = 1'b0;
    rom[468] = 1'b0;
    rom[469] = 1'b0;
    rom[470] = 1'b0;
    rom[471] = 1'b0;
    rom[472] = 1'b0;
    rom[473] = 1'b0;
    rom[474] = 1'b0;
    rom[475] = 1'b0;
    rom[476] = 1'b0;
    rom[477] = 1'b0;
    rom[478] = 1'b0;
    rom[479] = 1'b0;
    rom[480] = 1'b0;
    rom[481] = 1'b0;
    rom[482] = 1'b0;
    rom[483] = 1'b0;
    rom[484] = 1'b0;
    rom[485] = 1'b0;
    rom[486] = 1'b0;
    rom[487] = 1'b0;
    rom[488] = 1'b0;
    rom[489] = 1'b0;
    rom[490] = 1'b0;
    rom[491] = 1'b0;
    rom[492] = 1'b0;
    rom[493] = 1'b0;
    rom[494] = 1'b0;
    rom[495] = 1'b0;
    rom[496] = 1'b0;
    rom[497] = 1'b0;
    rom[498] = 1'b0;
    rom[499] = 1'b0;
    rom[500] = 1'b0;
    rom[501] = 1'b0;
    rom[502] = 1'b0;
    rom[503] = 1'b0;
    rom[504] = 1'b0;
    rom[505] = 1'b0;
    rom[506] = 1'b0;
    rom[507] = 1'b0;
    rom[508] = 1'b0;
    rom[509] = 1'b0;
    rom[510] = 1'b0;
    rom[511] = 1'b0;
end


always @(posedge clk)
begin
    addra_d <= addra;
    rom_pipea <= rom[addra_d];
    doa_d <= rom_pipea;
end
endmodule
