/*************************************************************************/
//// File        : pipe_mux_512_1.v
// Description : Implements a pipelined multiplexer to be used in high speed design
// This module has a delay of 4 clock cycles//
// -------------------------------------------------------------------
//
/***************************************************************************/


module pipe_mux_512_1
(
    input clk,
    input sync_reset,
    input valid_i,
    input [8:0] sel,
    input [511:0] input_word,
    output valid_o,
    output [8:0] sel_o,
    output output_word
);

(* KEEP = "TRUE" *) reg [8:0] sel_d0_0;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_1;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_2;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_3;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_4;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_5;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_6;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_7;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_8;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_9;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_10;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_11;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_12;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_13;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_14;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_15;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_16;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_17;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_18;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_19;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_20;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_21;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_22;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_23;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_24;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_25;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_26;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_27;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_28;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_29;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_30;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_31;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_32;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_33;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_34;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_35;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_36;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_37;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_38;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_39;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_40;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_41;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_42;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_43;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_44;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_45;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_46;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_47;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_48;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_49;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_50;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_51;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_52;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_53;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_54;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_55;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_56;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_57;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_58;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_59;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_60;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_61;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_62;
(* KEEP = "TRUE" *) reg [8:0] sel_d0_63;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_0;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_1;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_2;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_3;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_4;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_5;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_6;
(* KEEP = "TRUE" *) reg [8:0] sel_d1_7;
(* KEEP = "TRUE" *) reg [8:0] sel_d2_0;
(* KEEP = "TRUE" *) reg [8:0] sel_d3;
reg valid_d0;
reg valid_d1;
reg valid_d2;
reg valid_d3;
reg [0:0] mux_d0_0, next_mux_d0_0;
reg [0:0] mux_d0_1, next_mux_d0_1;
reg [0:0] mux_d0_2, next_mux_d0_2;
reg [0:0] mux_d0_3, next_mux_d0_3;
reg [0:0] mux_d0_4, next_mux_d0_4;
reg [0:0] mux_d0_5, next_mux_d0_5;
reg [0:0] mux_d0_6, next_mux_d0_6;
reg [0:0] mux_d0_7, next_mux_d0_7;
reg [0:0] mux_d0_8, next_mux_d0_8;
reg [0:0] mux_d0_9, next_mux_d0_9;
reg [0:0] mux_d0_10, next_mux_d0_10;
reg [0:0] mux_d0_11, next_mux_d0_11;
reg [0:0] mux_d0_12, next_mux_d0_12;
reg [0:0] mux_d0_13, next_mux_d0_13;
reg [0:0] mux_d0_14, next_mux_d0_14;
reg [0:0] mux_d0_15, next_mux_d0_15;
reg [0:0] mux_d0_16, next_mux_d0_16;
reg [0:0] mux_d0_17, next_mux_d0_17;
reg [0:0] mux_d0_18, next_mux_d0_18;
reg [0:0] mux_d0_19, next_mux_d0_19;
reg [0:0] mux_d0_20, next_mux_d0_20;
reg [0:0] mux_d0_21, next_mux_d0_21;
reg [0:0] mux_d0_22, next_mux_d0_22;
reg [0:0] mux_d0_23, next_mux_d0_23;
reg [0:0] mux_d0_24, next_mux_d0_24;
reg [0:0] mux_d0_25, next_mux_d0_25;
reg [0:0] mux_d0_26, next_mux_d0_26;
reg [0:0] mux_d0_27, next_mux_d0_27;
reg [0:0] mux_d0_28, next_mux_d0_28;
reg [0:0] mux_d0_29, next_mux_d0_29;
reg [0:0] mux_d0_30, next_mux_d0_30;
reg [0:0] mux_d0_31, next_mux_d0_31;
reg [0:0] mux_d0_32, next_mux_d0_32;
reg [0:0] mux_d0_33, next_mux_d0_33;
reg [0:0] mux_d0_34, next_mux_d0_34;
reg [0:0] mux_d0_35, next_mux_d0_35;
reg [0:0] mux_d0_36, next_mux_d0_36;
reg [0:0] mux_d0_37, next_mux_d0_37;
reg [0:0] mux_d0_38, next_mux_d0_38;
reg [0:0] mux_d0_39, next_mux_d0_39;
reg [0:0] mux_d0_40, next_mux_d0_40;
reg [0:0] mux_d0_41, next_mux_d0_41;
reg [0:0] mux_d0_42, next_mux_d0_42;
reg [0:0] mux_d0_43, next_mux_d0_43;
reg [0:0] mux_d0_44, next_mux_d0_44;
reg [0:0] mux_d0_45, next_mux_d0_45;
reg [0:0] mux_d0_46, next_mux_d0_46;
reg [0:0] mux_d0_47, next_mux_d0_47;
reg [0:0] mux_d0_48, next_mux_d0_48;
reg [0:0] mux_d0_49, next_mux_d0_49;
reg [0:0] mux_d0_50, next_mux_d0_50;
reg [0:0] mux_d0_51, next_mux_d0_51;
reg [0:0] mux_d0_52, next_mux_d0_52;
reg [0:0] mux_d0_53, next_mux_d0_53;
reg [0:0] mux_d0_54, next_mux_d0_54;
reg [0:0] mux_d0_55, next_mux_d0_55;
reg [0:0] mux_d0_56, next_mux_d0_56;
reg [0:0] mux_d0_57, next_mux_d0_57;
reg [0:0] mux_d0_58, next_mux_d0_58;
reg [0:0] mux_d0_59, next_mux_d0_59;
reg [0:0] mux_d0_60, next_mux_d0_60;
reg [0:0] mux_d0_61, next_mux_d0_61;
reg [0:0] mux_d0_62, next_mux_d0_62;
reg [0:0] mux_d0_63, next_mux_d0_63;
reg [0:0] mux_d1_0, next_mux_d1_0;
reg [0:0] mux_d1_1, next_mux_d1_1;
reg [0:0] mux_d1_2, next_mux_d1_2;
reg [0:0] mux_d1_3, next_mux_d1_3;
reg [0:0] mux_d1_4, next_mux_d1_4;
reg [0:0] mux_d1_5, next_mux_d1_5;
reg [0:0] mux_d1_6, next_mux_d1_6;
reg [0:0] mux_d1_7, next_mux_d1_7;
reg [0:0] mux_d2_0, next_mux_d2_0;
reg [511:0] input_word_d;

assign output_word = mux_d2_0;
assign valid_o = valid_d3;
assign sel_o = sel_d3;

always @(posedge clk) begin
    if (sync_reset) begin
        valid_d0  <= 0;
        valid_d1  <= 0;
        valid_d2  <= 0;
        valid_d3  <= 0;
    end else begin
        valid_d0  <= valid_i;
        valid_d1  <= valid_d0;
        valid_d2  <= valid_d1;
        valid_d3  <= valid_d2;
    end
end


always @(posedge clk) begin
    input_word_d <= input_word;
    mux_d0_0 <= next_mux_d0_0;
    mux_d0_1 <= next_mux_d0_1;
    mux_d0_2 <= next_mux_d0_2;
    mux_d0_3 <= next_mux_d0_3;
    mux_d0_4 <= next_mux_d0_4;
    mux_d0_5 <= next_mux_d0_5;
    mux_d0_6 <= next_mux_d0_6;
    mux_d0_7 <= next_mux_d0_7;
    mux_d0_8 <= next_mux_d0_8;
    mux_d0_9 <= next_mux_d0_9;
    mux_d0_10 <= next_mux_d0_10;
    mux_d0_11 <= next_mux_d0_11;
    mux_d0_12 <= next_mux_d0_12;
    mux_d0_13 <= next_mux_d0_13;
    mux_d0_14 <= next_mux_d0_14;
    mux_d0_15 <= next_mux_d0_15;
    mux_d0_16 <= next_mux_d0_16;
    mux_d0_17 <= next_mux_d0_17;
    mux_d0_18 <= next_mux_d0_18;
    mux_d0_19 <= next_mux_d0_19;
    mux_d0_20 <= next_mux_d0_20;
    mux_d0_21 <= next_mux_d0_21;
    mux_d0_22 <= next_mux_d0_22;
    mux_d0_23 <= next_mux_d0_23;
    mux_d0_24 <= next_mux_d0_24;
    mux_d0_25 <= next_mux_d0_25;
    mux_d0_26 <= next_mux_d0_26;
    mux_d0_27 <= next_mux_d0_27;
    mux_d0_28 <= next_mux_d0_28;
    mux_d0_29 <= next_mux_d0_29;
    mux_d0_30 <= next_mux_d0_30;
    mux_d0_31 <= next_mux_d0_31;
    mux_d0_32 <= next_mux_d0_32;
    mux_d0_33 <= next_mux_d0_33;
    mux_d0_34 <= next_mux_d0_34;
    mux_d0_35 <= next_mux_d0_35;
    mux_d0_36 <= next_mux_d0_36;
    mux_d0_37 <= next_mux_d0_37;
    mux_d0_38 <= next_mux_d0_38;
    mux_d0_39 <= next_mux_d0_39;
    mux_d0_40 <= next_mux_d0_40;
    mux_d0_41 <= next_mux_d0_41;
    mux_d0_42 <= next_mux_d0_42;
    mux_d0_43 <= next_mux_d0_43;
    mux_d0_44 <= next_mux_d0_44;
    mux_d0_45 <= next_mux_d0_45;
    mux_d0_46 <= next_mux_d0_46;
    mux_d0_47 <= next_mux_d0_47;
    mux_d0_48 <= next_mux_d0_48;
    mux_d0_49 <= next_mux_d0_49;
    mux_d0_50 <= next_mux_d0_50;
    mux_d0_51 <= next_mux_d0_51;
    mux_d0_52 <= next_mux_d0_52;
    mux_d0_53 <= next_mux_d0_53;
    mux_d0_54 <= next_mux_d0_54;
    mux_d0_55 <= next_mux_d0_55;
    mux_d0_56 <= next_mux_d0_56;
    mux_d0_57 <= next_mux_d0_57;
    mux_d0_58 <= next_mux_d0_58;
    mux_d0_59 <= next_mux_d0_59;
    mux_d0_60 <= next_mux_d0_60;
    mux_d0_61 <= next_mux_d0_61;
    mux_d0_62 <= next_mux_d0_62;
    mux_d0_63 <= next_mux_d0_63;
    mux_d1_0 <= next_mux_d1_0;
    mux_d1_1 <= next_mux_d1_1;
    mux_d1_2 <= next_mux_d1_2;
    mux_d1_3 <= next_mux_d1_3;
    mux_d1_4 <= next_mux_d1_4;
    mux_d1_5 <= next_mux_d1_5;
    mux_d1_6 <= next_mux_d1_6;
    mux_d1_7 <= next_mux_d1_7;
    mux_d2_0 <= next_mux_d2_0;
    sel_d0_0 <= sel;
    sel_d0_1 <= sel;
    sel_d0_2 <= sel;
    sel_d0_3 <= sel;
    sel_d0_4 <= sel;
    sel_d0_5 <= sel;
    sel_d0_6 <= sel;
    sel_d0_7 <= sel;
    sel_d0_8 <= sel;
    sel_d0_9 <= sel;
    sel_d0_10 <= sel;
    sel_d0_11 <= sel;
    sel_d0_12 <= sel;
    sel_d0_13 <= sel;
    sel_d0_14 <= sel;
    sel_d0_15 <= sel;
    sel_d0_16 <= sel;
    sel_d0_17 <= sel;
    sel_d0_18 <= sel;
    sel_d0_19 <= sel;
    sel_d0_20 <= sel;
    sel_d0_21 <= sel;
    sel_d0_22 <= sel;
    sel_d0_23 <= sel;
    sel_d0_24 <= sel;
    sel_d0_25 <= sel;
    sel_d0_26 <= sel;
    sel_d0_27 <= sel;
    sel_d0_28 <= sel;
    sel_d0_29 <= sel;
    sel_d0_30 <= sel;
    sel_d0_31 <= sel;
    sel_d0_32 <= sel;
    sel_d0_33 <= sel;
    sel_d0_34 <= sel;
    sel_d0_35 <= sel;
    sel_d0_36 <= sel;
    sel_d0_37 <= sel;
    sel_d0_38 <= sel;
    sel_d0_39 <= sel;
    sel_d0_40 <= sel;
    sel_d0_41 <= sel;
    sel_d0_42 <= sel;
    sel_d0_43 <= sel;
    sel_d0_44 <= sel;
    sel_d0_45 <= sel;
    sel_d0_46 <= sel;
    sel_d0_47 <= sel;
    sel_d0_48 <= sel;
    sel_d0_49 <= sel;
    sel_d0_50 <= sel;
    sel_d0_51 <= sel;
    sel_d0_52 <= sel;
    sel_d0_53 <= sel;
    sel_d0_54 <= sel;
    sel_d0_55 <= sel;
    sel_d0_56 <= sel;
    sel_d0_57 <= sel;
    sel_d0_58 <= sel;
    sel_d0_59 <= sel;
    sel_d0_60 <= sel;
    sel_d0_61 <= sel;
    sel_d0_62 <= sel;
    sel_d0_63 <= sel;
    sel_d1_0 <= sel_d0_63;
    sel_d1_1 <= sel_d0_63;
    sel_d1_2 <= sel_d0_63;
    sel_d1_3 <= sel_d0_63;
    sel_d1_4 <= sel_d0_63;
    sel_d1_5 <= sel_d0_63;
    sel_d1_6 <= sel_d0_63;
    sel_d1_7 <= sel_d0_63;
    sel_d2_0 <= sel_d1_7;
    sel_d3 <= sel_d2_0;
end


always @*
begin
    next_mux_d0_0 = mux_d0_0;
    next_mux_d0_1 = mux_d0_1;
    next_mux_d0_2 = mux_d0_2;
    next_mux_d0_3 = mux_d0_3;
    next_mux_d0_4 = mux_d0_4;
    next_mux_d0_5 = mux_d0_5;
    next_mux_d0_6 = mux_d0_6;
    next_mux_d0_7 = mux_d0_7;
    next_mux_d0_8 = mux_d0_8;
    next_mux_d0_9 = mux_d0_9;
    next_mux_d0_10 = mux_d0_10;
    next_mux_d0_11 = mux_d0_11;
    next_mux_d0_12 = mux_d0_12;
    next_mux_d0_13 = mux_d0_13;
    next_mux_d0_14 = mux_d0_14;
    next_mux_d0_15 = mux_d0_15;
    next_mux_d0_16 = mux_d0_16;
    next_mux_d0_17 = mux_d0_17;
    next_mux_d0_18 = mux_d0_18;
    next_mux_d0_19 = mux_d0_19;
    next_mux_d0_20 = mux_d0_20;
    next_mux_d0_21 = mux_d0_21;
    next_mux_d0_22 = mux_d0_22;
    next_mux_d0_23 = mux_d0_23;
    next_mux_d0_24 = mux_d0_24;
    next_mux_d0_25 = mux_d0_25;
    next_mux_d0_26 = mux_d0_26;
    next_mux_d0_27 = mux_d0_27;
    next_mux_d0_28 = mux_d0_28;
    next_mux_d0_29 = mux_d0_29;
    next_mux_d0_30 = mux_d0_30;
    next_mux_d0_31 = mux_d0_31;
    next_mux_d0_32 = mux_d0_32;
    next_mux_d0_33 = mux_d0_33;
    next_mux_d0_34 = mux_d0_34;
    next_mux_d0_35 = mux_d0_35;
    next_mux_d0_36 = mux_d0_36;
    next_mux_d0_37 = mux_d0_37;
    next_mux_d0_38 = mux_d0_38;
    next_mux_d0_39 = mux_d0_39;
    next_mux_d0_40 = mux_d0_40;
    next_mux_d0_41 = mux_d0_41;
    next_mux_d0_42 = mux_d0_42;
    next_mux_d0_43 = mux_d0_43;
    next_mux_d0_44 = mux_d0_44;
    next_mux_d0_45 = mux_d0_45;
    next_mux_d0_46 = mux_d0_46;
    next_mux_d0_47 = mux_d0_47;
    next_mux_d0_48 = mux_d0_48;
    next_mux_d0_49 = mux_d0_49;
    next_mux_d0_50 = mux_d0_50;
    next_mux_d0_51 = mux_d0_51;
    next_mux_d0_52 = mux_d0_52;
    next_mux_d0_53 = mux_d0_53;
    next_mux_d0_54 = mux_d0_54;
    next_mux_d0_55 = mux_d0_55;
    next_mux_d0_56 = mux_d0_56;
    next_mux_d0_57 = mux_d0_57;
    next_mux_d0_58 = mux_d0_58;
    next_mux_d0_59 = mux_d0_59;
    next_mux_d0_60 = mux_d0_60;
    next_mux_d0_61 = mux_d0_61;
    next_mux_d0_62 = mux_d0_62;
    next_mux_d0_63 = mux_d0_63;
    next_mux_d1_0 = mux_d1_0;
    next_mux_d1_1 = mux_d1_1;
    next_mux_d1_2 = mux_d1_2;
    next_mux_d1_3 = mux_d1_3;
    next_mux_d1_4 = mux_d1_4;
    next_mux_d1_5 = mux_d1_5;
    next_mux_d1_6 = mux_d1_6;
    next_mux_d1_7 = mux_d1_7;
    next_mux_d2_0 = mux_d2_0;

    if (sel_d0_0[2:0] == 0) begin
        next_mux_d0_0 = input_word_d[0];
    end else if (sel_d0_0[2:0] == 1) begin
        next_mux_d0_0 = input_word_d[1];
    end else if (sel_d0_0[2:0] == 2) begin
        next_mux_d0_0 = input_word_d[2];
    end else if (sel_d0_0[2:0] == 3) begin
        next_mux_d0_0 = input_word_d[3];
    end else if (sel_d0_0[2:0] == 4) begin
        next_mux_d0_0 = input_word_d[4];
    end else if (sel_d0_0[2:0] == 5) begin
        next_mux_d0_0 = input_word_d[5];
    end else if (sel_d0_0[2:0] == 6) begin
        next_mux_d0_0 = input_word_d[6];
    end else begin
        next_mux_d0_0 = input_word_d[7];
    end

    if (sel_d0_1[2:0] == 0) begin
        next_mux_d0_1 = input_word_d[8];
    end else if (sel_d0_1[2:0] == 1) begin
        next_mux_d0_1 = input_word_d[9];
    end else if (sel_d0_1[2:0] == 2) begin
        next_mux_d0_1 = input_word_d[10];
    end else if (sel_d0_1[2:0] == 3) begin
        next_mux_d0_1 = input_word_d[11];
    end else if (sel_d0_1[2:0] == 4) begin
        next_mux_d0_1 = input_word_d[12];
    end else if (sel_d0_1[2:0] == 5) begin
        next_mux_d0_1 = input_word_d[13];
    end else if (sel_d0_1[2:0] == 6) begin
        next_mux_d0_1 = input_word_d[14];
    end else begin
        next_mux_d0_1 = input_word_d[15];
    end

    if (sel_d0_2[2:0] == 0) begin
        next_mux_d0_2 = input_word_d[16];
    end else if (sel_d0_2[2:0] == 1) begin
        next_mux_d0_2 = input_word_d[17];
    end else if (sel_d0_2[2:0] == 2) begin
        next_mux_d0_2 = input_word_d[18];
    end else if (sel_d0_2[2:0] == 3) begin
        next_mux_d0_2 = input_word_d[19];
    end else if (sel_d0_2[2:0] == 4) begin
        next_mux_d0_2 = input_word_d[20];
    end else if (sel_d0_2[2:0] == 5) begin
        next_mux_d0_2 = input_word_d[21];
    end else if (sel_d0_2[2:0] == 6) begin
        next_mux_d0_2 = input_word_d[22];
    end else begin
        next_mux_d0_2 = input_word_d[23];
    end

    if (sel_d0_3[2:0] == 0) begin
        next_mux_d0_3 = input_word_d[24];
    end else if (sel_d0_3[2:0] == 1) begin
        next_mux_d0_3 = input_word_d[25];
    end else if (sel_d0_3[2:0] == 2) begin
        next_mux_d0_3 = input_word_d[26];
    end else if (sel_d0_3[2:0] == 3) begin
        next_mux_d0_3 = input_word_d[27];
    end else if (sel_d0_3[2:0] == 4) begin
        next_mux_d0_3 = input_word_d[28];
    end else if (sel_d0_3[2:0] == 5) begin
        next_mux_d0_3 = input_word_d[29];
    end else if (sel_d0_3[2:0] == 6) begin
        next_mux_d0_3 = input_word_d[30];
    end else begin
        next_mux_d0_3 = input_word_d[31];
    end

    if (sel_d0_4[2:0] == 0) begin
        next_mux_d0_4 = input_word_d[32];
    end else if (sel_d0_4[2:0] == 1) begin
        next_mux_d0_4 = input_word_d[33];
    end else if (sel_d0_4[2:0] == 2) begin
        next_mux_d0_4 = input_word_d[34];
    end else if (sel_d0_4[2:0] == 3) begin
        next_mux_d0_4 = input_word_d[35];
    end else if (sel_d0_4[2:0] == 4) begin
        next_mux_d0_4 = input_word_d[36];
    end else if (sel_d0_4[2:0] == 5) begin
        next_mux_d0_4 = input_word_d[37];
    end else if (sel_d0_4[2:0] == 6) begin
        next_mux_d0_4 = input_word_d[38];
    end else begin
        next_mux_d0_4 = input_word_d[39];
    end

    if (sel_d0_5[2:0] == 0) begin
        next_mux_d0_5 = input_word_d[40];
    end else if (sel_d0_5[2:0] == 1) begin
        next_mux_d0_5 = input_word_d[41];
    end else if (sel_d0_5[2:0] == 2) begin
        next_mux_d0_5 = input_word_d[42];
    end else if (sel_d0_5[2:0] == 3) begin
        next_mux_d0_5 = input_word_d[43];
    end else if (sel_d0_5[2:0] == 4) begin
        next_mux_d0_5 = input_word_d[44];
    end else if (sel_d0_5[2:0] == 5) begin
        next_mux_d0_5 = input_word_d[45];
    end else if (sel_d0_5[2:0] == 6) begin
        next_mux_d0_5 = input_word_d[46];
    end else begin
        next_mux_d0_5 = input_word_d[47];
    end

    if (sel_d0_6[2:0] == 0) begin
        next_mux_d0_6 = input_word_d[48];
    end else if (sel_d0_6[2:0] == 1) begin
        next_mux_d0_6 = input_word_d[49];
    end else if (sel_d0_6[2:0] == 2) begin
        next_mux_d0_6 = input_word_d[50];
    end else if (sel_d0_6[2:0] == 3) begin
        next_mux_d0_6 = input_word_d[51];
    end else if (sel_d0_6[2:0] == 4) begin
        next_mux_d0_6 = input_word_d[52];
    end else if (sel_d0_6[2:0] == 5) begin
        next_mux_d0_6 = input_word_d[53];
    end else if (sel_d0_6[2:0] == 6) begin
        next_mux_d0_6 = input_word_d[54];
    end else begin
        next_mux_d0_6 = input_word_d[55];
    end

    if (sel_d0_7[2:0] == 0) begin
        next_mux_d0_7 = input_word_d[56];
    end else if (sel_d0_7[2:0] == 1) begin
        next_mux_d0_7 = input_word_d[57];
    end else if (sel_d0_7[2:0] == 2) begin
        next_mux_d0_7 = input_word_d[58];
    end else if (sel_d0_7[2:0] == 3) begin
        next_mux_d0_7 = input_word_d[59];
    end else if (sel_d0_7[2:0] == 4) begin
        next_mux_d0_7 = input_word_d[60];
    end else if (sel_d0_7[2:0] == 5) begin
        next_mux_d0_7 = input_word_d[61];
    end else if (sel_d0_7[2:0] == 6) begin
        next_mux_d0_7 = input_word_d[62];
    end else begin
        next_mux_d0_7 = input_word_d[63];
    end

    if (sel_d0_8[2:0] == 0) begin
        next_mux_d0_8 = input_word_d[64];
    end else if (sel_d0_8[2:0] == 1) begin
        next_mux_d0_8 = input_word_d[65];
    end else if (sel_d0_8[2:0] == 2) begin
        next_mux_d0_8 = input_word_d[66];
    end else if (sel_d0_8[2:0] == 3) begin
        next_mux_d0_8 = input_word_d[67];
    end else if (sel_d0_8[2:0] == 4) begin
        next_mux_d0_8 = input_word_d[68];
    end else if (sel_d0_8[2:0] == 5) begin
        next_mux_d0_8 = input_word_d[69];
    end else if (sel_d0_8[2:0] == 6) begin
        next_mux_d0_8 = input_word_d[70];
    end else begin
        next_mux_d0_8 = input_word_d[71];
    end

    if (sel_d0_9[2:0] == 0) begin
        next_mux_d0_9 = input_word_d[72];
    end else if (sel_d0_9[2:0] == 1) begin
        next_mux_d0_9 = input_word_d[73];
    end else if (sel_d0_9[2:0] == 2) begin
        next_mux_d0_9 = input_word_d[74];
    end else if (sel_d0_9[2:0] == 3) begin
        next_mux_d0_9 = input_word_d[75];
    end else if (sel_d0_9[2:0] == 4) begin
        next_mux_d0_9 = input_word_d[76];
    end else if (sel_d0_9[2:0] == 5) begin
        next_mux_d0_9 = input_word_d[77];
    end else if (sel_d0_9[2:0] == 6) begin
        next_mux_d0_9 = input_word_d[78];
    end else begin
        next_mux_d0_9 = input_word_d[79];
    end

    if (sel_d0_10[2:0] == 0) begin
        next_mux_d0_10 = input_word_d[80];
    end else if (sel_d0_10[2:0] == 1) begin
        next_mux_d0_10 = input_word_d[81];
    end else if (sel_d0_10[2:0] == 2) begin
        next_mux_d0_10 = input_word_d[82];
    end else if (sel_d0_10[2:0] == 3) begin
        next_mux_d0_10 = input_word_d[83];
    end else if (sel_d0_10[2:0] == 4) begin
        next_mux_d0_10 = input_word_d[84];
    end else if (sel_d0_10[2:0] == 5) begin
        next_mux_d0_10 = input_word_d[85];
    end else if (sel_d0_10[2:0] == 6) begin
        next_mux_d0_10 = input_word_d[86];
    end else begin
        next_mux_d0_10 = input_word_d[87];
    end

    if (sel_d0_11[2:0] == 0) begin
        next_mux_d0_11 = input_word_d[88];
    end else if (sel_d0_11[2:0] == 1) begin
        next_mux_d0_11 = input_word_d[89];
    end else if (sel_d0_11[2:0] == 2) begin
        next_mux_d0_11 = input_word_d[90];
    end else if (sel_d0_11[2:0] == 3) begin
        next_mux_d0_11 = input_word_d[91];
    end else if (sel_d0_11[2:0] == 4) begin
        next_mux_d0_11 = input_word_d[92];
    end else if (sel_d0_11[2:0] == 5) begin
        next_mux_d0_11 = input_word_d[93];
    end else if (sel_d0_11[2:0] == 6) begin
        next_mux_d0_11 = input_word_d[94];
    end else begin
        next_mux_d0_11 = input_word_d[95];
    end

    if (sel_d0_12[2:0] == 0) begin
        next_mux_d0_12 = input_word_d[96];
    end else if (sel_d0_12[2:0] == 1) begin
        next_mux_d0_12 = input_word_d[97];
    end else if (sel_d0_12[2:0] == 2) begin
        next_mux_d0_12 = input_word_d[98];
    end else if (sel_d0_12[2:0] == 3) begin
        next_mux_d0_12 = input_word_d[99];
    end else if (sel_d0_12[2:0] == 4) begin
        next_mux_d0_12 = input_word_d[100];
    end else if (sel_d0_12[2:0] == 5) begin
        next_mux_d0_12 = input_word_d[101];
    end else if (sel_d0_12[2:0] == 6) begin
        next_mux_d0_12 = input_word_d[102];
    end else begin
        next_mux_d0_12 = input_word_d[103];
    end

    if (sel_d0_13[2:0] == 0) begin
        next_mux_d0_13 = input_word_d[104];
    end else if (sel_d0_13[2:0] == 1) begin
        next_mux_d0_13 = input_word_d[105];
    end else if (sel_d0_13[2:0] == 2) begin
        next_mux_d0_13 = input_word_d[106];
    end else if (sel_d0_13[2:0] == 3) begin
        next_mux_d0_13 = input_word_d[107];
    end else if (sel_d0_13[2:0] == 4) begin
        next_mux_d0_13 = input_word_d[108];
    end else if (sel_d0_13[2:0] == 5) begin
        next_mux_d0_13 = input_word_d[109];
    end else if (sel_d0_13[2:0] == 6) begin
        next_mux_d0_13 = input_word_d[110];
    end else begin
        next_mux_d0_13 = input_word_d[111];
    end

    if (sel_d0_14[2:0] == 0) begin
        next_mux_d0_14 = input_word_d[112];
    end else if (sel_d0_14[2:0] == 1) begin
        next_mux_d0_14 = input_word_d[113];
    end else if (sel_d0_14[2:0] == 2) begin
        next_mux_d0_14 = input_word_d[114];
    end else if (sel_d0_14[2:0] == 3) begin
        next_mux_d0_14 = input_word_d[115];
    end else if (sel_d0_14[2:0] == 4) begin
        next_mux_d0_14 = input_word_d[116];
    end else if (sel_d0_14[2:0] == 5) begin
        next_mux_d0_14 = input_word_d[117];
    end else if (sel_d0_14[2:0] == 6) begin
        next_mux_d0_14 = input_word_d[118];
    end else begin
        next_mux_d0_14 = input_word_d[119];
    end

    if (sel_d0_15[2:0] == 0) begin
        next_mux_d0_15 = input_word_d[120];
    end else if (sel_d0_15[2:0] == 1) begin
        next_mux_d0_15 = input_word_d[121];
    end else if (sel_d0_15[2:0] == 2) begin
        next_mux_d0_15 = input_word_d[122];
    end else if (sel_d0_15[2:0] == 3) begin
        next_mux_d0_15 = input_word_d[123];
    end else if (sel_d0_15[2:0] == 4) begin
        next_mux_d0_15 = input_word_d[124];
    end else if (sel_d0_15[2:0] == 5) begin
        next_mux_d0_15 = input_word_d[125];
    end else if (sel_d0_15[2:0] == 6) begin
        next_mux_d0_15 = input_word_d[126];
    end else begin
        next_mux_d0_15 = input_word_d[127];
    end

    if (sel_d0_16[2:0] == 0) begin
        next_mux_d0_16 = input_word_d[128];
    end else if (sel_d0_16[2:0] == 1) begin
        next_mux_d0_16 = input_word_d[129];
    end else if (sel_d0_16[2:0] == 2) begin
        next_mux_d0_16 = input_word_d[130];
    end else if (sel_d0_16[2:0] == 3) begin
        next_mux_d0_16 = input_word_d[131];
    end else if (sel_d0_16[2:0] == 4) begin
        next_mux_d0_16 = input_word_d[132];
    end else if (sel_d0_16[2:0] == 5) begin
        next_mux_d0_16 = input_word_d[133];
    end else if (sel_d0_16[2:0] == 6) begin
        next_mux_d0_16 = input_word_d[134];
    end else begin
        next_mux_d0_16 = input_word_d[135];
    end

    if (sel_d0_17[2:0] == 0) begin
        next_mux_d0_17 = input_word_d[136];
    end else if (sel_d0_17[2:0] == 1) begin
        next_mux_d0_17 = input_word_d[137];
    end else if (sel_d0_17[2:0] == 2) begin
        next_mux_d0_17 = input_word_d[138];
    end else if (sel_d0_17[2:0] == 3) begin
        next_mux_d0_17 = input_word_d[139];
    end else if (sel_d0_17[2:0] == 4) begin
        next_mux_d0_17 = input_word_d[140];
    end else if (sel_d0_17[2:0] == 5) begin
        next_mux_d0_17 = input_word_d[141];
    end else if (sel_d0_17[2:0] == 6) begin
        next_mux_d0_17 = input_word_d[142];
    end else begin
        next_mux_d0_17 = input_word_d[143];
    end

    if (sel_d0_18[2:0] == 0) begin
        next_mux_d0_18 = input_word_d[144];
    end else if (sel_d0_18[2:0] == 1) begin
        next_mux_d0_18 = input_word_d[145];
    end else if (sel_d0_18[2:0] == 2) begin
        next_mux_d0_18 = input_word_d[146];
    end else if (sel_d0_18[2:0] == 3) begin
        next_mux_d0_18 = input_word_d[147];
    end else if (sel_d0_18[2:0] == 4) begin
        next_mux_d0_18 = input_word_d[148];
    end else if (sel_d0_18[2:0] == 5) begin
        next_mux_d0_18 = input_word_d[149];
    end else if (sel_d0_18[2:0] == 6) begin
        next_mux_d0_18 = input_word_d[150];
    end else begin
        next_mux_d0_18 = input_word_d[151];
    end

    if (sel_d0_19[2:0] == 0) begin
        next_mux_d0_19 = input_word_d[152];
    end else if (sel_d0_19[2:0] == 1) begin
        next_mux_d0_19 = input_word_d[153];
    end else if (sel_d0_19[2:0] == 2) begin
        next_mux_d0_19 = input_word_d[154];
    end else if (sel_d0_19[2:0] == 3) begin
        next_mux_d0_19 = input_word_d[155];
    end else if (sel_d0_19[2:0] == 4) begin
        next_mux_d0_19 = input_word_d[156];
    end else if (sel_d0_19[2:0] == 5) begin
        next_mux_d0_19 = input_word_d[157];
    end else if (sel_d0_19[2:0] == 6) begin
        next_mux_d0_19 = input_word_d[158];
    end else begin
        next_mux_d0_19 = input_word_d[159];
    end

    if (sel_d0_20[2:0] == 0) begin
        next_mux_d0_20 = input_word_d[160];
    end else if (sel_d0_20[2:0] == 1) begin
        next_mux_d0_20 = input_word_d[161];
    end else if (sel_d0_20[2:0] == 2) begin
        next_mux_d0_20 = input_word_d[162];
    end else if (sel_d0_20[2:0] == 3) begin
        next_mux_d0_20 = input_word_d[163];
    end else if (sel_d0_20[2:0] == 4) begin
        next_mux_d0_20 = input_word_d[164];
    end else if (sel_d0_20[2:0] == 5) begin
        next_mux_d0_20 = input_word_d[165];
    end else if (sel_d0_20[2:0] == 6) begin
        next_mux_d0_20 = input_word_d[166];
    end else begin
        next_mux_d0_20 = input_word_d[167];
    end

    if (sel_d0_21[2:0] == 0) begin
        next_mux_d0_21 = input_word_d[168];
    end else if (sel_d0_21[2:0] == 1) begin
        next_mux_d0_21 = input_word_d[169];
    end else if (sel_d0_21[2:0] == 2) begin
        next_mux_d0_21 = input_word_d[170];
    end else if (sel_d0_21[2:0] == 3) begin
        next_mux_d0_21 = input_word_d[171];
    end else if (sel_d0_21[2:0] == 4) begin
        next_mux_d0_21 = input_word_d[172];
    end else if (sel_d0_21[2:0] == 5) begin
        next_mux_d0_21 = input_word_d[173];
    end else if (sel_d0_21[2:0] == 6) begin
        next_mux_d0_21 = input_word_d[174];
    end else begin
        next_mux_d0_21 = input_word_d[175];
    end

    if (sel_d0_22[2:0] == 0) begin
        next_mux_d0_22 = input_word_d[176];
    end else if (sel_d0_22[2:0] == 1) begin
        next_mux_d0_22 = input_word_d[177];
    end else if (sel_d0_22[2:0] == 2) begin
        next_mux_d0_22 = input_word_d[178];
    end else if (sel_d0_22[2:0] == 3) begin
        next_mux_d0_22 = input_word_d[179];
    end else if (sel_d0_22[2:0] == 4) begin
        next_mux_d0_22 = input_word_d[180];
    end else if (sel_d0_22[2:0] == 5) begin
        next_mux_d0_22 = input_word_d[181];
    end else if (sel_d0_22[2:0] == 6) begin
        next_mux_d0_22 = input_word_d[182];
    end else begin
        next_mux_d0_22 = input_word_d[183];
    end

    if (sel_d0_23[2:0] == 0) begin
        next_mux_d0_23 = input_word_d[184];
    end else if (sel_d0_23[2:0] == 1) begin
        next_mux_d0_23 = input_word_d[185];
    end else if (sel_d0_23[2:0] == 2) begin
        next_mux_d0_23 = input_word_d[186];
    end else if (sel_d0_23[2:0] == 3) begin
        next_mux_d0_23 = input_word_d[187];
    end else if (sel_d0_23[2:0] == 4) begin
        next_mux_d0_23 = input_word_d[188];
    end else if (sel_d0_23[2:0] == 5) begin
        next_mux_d0_23 = input_word_d[189];
    end else if (sel_d0_23[2:0] == 6) begin
        next_mux_d0_23 = input_word_d[190];
    end else begin
        next_mux_d0_23 = input_word_d[191];
    end

    if (sel_d0_24[2:0] == 0) begin
        next_mux_d0_24 = input_word_d[192];
    end else if (sel_d0_24[2:0] == 1) begin
        next_mux_d0_24 = input_word_d[193];
    end else if (sel_d0_24[2:0] == 2) begin
        next_mux_d0_24 = input_word_d[194];
    end else if (sel_d0_24[2:0] == 3) begin
        next_mux_d0_24 = input_word_d[195];
    end else if (sel_d0_24[2:0] == 4) begin
        next_mux_d0_24 = input_word_d[196];
    end else if (sel_d0_24[2:0] == 5) begin
        next_mux_d0_24 = input_word_d[197];
    end else if (sel_d0_24[2:0] == 6) begin
        next_mux_d0_24 = input_word_d[198];
    end else begin
        next_mux_d0_24 = input_word_d[199];
    end

    if (sel_d0_25[2:0] == 0) begin
        next_mux_d0_25 = input_word_d[200];
    end else if (sel_d0_25[2:0] == 1) begin
        next_mux_d0_25 = input_word_d[201];
    end else if (sel_d0_25[2:0] == 2) begin
        next_mux_d0_25 = input_word_d[202];
    end else if (sel_d0_25[2:0] == 3) begin
        next_mux_d0_25 = input_word_d[203];
    end else if (sel_d0_25[2:0] == 4) begin
        next_mux_d0_25 = input_word_d[204];
    end else if (sel_d0_25[2:0] == 5) begin
        next_mux_d0_25 = input_word_d[205];
    end else if (sel_d0_25[2:0] == 6) begin
        next_mux_d0_25 = input_word_d[206];
    end else begin
        next_mux_d0_25 = input_word_d[207];
    end

    if (sel_d0_26[2:0] == 0) begin
        next_mux_d0_26 = input_word_d[208];
    end else if (sel_d0_26[2:0] == 1) begin
        next_mux_d0_26 = input_word_d[209];
    end else if (sel_d0_26[2:0] == 2) begin
        next_mux_d0_26 = input_word_d[210];
    end else if (sel_d0_26[2:0] == 3) begin
        next_mux_d0_26 = input_word_d[211];
    end else if (sel_d0_26[2:0] == 4) begin
        next_mux_d0_26 = input_word_d[212];
    end else if (sel_d0_26[2:0] == 5) begin
        next_mux_d0_26 = input_word_d[213];
    end else if (sel_d0_26[2:0] == 6) begin
        next_mux_d0_26 = input_word_d[214];
    end else begin
        next_mux_d0_26 = input_word_d[215];
    end

    if (sel_d0_27[2:0] == 0) begin
        next_mux_d0_27 = input_word_d[216];
    end else if (sel_d0_27[2:0] == 1) begin
        next_mux_d0_27 = input_word_d[217];
    end else if (sel_d0_27[2:0] == 2) begin
        next_mux_d0_27 = input_word_d[218];
    end else if (sel_d0_27[2:0] == 3) begin
        next_mux_d0_27 = input_word_d[219];
    end else if (sel_d0_27[2:0] == 4) begin
        next_mux_d0_27 = input_word_d[220];
    end else if (sel_d0_27[2:0] == 5) begin
        next_mux_d0_27 = input_word_d[221];
    end else if (sel_d0_27[2:0] == 6) begin
        next_mux_d0_27 = input_word_d[222];
    end else begin
        next_mux_d0_27 = input_word_d[223];
    end

    if (sel_d0_28[2:0] == 0) begin
        next_mux_d0_28 = input_word_d[224];
    end else if (sel_d0_28[2:0] == 1) begin
        next_mux_d0_28 = input_word_d[225];
    end else if (sel_d0_28[2:0] == 2) begin
        next_mux_d0_28 = input_word_d[226];
    end else if (sel_d0_28[2:0] == 3) begin
        next_mux_d0_28 = input_word_d[227];
    end else if (sel_d0_28[2:0] == 4) begin
        next_mux_d0_28 = input_word_d[228];
    end else if (sel_d0_28[2:0] == 5) begin
        next_mux_d0_28 = input_word_d[229];
    end else if (sel_d0_28[2:0] == 6) begin
        next_mux_d0_28 = input_word_d[230];
    end else begin
        next_mux_d0_28 = input_word_d[231];
    end

    if (sel_d0_29[2:0] == 0) begin
        next_mux_d0_29 = input_word_d[232];
    end else if (sel_d0_29[2:0] == 1) begin
        next_mux_d0_29 = input_word_d[233];
    end else if (sel_d0_29[2:0] == 2) begin
        next_mux_d0_29 = input_word_d[234];
    end else if (sel_d0_29[2:0] == 3) begin
        next_mux_d0_29 = input_word_d[235];
    end else if (sel_d0_29[2:0] == 4) begin
        next_mux_d0_29 = input_word_d[236];
    end else if (sel_d0_29[2:0] == 5) begin
        next_mux_d0_29 = input_word_d[237];
    end else if (sel_d0_29[2:0] == 6) begin
        next_mux_d0_29 = input_word_d[238];
    end else begin
        next_mux_d0_29 = input_word_d[239];
    end

    if (sel_d0_30[2:0] == 0) begin
        next_mux_d0_30 = input_word_d[240];
    end else if (sel_d0_30[2:0] == 1) begin
        next_mux_d0_30 = input_word_d[241];
    end else if (sel_d0_30[2:0] == 2) begin
        next_mux_d0_30 = input_word_d[242];
    end else if (sel_d0_30[2:0] == 3) begin
        next_mux_d0_30 = input_word_d[243];
    end else if (sel_d0_30[2:0] == 4) begin
        next_mux_d0_30 = input_word_d[244];
    end else if (sel_d0_30[2:0] == 5) begin
        next_mux_d0_30 = input_word_d[245];
    end else if (sel_d0_30[2:0] == 6) begin
        next_mux_d0_30 = input_word_d[246];
    end else begin
        next_mux_d0_30 = input_word_d[247];
    end

    if (sel_d0_31[2:0] == 0) begin
        next_mux_d0_31 = input_word_d[248];
    end else if (sel_d0_31[2:0] == 1) begin
        next_mux_d0_31 = input_word_d[249];
    end else if (sel_d0_31[2:0] == 2) begin
        next_mux_d0_31 = input_word_d[250];
    end else if (sel_d0_31[2:0] == 3) begin
        next_mux_d0_31 = input_word_d[251];
    end else if (sel_d0_31[2:0] == 4) begin
        next_mux_d0_31 = input_word_d[252];
    end else if (sel_d0_31[2:0] == 5) begin
        next_mux_d0_31 = input_word_d[253];
    end else if (sel_d0_31[2:0] == 6) begin
        next_mux_d0_31 = input_word_d[254];
    end else begin
        next_mux_d0_31 = input_word_d[255];
    end

    if (sel_d0_32[2:0] == 0) begin
        next_mux_d0_32 = input_word_d[256];
    end else if (sel_d0_32[2:0] == 1) begin
        next_mux_d0_32 = input_word_d[257];
    end else if (sel_d0_32[2:0] == 2) begin
        next_mux_d0_32 = input_word_d[258];
    end else if (sel_d0_32[2:0] == 3) begin
        next_mux_d0_32 = input_word_d[259];
    end else if (sel_d0_32[2:0] == 4) begin
        next_mux_d0_32 = input_word_d[260];
    end else if (sel_d0_32[2:0] == 5) begin
        next_mux_d0_32 = input_word_d[261];
    end else if (sel_d0_32[2:0] == 6) begin
        next_mux_d0_32 = input_word_d[262];
    end else begin
        next_mux_d0_32 = input_word_d[263];
    end

    if (sel_d0_33[2:0] == 0) begin
        next_mux_d0_33 = input_word_d[264];
    end else if (sel_d0_33[2:0] == 1) begin
        next_mux_d0_33 = input_word_d[265];
    end else if (sel_d0_33[2:0] == 2) begin
        next_mux_d0_33 = input_word_d[266];
    end else if (sel_d0_33[2:0] == 3) begin
        next_mux_d0_33 = input_word_d[267];
    end else if (sel_d0_33[2:0] == 4) begin
        next_mux_d0_33 = input_word_d[268];
    end else if (sel_d0_33[2:0] == 5) begin
        next_mux_d0_33 = input_word_d[269];
    end else if (sel_d0_33[2:0] == 6) begin
        next_mux_d0_33 = input_word_d[270];
    end else begin
        next_mux_d0_33 = input_word_d[271];
    end

    if (sel_d0_34[2:0] == 0) begin
        next_mux_d0_34 = input_word_d[272];
    end else if (sel_d0_34[2:0] == 1) begin
        next_mux_d0_34 = input_word_d[273];
    end else if (sel_d0_34[2:0] == 2) begin
        next_mux_d0_34 = input_word_d[274];
    end else if (sel_d0_34[2:0] == 3) begin
        next_mux_d0_34 = input_word_d[275];
    end else if (sel_d0_34[2:0] == 4) begin
        next_mux_d0_34 = input_word_d[276];
    end else if (sel_d0_34[2:0] == 5) begin
        next_mux_d0_34 = input_word_d[277];
    end else if (sel_d0_34[2:0] == 6) begin
        next_mux_d0_34 = input_word_d[278];
    end else begin
        next_mux_d0_34 = input_word_d[279];
    end

    if (sel_d0_35[2:0] == 0) begin
        next_mux_d0_35 = input_word_d[280];
    end else if (sel_d0_35[2:0] == 1) begin
        next_mux_d0_35 = input_word_d[281];
    end else if (sel_d0_35[2:0] == 2) begin
        next_mux_d0_35 = input_word_d[282];
    end else if (sel_d0_35[2:0] == 3) begin
        next_mux_d0_35 = input_word_d[283];
    end else if (sel_d0_35[2:0] == 4) begin
        next_mux_d0_35 = input_word_d[284];
    end else if (sel_d0_35[2:0] == 5) begin
        next_mux_d0_35 = input_word_d[285];
    end else if (sel_d0_35[2:0] == 6) begin
        next_mux_d0_35 = input_word_d[286];
    end else begin
        next_mux_d0_35 = input_word_d[287];
    end

    if (sel_d0_36[2:0] == 0) begin
        next_mux_d0_36 = input_word_d[288];
    end else if (sel_d0_36[2:0] == 1) begin
        next_mux_d0_36 = input_word_d[289];
    end else if (sel_d0_36[2:0] == 2) begin
        next_mux_d0_36 = input_word_d[290];
    end else if (sel_d0_36[2:0] == 3) begin
        next_mux_d0_36 = input_word_d[291];
    end else if (sel_d0_36[2:0] == 4) begin
        next_mux_d0_36 = input_word_d[292];
    end else if (sel_d0_36[2:0] == 5) begin
        next_mux_d0_36 = input_word_d[293];
    end else if (sel_d0_36[2:0] == 6) begin
        next_mux_d0_36 = input_word_d[294];
    end else begin
        next_mux_d0_36 = input_word_d[295];
    end

    if (sel_d0_37[2:0] == 0) begin
        next_mux_d0_37 = input_word_d[296];
    end else if (sel_d0_37[2:0] == 1) begin
        next_mux_d0_37 = input_word_d[297];
    end else if (sel_d0_37[2:0] == 2) begin
        next_mux_d0_37 = input_word_d[298];
    end else if (sel_d0_37[2:0] == 3) begin
        next_mux_d0_37 = input_word_d[299];
    end else if (sel_d0_37[2:0] == 4) begin
        next_mux_d0_37 = input_word_d[300];
    end else if (sel_d0_37[2:0] == 5) begin
        next_mux_d0_37 = input_word_d[301];
    end else if (sel_d0_37[2:0] == 6) begin
        next_mux_d0_37 = input_word_d[302];
    end else begin
        next_mux_d0_37 = input_word_d[303];
    end

    if (sel_d0_38[2:0] == 0) begin
        next_mux_d0_38 = input_word_d[304];
    end else if (sel_d0_38[2:0] == 1) begin
        next_mux_d0_38 = input_word_d[305];
    end else if (sel_d0_38[2:0] == 2) begin
        next_mux_d0_38 = input_word_d[306];
    end else if (sel_d0_38[2:0] == 3) begin
        next_mux_d0_38 = input_word_d[307];
    end else if (sel_d0_38[2:0] == 4) begin
        next_mux_d0_38 = input_word_d[308];
    end else if (sel_d0_38[2:0] == 5) begin
        next_mux_d0_38 = input_word_d[309];
    end else if (sel_d0_38[2:0] == 6) begin
        next_mux_d0_38 = input_word_d[310];
    end else begin
        next_mux_d0_38 = input_word_d[311];
    end

    if (sel_d0_39[2:0] == 0) begin
        next_mux_d0_39 = input_word_d[312];
    end else if (sel_d0_39[2:0] == 1) begin
        next_mux_d0_39 = input_word_d[313];
    end else if (sel_d0_39[2:0] == 2) begin
        next_mux_d0_39 = input_word_d[314];
    end else if (sel_d0_39[2:0] == 3) begin
        next_mux_d0_39 = input_word_d[315];
    end else if (sel_d0_39[2:0] == 4) begin
        next_mux_d0_39 = input_word_d[316];
    end else if (sel_d0_39[2:0] == 5) begin
        next_mux_d0_39 = input_word_d[317];
    end else if (sel_d0_39[2:0] == 6) begin
        next_mux_d0_39 = input_word_d[318];
    end else begin
        next_mux_d0_39 = input_word_d[319];
    end

    if (sel_d0_40[2:0] == 0) begin
        next_mux_d0_40 = input_word_d[320];
    end else if (sel_d0_40[2:0] == 1) begin
        next_mux_d0_40 = input_word_d[321];
    end else if (sel_d0_40[2:0] == 2) begin
        next_mux_d0_40 = input_word_d[322];
    end else if (sel_d0_40[2:0] == 3) begin
        next_mux_d0_40 = input_word_d[323];
    end else if (sel_d0_40[2:0] == 4) begin
        next_mux_d0_40 = input_word_d[324];
    end else if (sel_d0_40[2:0] == 5) begin
        next_mux_d0_40 = input_word_d[325];
    end else if (sel_d0_40[2:0] == 6) begin
        next_mux_d0_40 = input_word_d[326];
    end else begin
        next_mux_d0_40 = input_word_d[327];
    end

    if (sel_d0_41[2:0] == 0) begin
        next_mux_d0_41 = input_word_d[328];
    end else if (sel_d0_41[2:0] == 1) begin
        next_mux_d0_41 = input_word_d[329];
    end else if (sel_d0_41[2:0] == 2) begin
        next_mux_d0_41 = input_word_d[330];
    end else if (sel_d0_41[2:0] == 3) begin
        next_mux_d0_41 = input_word_d[331];
    end else if (sel_d0_41[2:0] == 4) begin
        next_mux_d0_41 = input_word_d[332];
    end else if (sel_d0_41[2:0] == 5) begin
        next_mux_d0_41 = input_word_d[333];
    end else if (sel_d0_41[2:0] == 6) begin
        next_mux_d0_41 = input_word_d[334];
    end else begin
        next_mux_d0_41 = input_word_d[335];
    end

    if (sel_d0_42[2:0] == 0) begin
        next_mux_d0_42 = input_word_d[336];
    end else if (sel_d0_42[2:0] == 1) begin
        next_mux_d0_42 = input_word_d[337];
    end else if (sel_d0_42[2:0] == 2) begin
        next_mux_d0_42 = input_word_d[338];
    end else if (sel_d0_42[2:0] == 3) begin
        next_mux_d0_42 = input_word_d[339];
    end else if (sel_d0_42[2:0] == 4) begin
        next_mux_d0_42 = input_word_d[340];
    end else if (sel_d0_42[2:0] == 5) begin
        next_mux_d0_42 = input_word_d[341];
    end else if (sel_d0_42[2:0] == 6) begin
        next_mux_d0_42 = input_word_d[342];
    end else begin
        next_mux_d0_42 = input_word_d[343];
    end

    if (sel_d0_43[2:0] == 0) begin
        next_mux_d0_43 = input_word_d[344];
    end else if (sel_d0_43[2:0] == 1) begin
        next_mux_d0_43 = input_word_d[345];
    end else if (sel_d0_43[2:0] == 2) begin
        next_mux_d0_43 = input_word_d[346];
    end else if (sel_d0_43[2:0] == 3) begin
        next_mux_d0_43 = input_word_d[347];
    end else if (sel_d0_43[2:0] == 4) begin
        next_mux_d0_43 = input_word_d[348];
    end else if (sel_d0_43[2:0] == 5) begin
        next_mux_d0_43 = input_word_d[349];
    end else if (sel_d0_43[2:0] == 6) begin
        next_mux_d0_43 = input_word_d[350];
    end else begin
        next_mux_d0_43 = input_word_d[351];
    end

    if (sel_d0_44[2:0] == 0) begin
        next_mux_d0_44 = input_word_d[352];
    end else if (sel_d0_44[2:0] == 1) begin
        next_mux_d0_44 = input_word_d[353];
    end else if (sel_d0_44[2:0] == 2) begin
        next_mux_d0_44 = input_word_d[354];
    end else if (sel_d0_44[2:0] == 3) begin
        next_mux_d0_44 = input_word_d[355];
    end else if (sel_d0_44[2:0] == 4) begin
        next_mux_d0_44 = input_word_d[356];
    end else if (sel_d0_44[2:0] == 5) begin
        next_mux_d0_44 = input_word_d[357];
    end else if (sel_d0_44[2:0] == 6) begin
        next_mux_d0_44 = input_word_d[358];
    end else begin
        next_mux_d0_44 = input_word_d[359];
    end

    if (sel_d0_45[2:0] == 0) begin
        next_mux_d0_45 = input_word_d[360];
    end else if (sel_d0_45[2:0] == 1) begin
        next_mux_d0_45 = input_word_d[361];
    end else if (sel_d0_45[2:0] == 2) begin
        next_mux_d0_45 = input_word_d[362];
    end else if (sel_d0_45[2:0] == 3) begin
        next_mux_d0_45 = input_word_d[363];
    end else if (sel_d0_45[2:0] == 4) begin
        next_mux_d0_45 = input_word_d[364];
    end else if (sel_d0_45[2:0] == 5) begin
        next_mux_d0_45 = input_word_d[365];
    end else if (sel_d0_45[2:0] == 6) begin
        next_mux_d0_45 = input_word_d[366];
    end else begin
        next_mux_d0_45 = input_word_d[367];
    end

    if (sel_d0_46[2:0] == 0) begin
        next_mux_d0_46 = input_word_d[368];
    end else if (sel_d0_46[2:0] == 1) begin
        next_mux_d0_46 = input_word_d[369];
    end else if (sel_d0_46[2:0] == 2) begin
        next_mux_d0_46 = input_word_d[370];
    end else if (sel_d0_46[2:0] == 3) begin
        next_mux_d0_46 = input_word_d[371];
    end else if (sel_d0_46[2:0] == 4) begin
        next_mux_d0_46 = input_word_d[372];
    end else if (sel_d0_46[2:0] == 5) begin
        next_mux_d0_46 = input_word_d[373];
    end else if (sel_d0_46[2:0] == 6) begin
        next_mux_d0_46 = input_word_d[374];
    end else begin
        next_mux_d0_46 = input_word_d[375];
    end

    if (sel_d0_47[2:0] == 0) begin
        next_mux_d0_47 = input_word_d[376];
    end else if (sel_d0_47[2:0] == 1) begin
        next_mux_d0_47 = input_word_d[377];
    end else if (sel_d0_47[2:0] == 2) begin
        next_mux_d0_47 = input_word_d[378];
    end else if (sel_d0_47[2:0] == 3) begin
        next_mux_d0_47 = input_word_d[379];
    end else if (sel_d0_47[2:0] == 4) begin
        next_mux_d0_47 = input_word_d[380];
    end else if (sel_d0_47[2:0] == 5) begin
        next_mux_d0_47 = input_word_d[381];
    end else if (sel_d0_47[2:0] == 6) begin
        next_mux_d0_47 = input_word_d[382];
    end else begin
        next_mux_d0_47 = input_word_d[383];
    end

    if (sel_d0_48[2:0] == 0) begin
        next_mux_d0_48 = input_word_d[384];
    end else if (sel_d0_48[2:0] == 1) begin
        next_mux_d0_48 = input_word_d[385];
    end else if (sel_d0_48[2:0] == 2) begin
        next_mux_d0_48 = input_word_d[386];
    end else if (sel_d0_48[2:0] == 3) begin
        next_mux_d0_48 = input_word_d[387];
    end else if (sel_d0_48[2:0] == 4) begin
        next_mux_d0_48 = input_word_d[388];
    end else if (sel_d0_48[2:0] == 5) begin
        next_mux_d0_48 = input_word_d[389];
    end else if (sel_d0_48[2:0] == 6) begin
        next_mux_d0_48 = input_word_d[390];
    end else begin
        next_mux_d0_48 = input_word_d[391];
    end

    if (sel_d0_49[2:0] == 0) begin
        next_mux_d0_49 = input_word_d[392];
    end else if (sel_d0_49[2:0] == 1) begin
        next_mux_d0_49 = input_word_d[393];
    end else if (sel_d0_49[2:0] == 2) begin
        next_mux_d0_49 = input_word_d[394];
    end else if (sel_d0_49[2:0] == 3) begin
        next_mux_d0_49 = input_word_d[395];
    end else if (sel_d0_49[2:0] == 4) begin
        next_mux_d0_49 = input_word_d[396];
    end else if (sel_d0_49[2:0] == 5) begin
        next_mux_d0_49 = input_word_d[397];
    end else if (sel_d0_49[2:0] == 6) begin
        next_mux_d0_49 = input_word_d[398];
    end else begin
        next_mux_d0_49 = input_word_d[399];
    end

    if (sel_d0_50[2:0] == 0) begin
        next_mux_d0_50 = input_word_d[400];
    end else if (sel_d0_50[2:0] == 1) begin
        next_mux_d0_50 = input_word_d[401];
    end else if (sel_d0_50[2:0] == 2) begin
        next_mux_d0_50 = input_word_d[402];
    end else if (sel_d0_50[2:0] == 3) begin
        next_mux_d0_50 = input_word_d[403];
    end else if (sel_d0_50[2:0] == 4) begin
        next_mux_d0_50 = input_word_d[404];
    end else if (sel_d0_50[2:0] == 5) begin
        next_mux_d0_50 = input_word_d[405];
    end else if (sel_d0_50[2:0] == 6) begin
        next_mux_d0_50 = input_word_d[406];
    end else begin
        next_mux_d0_50 = input_word_d[407];
    end

    if (sel_d0_51[2:0] == 0) begin
        next_mux_d0_51 = input_word_d[408];
    end else if (sel_d0_51[2:0] == 1) begin
        next_mux_d0_51 = input_word_d[409];
    end else if (sel_d0_51[2:0] == 2) begin
        next_mux_d0_51 = input_word_d[410];
    end else if (sel_d0_51[2:0] == 3) begin
        next_mux_d0_51 = input_word_d[411];
    end else if (sel_d0_51[2:0] == 4) begin
        next_mux_d0_51 = input_word_d[412];
    end else if (sel_d0_51[2:0] == 5) begin
        next_mux_d0_51 = input_word_d[413];
    end else if (sel_d0_51[2:0] == 6) begin
        next_mux_d0_51 = input_word_d[414];
    end else begin
        next_mux_d0_51 = input_word_d[415];
    end

    if (sel_d0_52[2:0] == 0) begin
        next_mux_d0_52 = input_word_d[416];
    end else if (sel_d0_52[2:0] == 1) begin
        next_mux_d0_52 = input_word_d[417];
    end else if (sel_d0_52[2:0] == 2) begin
        next_mux_d0_52 = input_word_d[418];
    end else if (sel_d0_52[2:0] == 3) begin
        next_mux_d0_52 = input_word_d[419];
    end else if (sel_d0_52[2:0] == 4) begin
        next_mux_d0_52 = input_word_d[420];
    end else if (sel_d0_52[2:0] == 5) begin
        next_mux_d0_52 = input_word_d[421];
    end else if (sel_d0_52[2:0] == 6) begin
        next_mux_d0_52 = input_word_d[422];
    end else begin
        next_mux_d0_52 = input_word_d[423];
    end

    if (sel_d0_53[2:0] == 0) begin
        next_mux_d0_53 = input_word_d[424];
    end else if (sel_d0_53[2:0] == 1) begin
        next_mux_d0_53 = input_word_d[425];
    end else if (sel_d0_53[2:0] == 2) begin
        next_mux_d0_53 = input_word_d[426];
    end else if (sel_d0_53[2:0] == 3) begin
        next_mux_d0_53 = input_word_d[427];
    end else if (sel_d0_53[2:0] == 4) begin
        next_mux_d0_53 = input_word_d[428];
    end else if (sel_d0_53[2:0] == 5) begin
        next_mux_d0_53 = input_word_d[429];
    end else if (sel_d0_53[2:0] == 6) begin
        next_mux_d0_53 = input_word_d[430];
    end else begin
        next_mux_d0_53 = input_word_d[431];
    end

    if (sel_d0_54[2:0] == 0) begin
        next_mux_d0_54 = input_word_d[432];
    end else if (sel_d0_54[2:0] == 1) begin
        next_mux_d0_54 = input_word_d[433];
    end else if (sel_d0_54[2:0] == 2) begin
        next_mux_d0_54 = input_word_d[434];
    end else if (sel_d0_54[2:0] == 3) begin
        next_mux_d0_54 = input_word_d[435];
    end else if (sel_d0_54[2:0] == 4) begin
        next_mux_d0_54 = input_word_d[436];
    end else if (sel_d0_54[2:0] == 5) begin
        next_mux_d0_54 = input_word_d[437];
    end else if (sel_d0_54[2:0] == 6) begin
        next_mux_d0_54 = input_word_d[438];
    end else begin
        next_mux_d0_54 = input_word_d[439];
    end

    if (sel_d0_55[2:0] == 0) begin
        next_mux_d0_55 = input_word_d[440];
    end else if (sel_d0_55[2:0] == 1) begin
        next_mux_d0_55 = input_word_d[441];
    end else if (sel_d0_55[2:0] == 2) begin
        next_mux_d0_55 = input_word_d[442];
    end else if (sel_d0_55[2:0] == 3) begin
        next_mux_d0_55 = input_word_d[443];
    end else if (sel_d0_55[2:0] == 4) begin
        next_mux_d0_55 = input_word_d[444];
    end else if (sel_d0_55[2:0] == 5) begin
        next_mux_d0_55 = input_word_d[445];
    end else if (sel_d0_55[2:0] == 6) begin
        next_mux_d0_55 = input_word_d[446];
    end else begin
        next_mux_d0_55 = input_word_d[447];
    end

    if (sel_d0_56[2:0] == 0) begin
        next_mux_d0_56 = input_word_d[448];
    end else if (sel_d0_56[2:0] == 1) begin
        next_mux_d0_56 = input_word_d[449];
    end else if (sel_d0_56[2:0] == 2) begin
        next_mux_d0_56 = input_word_d[450];
    end else if (sel_d0_56[2:0] == 3) begin
        next_mux_d0_56 = input_word_d[451];
    end else if (sel_d0_56[2:0] == 4) begin
        next_mux_d0_56 = input_word_d[452];
    end else if (sel_d0_56[2:0] == 5) begin
        next_mux_d0_56 = input_word_d[453];
    end else if (sel_d0_56[2:0] == 6) begin
        next_mux_d0_56 = input_word_d[454];
    end else begin
        next_mux_d0_56 = input_word_d[455];
    end

    if (sel_d0_57[2:0] == 0) begin
        next_mux_d0_57 = input_word_d[456];
    end else if (sel_d0_57[2:0] == 1) begin
        next_mux_d0_57 = input_word_d[457];
    end else if (sel_d0_57[2:0] == 2) begin
        next_mux_d0_57 = input_word_d[458];
    end else if (sel_d0_57[2:0] == 3) begin
        next_mux_d0_57 = input_word_d[459];
    end else if (sel_d0_57[2:0] == 4) begin
        next_mux_d0_57 = input_word_d[460];
    end else if (sel_d0_57[2:0] == 5) begin
        next_mux_d0_57 = input_word_d[461];
    end else if (sel_d0_57[2:0] == 6) begin
        next_mux_d0_57 = input_word_d[462];
    end else begin
        next_mux_d0_57 = input_word_d[463];
    end

    if (sel_d0_58[2:0] == 0) begin
        next_mux_d0_58 = input_word_d[464];
    end else if (sel_d0_58[2:0] == 1) begin
        next_mux_d0_58 = input_word_d[465];
    end else if (sel_d0_58[2:0] == 2) begin
        next_mux_d0_58 = input_word_d[466];
    end else if (sel_d0_58[2:0] == 3) begin
        next_mux_d0_58 = input_word_d[467];
    end else if (sel_d0_58[2:0] == 4) begin
        next_mux_d0_58 = input_word_d[468];
    end else if (sel_d0_58[2:0] == 5) begin
        next_mux_d0_58 = input_word_d[469];
    end else if (sel_d0_58[2:0] == 6) begin
        next_mux_d0_58 = input_word_d[470];
    end else begin
        next_mux_d0_58 = input_word_d[471];
    end

    if (sel_d0_59[2:0] == 0) begin
        next_mux_d0_59 = input_word_d[472];
    end else if (sel_d0_59[2:0] == 1) begin
        next_mux_d0_59 = input_word_d[473];
    end else if (sel_d0_59[2:0] == 2) begin
        next_mux_d0_59 = input_word_d[474];
    end else if (sel_d0_59[2:0] == 3) begin
        next_mux_d0_59 = input_word_d[475];
    end else if (sel_d0_59[2:0] == 4) begin
        next_mux_d0_59 = input_word_d[476];
    end else if (sel_d0_59[2:0] == 5) begin
        next_mux_d0_59 = input_word_d[477];
    end else if (sel_d0_59[2:0] == 6) begin
        next_mux_d0_59 = input_word_d[478];
    end else begin
        next_mux_d0_59 = input_word_d[479];
    end

    if (sel_d0_60[2:0] == 0) begin
        next_mux_d0_60 = input_word_d[480];
    end else if (sel_d0_60[2:0] == 1) begin
        next_mux_d0_60 = input_word_d[481];
    end else if (sel_d0_60[2:0] == 2) begin
        next_mux_d0_60 = input_word_d[482];
    end else if (sel_d0_60[2:0] == 3) begin
        next_mux_d0_60 = input_word_d[483];
    end else if (sel_d0_60[2:0] == 4) begin
        next_mux_d0_60 = input_word_d[484];
    end else if (sel_d0_60[2:0] == 5) begin
        next_mux_d0_60 = input_word_d[485];
    end else if (sel_d0_60[2:0] == 6) begin
        next_mux_d0_60 = input_word_d[486];
    end else begin
        next_mux_d0_60 = input_word_d[487];
    end

    if (sel_d0_61[2:0] == 0) begin
        next_mux_d0_61 = input_word_d[488];
    end else if (sel_d0_61[2:0] == 1) begin
        next_mux_d0_61 = input_word_d[489];
    end else if (sel_d0_61[2:0] == 2) begin
        next_mux_d0_61 = input_word_d[490];
    end else if (sel_d0_61[2:0] == 3) begin
        next_mux_d0_61 = input_word_d[491];
    end else if (sel_d0_61[2:0] == 4) begin
        next_mux_d0_61 = input_word_d[492];
    end else if (sel_d0_61[2:0] == 5) begin
        next_mux_d0_61 = input_word_d[493];
    end else if (sel_d0_61[2:0] == 6) begin
        next_mux_d0_61 = input_word_d[494];
    end else begin
        next_mux_d0_61 = input_word_d[495];
    end

    if (sel_d0_62[2:0] == 0) begin
        next_mux_d0_62 = input_word_d[496];
    end else if (sel_d0_62[2:0] == 1) begin
        next_mux_d0_62 = input_word_d[497];
    end else if (sel_d0_62[2:0] == 2) begin
        next_mux_d0_62 = input_word_d[498];
    end else if (sel_d0_62[2:0] == 3) begin
        next_mux_d0_62 = input_word_d[499];
    end else if (sel_d0_62[2:0] == 4) begin
        next_mux_d0_62 = input_word_d[500];
    end else if (sel_d0_62[2:0] == 5) begin
        next_mux_d0_62 = input_word_d[501];
    end else if (sel_d0_62[2:0] == 6) begin
        next_mux_d0_62 = input_word_d[502];
    end else begin
        next_mux_d0_62 = input_word_d[503];
    end

    if (sel_d0_63[2:0] == 0) begin
        next_mux_d0_63 = input_word_d[504];
    end else if (sel_d0_63[2:0] == 1) begin
        next_mux_d0_63 = input_word_d[505];
    end else if (sel_d0_63[2:0] == 2) begin
        next_mux_d0_63 = input_word_d[506];
    end else if (sel_d0_63[2:0] == 3) begin
        next_mux_d0_63 = input_word_d[507];
    end else if (sel_d0_63[2:0] == 4) begin
        next_mux_d0_63 = input_word_d[508];
    end else if (sel_d0_63[2:0] == 5) begin
        next_mux_d0_63 = input_word_d[509];
    end else if (sel_d0_63[2:0] == 6) begin
        next_mux_d0_63 = input_word_d[510];
    end else begin
        next_mux_d0_63 = input_word_d[511];
    end

    if (sel_d1_0[5:3] == 0) begin
        next_mux_d1_0 = mux_d0_0;
    end else if (sel_d1_0[5:3] == 1) begin
        next_mux_d1_0 = mux_d0_1;
    end else if (sel_d1_0[5:3] == 2) begin
        next_mux_d1_0 = mux_d0_2;
    end else if (sel_d1_0[5:3] == 3) begin
        next_mux_d1_0 = mux_d0_3;
    end else if (sel_d1_0[5:3] == 4) begin
        next_mux_d1_0 = mux_d0_4;
    end else if (sel_d1_0[5:3] == 5) begin
        next_mux_d1_0 = mux_d0_5;
    end else if (sel_d1_0[5:3] == 6) begin
        next_mux_d1_0 = mux_d0_6;
    end else begin
        next_mux_d1_0 = mux_d0_7;
    end

    if (sel_d1_1[5:3] == 0) begin
        next_mux_d1_1 = mux_d0_8;
    end else if (sel_d1_1[5:3] == 1) begin
        next_mux_d1_1 = mux_d0_9;
    end else if (sel_d1_1[5:3] == 2) begin
        next_mux_d1_1 = mux_d0_10;
    end else if (sel_d1_1[5:3] == 3) begin
        next_mux_d1_1 = mux_d0_11;
    end else if (sel_d1_1[5:3] == 4) begin
        next_mux_d1_1 = mux_d0_12;
    end else if (sel_d1_1[5:3] == 5) begin
        next_mux_d1_1 = mux_d0_13;
    end else if (sel_d1_1[5:3] == 6) begin
        next_mux_d1_1 = mux_d0_14;
    end else begin
        next_mux_d1_1 = mux_d0_15;
    end

    if (sel_d1_2[5:3] == 0) begin
        next_mux_d1_2 = mux_d0_16;
    end else if (sel_d1_2[5:3] == 1) begin
        next_mux_d1_2 = mux_d0_17;
    end else if (sel_d1_2[5:3] == 2) begin
        next_mux_d1_2 = mux_d0_18;
    end else if (sel_d1_2[5:3] == 3) begin
        next_mux_d1_2 = mux_d0_19;
    end else if (sel_d1_2[5:3] == 4) begin
        next_mux_d1_2 = mux_d0_20;
    end else if (sel_d1_2[5:3] == 5) begin
        next_mux_d1_2 = mux_d0_21;
    end else if (sel_d1_2[5:3] == 6) begin
        next_mux_d1_2 = mux_d0_22;
    end else begin
        next_mux_d1_2 = mux_d0_23;
    end

    if (sel_d1_3[5:3] == 0) begin
        next_mux_d1_3 = mux_d0_24;
    end else if (sel_d1_3[5:3] == 1) begin
        next_mux_d1_3 = mux_d0_25;
    end else if (sel_d1_3[5:3] == 2) begin
        next_mux_d1_3 = mux_d0_26;
    end else if (sel_d1_3[5:3] == 3) begin
        next_mux_d1_3 = mux_d0_27;
    end else if (sel_d1_3[5:3] == 4) begin
        next_mux_d1_3 = mux_d0_28;
    end else if (sel_d1_3[5:3] == 5) begin
        next_mux_d1_3 = mux_d0_29;
    end else if (sel_d1_3[5:3] == 6) begin
        next_mux_d1_3 = mux_d0_30;
    end else begin
        next_mux_d1_3 = mux_d0_31;
    end

    if (sel_d1_4[5:3] == 0) begin
        next_mux_d1_4 = mux_d0_32;
    end else if (sel_d1_4[5:3] == 1) begin
        next_mux_d1_4 = mux_d0_33;
    end else if (sel_d1_4[5:3] == 2) begin
        next_mux_d1_4 = mux_d0_34;
    end else if (sel_d1_4[5:3] == 3) begin
        next_mux_d1_4 = mux_d0_35;
    end else if (sel_d1_4[5:3] == 4) begin
        next_mux_d1_4 = mux_d0_36;
    end else if (sel_d1_4[5:3] == 5) begin
        next_mux_d1_4 = mux_d0_37;
    end else if (sel_d1_4[5:3] == 6) begin
        next_mux_d1_4 = mux_d0_38;
    end else begin
        next_mux_d1_4 = mux_d0_39;
    end

    if (sel_d1_5[5:3] == 0) begin
        next_mux_d1_5 = mux_d0_40;
    end else if (sel_d1_5[5:3] == 1) begin
        next_mux_d1_5 = mux_d0_41;
    end else if (sel_d1_5[5:3] == 2) begin
        next_mux_d1_5 = mux_d0_42;
    end else if (sel_d1_5[5:3] == 3) begin
        next_mux_d1_5 = mux_d0_43;
    end else if (sel_d1_5[5:3] == 4) begin
        next_mux_d1_5 = mux_d0_44;
    end else if (sel_d1_5[5:3] == 5) begin
        next_mux_d1_5 = mux_d0_45;
    end else if (sel_d1_5[5:3] == 6) begin
        next_mux_d1_5 = mux_d0_46;
    end else begin
        next_mux_d1_5 = mux_d0_47;
    end

    if (sel_d1_6[5:3] == 0) begin
        next_mux_d1_6 = mux_d0_48;
    end else if (sel_d1_6[5:3] == 1) begin
        next_mux_d1_6 = mux_d0_49;
    end else if (sel_d1_6[5:3] == 2) begin
        next_mux_d1_6 = mux_d0_50;
    end else if (sel_d1_6[5:3] == 3) begin
        next_mux_d1_6 = mux_d0_51;
    end else if (sel_d1_6[5:3] == 4) begin
        next_mux_d1_6 = mux_d0_52;
    end else if (sel_d1_6[5:3] == 5) begin
        next_mux_d1_6 = mux_d0_53;
    end else if (sel_d1_6[5:3] == 6) begin
        next_mux_d1_6 = mux_d0_54;
    end else begin
        next_mux_d1_6 = mux_d0_55;
    end

    if (sel_d1_7[5:3] == 0) begin
        next_mux_d1_7 = mux_d0_56;
    end else if (sel_d1_7[5:3] == 1) begin
        next_mux_d1_7 = mux_d0_57;
    end else if (sel_d1_7[5:3] == 2) begin
        next_mux_d1_7 = mux_d0_58;
    end else if (sel_d1_7[5:3] == 3) begin
        next_mux_d1_7 = mux_d0_59;
    end else if (sel_d1_7[5:3] == 4) begin
        next_mux_d1_7 = mux_d0_60;
    end else if (sel_d1_7[5:3] == 5) begin
        next_mux_d1_7 = mux_d0_61;
    end else if (sel_d1_7[5:3] == 6) begin
        next_mux_d1_7 = mux_d0_62;
    end else begin
        next_mux_d1_7 = mux_d0_63;
    end

    if (sel_d2_0[8:6] == 0) begin
        next_mux_d2_0 = mux_d1_0;
    end else if (sel_d2_0[8:6] == 1) begin
        next_mux_d2_0 = mux_d1_1;
    end else if (sel_d2_0[8:6] == 2) begin
        next_mux_d2_0 = mux_d1_2;
    end else if (sel_d2_0[8:6] == 3) begin
        next_mux_d2_0 = mux_d1_3;
    end else if (sel_d2_0[8:6] == 4) begin
        next_mux_d2_0 = mux_d1_4;
    end else if (sel_d2_0[8:6] == 5) begin
        next_mux_d2_0 = mux_d1_5;
    end else if (sel_d2_0[8:6] == 6) begin
        next_mux_d2_0 = mux_d1_6;
    end else begin
        next_mux_d2_0 = mux_d1_7;
    end

end

endmodule
