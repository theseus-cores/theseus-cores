//
// Macros used only in simulation.
//
//
`ifdef SIM_BIN_WRITE
`undef SIM_BIN_WRITE
`endif
