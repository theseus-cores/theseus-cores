/*************************************************************************/
//// File        : pipe_mux_2048_1.v
// Description : Implements a pipelined multiplexer to be used in high speed design
// This module has a delay of 5 clock cycles//
// -------------------------------------------------------------------
//
/***************************************************************************/


module pipe_mux_2048_1
(
    input clk,
    input sync_reset,
    input valid_i,
    input [10:0] sel,
    input [2047:0] input_word,
    output valid_o,
    output [10:0] sel_o,
    output output_word
);

(* KEEP = "TRUE" *) reg [10:0] sel_d0_0;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_1;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_2;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_3;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_4;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_5;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_6;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_7;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_8;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_9;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_10;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_11;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_12;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_13;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_14;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_15;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_16;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_17;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_18;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_19;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_20;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_21;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_22;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_23;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_24;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_25;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_26;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_27;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_28;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_29;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_30;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_31;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_32;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_33;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_34;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_35;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_36;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_37;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_38;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_39;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_40;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_41;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_42;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_43;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_44;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_45;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_46;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_47;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_48;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_49;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_50;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_51;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_52;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_53;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_54;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_55;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_56;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_57;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_58;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_59;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_60;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_61;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_62;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_63;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_64;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_65;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_66;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_67;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_68;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_69;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_70;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_71;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_72;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_73;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_74;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_75;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_76;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_77;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_78;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_79;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_80;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_81;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_82;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_83;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_84;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_85;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_86;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_87;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_88;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_89;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_90;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_91;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_92;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_93;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_94;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_95;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_96;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_97;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_98;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_99;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_100;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_101;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_102;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_103;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_104;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_105;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_106;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_107;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_108;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_109;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_110;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_111;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_112;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_113;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_114;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_115;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_116;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_117;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_118;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_119;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_120;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_121;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_122;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_123;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_124;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_125;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_126;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_127;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_128;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_129;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_130;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_131;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_132;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_133;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_134;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_135;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_136;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_137;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_138;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_139;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_140;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_141;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_142;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_143;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_144;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_145;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_146;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_147;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_148;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_149;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_150;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_151;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_152;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_153;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_154;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_155;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_156;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_157;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_158;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_159;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_160;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_161;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_162;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_163;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_164;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_165;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_166;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_167;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_168;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_169;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_170;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_171;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_172;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_173;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_174;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_175;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_176;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_177;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_178;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_179;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_180;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_181;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_182;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_183;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_184;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_185;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_186;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_187;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_188;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_189;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_190;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_191;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_192;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_193;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_194;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_195;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_196;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_197;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_198;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_199;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_200;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_201;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_202;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_203;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_204;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_205;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_206;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_207;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_208;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_209;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_210;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_211;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_212;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_213;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_214;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_215;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_216;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_217;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_218;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_219;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_220;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_221;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_222;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_223;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_224;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_225;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_226;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_227;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_228;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_229;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_230;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_231;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_232;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_233;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_234;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_235;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_236;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_237;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_238;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_239;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_240;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_241;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_242;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_243;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_244;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_245;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_246;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_247;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_248;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_249;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_250;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_251;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_252;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_253;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_254;
(* KEEP = "TRUE" *) reg [10:0] sel_d0_255;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_0;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_1;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_2;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_3;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_4;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_5;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_6;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_7;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_8;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_9;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_10;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_11;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_12;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_13;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_14;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_15;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_16;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_17;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_18;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_19;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_20;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_21;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_22;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_23;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_24;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_25;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_26;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_27;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_28;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_29;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_30;
(* KEEP = "TRUE" *) reg [10:0] sel_d1_31;
(* KEEP = "TRUE" *) reg [10:0] sel_d2_0;
(* KEEP = "TRUE" *) reg [10:0] sel_d2_1;
(* KEEP = "TRUE" *) reg [10:0] sel_d2_2;
(* KEEP = "TRUE" *) reg [10:0] sel_d2_3;
(* KEEP = "TRUE" *) reg [10:0] sel_d3_0;
(* KEEP = "TRUE" *) reg [10:0] sel_d4;
reg valid_d0;
reg valid_d1;
reg valid_d2;
reg valid_d3;
reg valid_d4;
reg [0:0] mux_d0_0, next_mux_d0_0;
reg [0:0] mux_d0_1, next_mux_d0_1;
reg [0:0] mux_d0_2, next_mux_d0_2;
reg [0:0] mux_d0_3, next_mux_d0_3;
reg [0:0] mux_d0_4, next_mux_d0_4;
reg [0:0] mux_d0_5, next_mux_d0_5;
reg [0:0] mux_d0_6, next_mux_d0_6;
reg [0:0] mux_d0_7, next_mux_d0_7;
reg [0:0] mux_d0_8, next_mux_d0_8;
reg [0:0] mux_d0_9, next_mux_d0_9;
reg [0:0] mux_d0_10, next_mux_d0_10;
reg [0:0] mux_d0_11, next_mux_d0_11;
reg [0:0] mux_d0_12, next_mux_d0_12;
reg [0:0] mux_d0_13, next_mux_d0_13;
reg [0:0] mux_d0_14, next_mux_d0_14;
reg [0:0] mux_d0_15, next_mux_d0_15;
reg [0:0] mux_d0_16, next_mux_d0_16;
reg [0:0] mux_d0_17, next_mux_d0_17;
reg [0:0] mux_d0_18, next_mux_d0_18;
reg [0:0] mux_d0_19, next_mux_d0_19;
reg [0:0] mux_d0_20, next_mux_d0_20;
reg [0:0] mux_d0_21, next_mux_d0_21;
reg [0:0] mux_d0_22, next_mux_d0_22;
reg [0:0] mux_d0_23, next_mux_d0_23;
reg [0:0] mux_d0_24, next_mux_d0_24;
reg [0:0] mux_d0_25, next_mux_d0_25;
reg [0:0] mux_d0_26, next_mux_d0_26;
reg [0:0] mux_d0_27, next_mux_d0_27;
reg [0:0] mux_d0_28, next_mux_d0_28;
reg [0:0] mux_d0_29, next_mux_d0_29;
reg [0:0] mux_d0_30, next_mux_d0_30;
reg [0:0] mux_d0_31, next_mux_d0_31;
reg [0:0] mux_d0_32, next_mux_d0_32;
reg [0:0] mux_d0_33, next_mux_d0_33;
reg [0:0] mux_d0_34, next_mux_d0_34;
reg [0:0] mux_d0_35, next_mux_d0_35;
reg [0:0] mux_d0_36, next_mux_d0_36;
reg [0:0] mux_d0_37, next_mux_d0_37;
reg [0:0] mux_d0_38, next_mux_d0_38;
reg [0:0] mux_d0_39, next_mux_d0_39;
reg [0:0] mux_d0_40, next_mux_d0_40;
reg [0:0] mux_d0_41, next_mux_d0_41;
reg [0:0] mux_d0_42, next_mux_d0_42;
reg [0:0] mux_d0_43, next_mux_d0_43;
reg [0:0] mux_d0_44, next_mux_d0_44;
reg [0:0] mux_d0_45, next_mux_d0_45;
reg [0:0] mux_d0_46, next_mux_d0_46;
reg [0:0] mux_d0_47, next_mux_d0_47;
reg [0:0] mux_d0_48, next_mux_d0_48;
reg [0:0] mux_d0_49, next_mux_d0_49;
reg [0:0] mux_d0_50, next_mux_d0_50;
reg [0:0] mux_d0_51, next_mux_d0_51;
reg [0:0] mux_d0_52, next_mux_d0_52;
reg [0:0] mux_d0_53, next_mux_d0_53;
reg [0:0] mux_d0_54, next_mux_d0_54;
reg [0:0] mux_d0_55, next_mux_d0_55;
reg [0:0] mux_d0_56, next_mux_d0_56;
reg [0:0] mux_d0_57, next_mux_d0_57;
reg [0:0] mux_d0_58, next_mux_d0_58;
reg [0:0] mux_d0_59, next_mux_d0_59;
reg [0:0] mux_d0_60, next_mux_d0_60;
reg [0:0] mux_d0_61, next_mux_d0_61;
reg [0:0] mux_d0_62, next_mux_d0_62;
reg [0:0] mux_d0_63, next_mux_d0_63;
reg [0:0] mux_d0_64, next_mux_d0_64;
reg [0:0] mux_d0_65, next_mux_d0_65;
reg [0:0] mux_d0_66, next_mux_d0_66;
reg [0:0] mux_d0_67, next_mux_d0_67;
reg [0:0] mux_d0_68, next_mux_d0_68;
reg [0:0] mux_d0_69, next_mux_d0_69;
reg [0:0] mux_d0_70, next_mux_d0_70;
reg [0:0] mux_d0_71, next_mux_d0_71;
reg [0:0] mux_d0_72, next_mux_d0_72;
reg [0:0] mux_d0_73, next_mux_d0_73;
reg [0:0] mux_d0_74, next_mux_d0_74;
reg [0:0] mux_d0_75, next_mux_d0_75;
reg [0:0] mux_d0_76, next_mux_d0_76;
reg [0:0] mux_d0_77, next_mux_d0_77;
reg [0:0] mux_d0_78, next_mux_d0_78;
reg [0:0] mux_d0_79, next_mux_d0_79;
reg [0:0] mux_d0_80, next_mux_d0_80;
reg [0:0] mux_d0_81, next_mux_d0_81;
reg [0:0] mux_d0_82, next_mux_d0_82;
reg [0:0] mux_d0_83, next_mux_d0_83;
reg [0:0] mux_d0_84, next_mux_d0_84;
reg [0:0] mux_d0_85, next_mux_d0_85;
reg [0:0] mux_d0_86, next_mux_d0_86;
reg [0:0] mux_d0_87, next_mux_d0_87;
reg [0:0] mux_d0_88, next_mux_d0_88;
reg [0:0] mux_d0_89, next_mux_d0_89;
reg [0:0] mux_d0_90, next_mux_d0_90;
reg [0:0] mux_d0_91, next_mux_d0_91;
reg [0:0] mux_d0_92, next_mux_d0_92;
reg [0:0] mux_d0_93, next_mux_d0_93;
reg [0:0] mux_d0_94, next_mux_d0_94;
reg [0:0] mux_d0_95, next_mux_d0_95;
reg [0:0] mux_d0_96, next_mux_d0_96;
reg [0:0] mux_d0_97, next_mux_d0_97;
reg [0:0] mux_d0_98, next_mux_d0_98;
reg [0:0] mux_d0_99, next_mux_d0_99;
reg [0:0] mux_d0_100, next_mux_d0_100;
reg [0:0] mux_d0_101, next_mux_d0_101;
reg [0:0] mux_d0_102, next_mux_d0_102;
reg [0:0] mux_d0_103, next_mux_d0_103;
reg [0:0] mux_d0_104, next_mux_d0_104;
reg [0:0] mux_d0_105, next_mux_d0_105;
reg [0:0] mux_d0_106, next_mux_d0_106;
reg [0:0] mux_d0_107, next_mux_d0_107;
reg [0:0] mux_d0_108, next_mux_d0_108;
reg [0:0] mux_d0_109, next_mux_d0_109;
reg [0:0] mux_d0_110, next_mux_d0_110;
reg [0:0] mux_d0_111, next_mux_d0_111;
reg [0:0] mux_d0_112, next_mux_d0_112;
reg [0:0] mux_d0_113, next_mux_d0_113;
reg [0:0] mux_d0_114, next_mux_d0_114;
reg [0:0] mux_d0_115, next_mux_d0_115;
reg [0:0] mux_d0_116, next_mux_d0_116;
reg [0:0] mux_d0_117, next_mux_d0_117;
reg [0:0] mux_d0_118, next_mux_d0_118;
reg [0:0] mux_d0_119, next_mux_d0_119;
reg [0:0] mux_d0_120, next_mux_d0_120;
reg [0:0] mux_d0_121, next_mux_d0_121;
reg [0:0] mux_d0_122, next_mux_d0_122;
reg [0:0] mux_d0_123, next_mux_d0_123;
reg [0:0] mux_d0_124, next_mux_d0_124;
reg [0:0] mux_d0_125, next_mux_d0_125;
reg [0:0] mux_d0_126, next_mux_d0_126;
reg [0:0] mux_d0_127, next_mux_d0_127;
reg [0:0] mux_d0_128, next_mux_d0_128;
reg [0:0] mux_d0_129, next_mux_d0_129;
reg [0:0] mux_d0_130, next_mux_d0_130;
reg [0:0] mux_d0_131, next_mux_d0_131;
reg [0:0] mux_d0_132, next_mux_d0_132;
reg [0:0] mux_d0_133, next_mux_d0_133;
reg [0:0] mux_d0_134, next_mux_d0_134;
reg [0:0] mux_d0_135, next_mux_d0_135;
reg [0:0] mux_d0_136, next_mux_d0_136;
reg [0:0] mux_d0_137, next_mux_d0_137;
reg [0:0] mux_d0_138, next_mux_d0_138;
reg [0:0] mux_d0_139, next_mux_d0_139;
reg [0:0] mux_d0_140, next_mux_d0_140;
reg [0:0] mux_d0_141, next_mux_d0_141;
reg [0:0] mux_d0_142, next_mux_d0_142;
reg [0:0] mux_d0_143, next_mux_d0_143;
reg [0:0] mux_d0_144, next_mux_d0_144;
reg [0:0] mux_d0_145, next_mux_d0_145;
reg [0:0] mux_d0_146, next_mux_d0_146;
reg [0:0] mux_d0_147, next_mux_d0_147;
reg [0:0] mux_d0_148, next_mux_d0_148;
reg [0:0] mux_d0_149, next_mux_d0_149;
reg [0:0] mux_d0_150, next_mux_d0_150;
reg [0:0] mux_d0_151, next_mux_d0_151;
reg [0:0] mux_d0_152, next_mux_d0_152;
reg [0:0] mux_d0_153, next_mux_d0_153;
reg [0:0] mux_d0_154, next_mux_d0_154;
reg [0:0] mux_d0_155, next_mux_d0_155;
reg [0:0] mux_d0_156, next_mux_d0_156;
reg [0:0] mux_d0_157, next_mux_d0_157;
reg [0:0] mux_d0_158, next_mux_d0_158;
reg [0:0] mux_d0_159, next_mux_d0_159;
reg [0:0] mux_d0_160, next_mux_d0_160;
reg [0:0] mux_d0_161, next_mux_d0_161;
reg [0:0] mux_d0_162, next_mux_d0_162;
reg [0:0] mux_d0_163, next_mux_d0_163;
reg [0:0] mux_d0_164, next_mux_d0_164;
reg [0:0] mux_d0_165, next_mux_d0_165;
reg [0:0] mux_d0_166, next_mux_d0_166;
reg [0:0] mux_d0_167, next_mux_d0_167;
reg [0:0] mux_d0_168, next_mux_d0_168;
reg [0:0] mux_d0_169, next_mux_d0_169;
reg [0:0] mux_d0_170, next_mux_d0_170;
reg [0:0] mux_d0_171, next_mux_d0_171;
reg [0:0] mux_d0_172, next_mux_d0_172;
reg [0:0] mux_d0_173, next_mux_d0_173;
reg [0:0] mux_d0_174, next_mux_d0_174;
reg [0:0] mux_d0_175, next_mux_d0_175;
reg [0:0] mux_d0_176, next_mux_d0_176;
reg [0:0] mux_d0_177, next_mux_d0_177;
reg [0:0] mux_d0_178, next_mux_d0_178;
reg [0:0] mux_d0_179, next_mux_d0_179;
reg [0:0] mux_d0_180, next_mux_d0_180;
reg [0:0] mux_d0_181, next_mux_d0_181;
reg [0:0] mux_d0_182, next_mux_d0_182;
reg [0:0] mux_d0_183, next_mux_d0_183;
reg [0:0] mux_d0_184, next_mux_d0_184;
reg [0:0] mux_d0_185, next_mux_d0_185;
reg [0:0] mux_d0_186, next_mux_d0_186;
reg [0:0] mux_d0_187, next_mux_d0_187;
reg [0:0] mux_d0_188, next_mux_d0_188;
reg [0:0] mux_d0_189, next_mux_d0_189;
reg [0:0] mux_d0_190, next_mux_d0_190;
reg [0:0] mux_d0_191, next_mux_d0_191;
reg [0:0] mux_d0_192, next_mux_d0_192;
reg [0:0] mux_d0_193, next_mux_d0_193;
reg [0:0] mux_d0_194, next_mux_d0_194;
reg [0:0] mux_d0_195, next_mux_d0_195;
reg [0:0] mux_d0_196, next_mux_d0_196;
reg [0:0] mux_d0_197, next_mux_d0_197;
reg [0:0] mux_d0_198, next_mux_d0_198;
reg [0:0] mux_d0_199, next_mux_d0_199;
reg [0:0] mux_d0_200, next_mux_d0_200;
reg [0:0] mux_d0_201, next_mux_d0_201;
reg [0:0] mux_d0_202, next_mux_d0_202;
reg [0:0] mux_d0_203, next_mux_d0_203;
reg [0:0] mux_d0_204, next_mux_d0_204;
reg [0:0] mux_d0_205, next_mux_d0_205;
reg [0:0] mux_d0_206, next_mux_d0_206;
reg [0:0] mux_d0_207, next_mux_d0_207;
reg [0:0] mux_d0_208, next_mux_d0_208;
reg [0:0] mux_d0_209, next_mux_d0_209;
reg [0:0] mux_d0_210, next_mux_d0_210;
reg [0:0] mux_d0_211, next_mux_d0_211;
reg [0:0] mux_d0_212, next_mux_d0_212;
reg [0:0] mux_d0_213, next_mux_d0_213;
reg [0:0] mux_d0_214, next_mux_d0_214;
reg [0:0] mux_d0_215, next_mux_d0_215;
reg [0:0] mux_d0_216, next_mux_d0_216;
reg [0:0] mux_d0_217, next_mux_d0_217;
reg [0:0] mux_d0_218, next_mux_d0_218;
reg [0:0] mux_d0_219, next_mux_d0_219;
reg [0:0] mux_d0_220, next_mux_d0_220;
reg [0:0] mux_d0_221, next_mux_d0_221;
reg [0:0] mux_d0_222, next_mux_d0_222;
reg [0:0] mux_d0_223, next_mux_d0_223;
reg [0:0] mux_d0_224, next_mux_d0_224;
reg [0:0] mux_d0_225, next_mux_d0_225;
reg [0:0] mux_d0_226, next_mux_d0_226;
reg [0:0] mux_d0_227, next_mux_d0_227;
reg [0:0] mux_d0_228, next_mux_d0_228;
reg [0:0] mux_d0_229, next_mux_d0_229;
reg [0:0] mux_d0_230, next_mux_d0_230;
reg [0:0] mux_d0_231, next_mux_d0_231;
reg [0:0] mux_d0_232, next_mux_d0_232;
reg [0:0] mux_d0_233, next_mux_d0_233;
reg [0:0] mux_d0_234, next_mux_d0_234;
reg [0:0] mux_d0_235, next_mux_d0_235;
reg [0:0] mux_d0_236, next_mux_d0_236;
reg [0:0] mux_d0_237, next_mux_d0_237;
reg [0:0] mux_d0_238, next_mux_d0_238;
reg [0:0] mux_d0_239, next_mux_d0_239;
reg [0:0] mux_d0_240, next_mux_d0_240;
reg [0:0] mux_d0_241, next_mux_d0_241;
reg [0:0] mux_d0_242, next_mux_d0_242;
reg [0:0] mux_d0_243, next_mux_d0_243;
reg [0:0] mux_d0_244, next_mux_d0_244;
reg [0:0] mux_d0_245, next_mux_d0_245;
reg [0:0] mux_d0_246, next_mux_d0_246;
reg [0:0] mux_d0_247, next_mux_d0_247;
reg [0:0] mux_d0_248, next_mux_d0_248;
reg [0:0] mux_d0_249, next_mux_d0_249;
reg [0:0] mux_d0_250, next_mux_d0_250;
reg [0:0] mux_d0_251, next_mux_d0_251;
reg [0:0] mux_d0_252, next_mux_d0_252;
reg [0:0] mux_d0_253, next_mux_d0_253;
reg [0:0] mux_d0_254, next_mux_d0_254;
reg [0:0] mux_d0_255, next_mux_d0_255;
reg [0:0] mux_d1_0, next_mux_d1_0;
reg [0:0] mux_d1_1, next_mux_d1_1;
reg [0:0] mux_d1_2, next_mux_d1_2;
reg [0:0] mux_d1_3, next_mux_d1_3;
reg [0:0] mux_d1_4, next_mux_d1_4;
reg [0:0] mux_d1_5, next_mux_d1_5;
reg [0:0] mux_d1_6, next_mux_d1_6;
reg [0:0] mux_d1_7, next_mux_d1_7;
reg [0:0] mux_d1_8, next_mux_d1_8;
reg [0:0] mux_d1_9, next_mux_d1_9;
reg [0:0] mux_d1_10, next_mux_d1_10;
reg [0:0] mux_d1_11, next_mux_d1_11;
reg [0:0] mux_d1_12, next_mux_d1_12;
reg [0:0] mux_d1_13, next_mux_d1_13;
reg [0:0] mux_d1_14, next_mux_d1_14;
reg [0:0] mux_d1_15, next_mux_d1_15;
reg [0:0] mux_d1_16, next_mux_d1_16;
reg [0:0] mux_d1_17, next_mux_d1_17;
reg [0:0] mux_d1_18, next_mux_d1_18;
reg [0:0] mux_d1_19, next_mux_d1_19;
reg [0:0] mux_d1_20, next_mux_d1_20;
reg [0:0] mux_d1_21, next_mux_d1_21;
reg [0:0] mux_d1_22, next_mux_d1_22;
reg [0:0] mux_d1_23, next_mux_d1_23;
reg [0:0] mux_d1_24, next_mux_d1_24;
reg [0:0] mux_d1_25, next_mux_d1_25;
reg [0:0] mux_d1_26, next_mux_d1_26;
reg [0:0] mux_d1_27, next_mux_d1_27;
reg [0:0] mux_d1_28, next_mux_d1_28;
reg [0:0] mux_d1_29, next_mux_d1_29;
reg [0:0] mux_d1_30, next_mux_d1_30;
reg [0:0] mux_d1_31, next_mux_d1_31;
reg [0:0] mux_d2_0, next_mux_d2_0;
reg [0:0] mux_d2_1, next_mux_d2_1;
reg [0:0] mux_d2_2, next_mux_d2_2;
reg [0:0] mux_d2_3, next_mux_d2_3;
reg [0:0] mux_d3_0, next_mux_d3_0;
reg [2047:0] input_word_d;

assign output_word = mux_d3_0;
assign valid_o = valid_d4;
assign sel_o = sel_d4;

integer ii;

always @(posedge clk) begin
    if (sync_reset) begin
        valid_d0  <= 0;
        valid_d1  <= 0;
        valid_d2  <= 0;
        valid_d3  <= 0;
        valid_d4  <= 0;
    end else begin
        valid_d0  <= valid_i;
        valid_d1  <= valid_d0;
        valid_d2  <= valid_d1;
        valid_d3  <= valid_d2;
        valid_d4  <= valid_d3;
    end
end


always @(posedge clk) begin
    input_word_d <= input_word;
    mux_d0_0 <= next_mux_d0_0;
    mux_d0_1 <= next_mux_d0_1;
    mux_d0_2 <= next_mux_d0_2;
    mux_d0_3 <= next_mux_d0_3;
    mux_d0_4 <= next_mux_d0_4;
    mux_d0_5 <= next_mux_d0_5;
    mux_d0_6 <= next_mux_d0_6;
    mux_d0_7 <= next_mux_d0_7;
    mux_d0_8 <= next_mux_d0_8;
    mux_d0_9 <= next_mux_d0_9;
    mux_d0_10 <= next_mux_d0_10;
    mux_d0_11 <= next_mux_d0_11;
    mux_d0_12 <= next_mux_d0_12;
    mux_d0_13 <= next_mux_d0_13;
    mux_d0_14 <= next_mux_d0_14;
    mux_d0_15 <= next_mux_d0_15;
    mux_d0_16 <= next_mux_d0_16;
    mux_d0_17 <= next_mux_d0_17;
    mux_d0_18 <= next_mux_d0_18;
    mux_d0_19 <= next_mux_d0_19;
    mux_d0_20 <= next_mux_d0_20;
    mux_d0_21 <= next_mux_d0_21;
    mux_d0_22 <= next_mux_d0_22;
    mux_d0_23 <= next_mux_d0_23;
    mux_d0_24 <= next_mux_d0_24;
    mux_d0_25 <= next_mux_d0_25;
    mux_d0_26 <= next_mux_d0_26;
    mux_d0_27 <= next_mux_d0_27;
    mux_d0_28 <= next_mux_d0_28;
    mux_d0_29 <= next_mux_d0_29;
    mux_d0_30 <= next_mux_d0_30;
    mux_d0_31 <= next_mux_d0_31;
    mux_d0_32 <= next_mux_d0_32;
    mux_d0_33 <= next_mux_d0_33;
    mux_d0_34 <= next_mux_d0_34;
    mux_d0_35 <= next_mux_d0_35;
    mux_d0_36 <= next_mux_d0_36;
    mux_d0_37 <= next_mux_d0_37;
    mux_d0_38 <= next_mux_d0_38;
    mux_d0_39 <= next_mux_d0_39;
    mux_d0_40 <= next_mux_d0_40;
    mux_d0_41 <= next_mux_d0_41;
    mux_d0_42 <= next_mux_d0_42;
    mux_d0_43 <= next_mux_d0_43;
    mux_d0_44 <= next_mux_d0_44;
    mux_d0_45 <= next_mux_d0_45;
    mux_d0_46 <= next_mux_d0_46;
    mux_d0_47 <= next_mux_d0_47;
    mux_d0_48 <= next_mux_d0_48;
    mux_d0_49 <= next_mux_d0_49;
    mux_d0_50 <= next_mux_d0_50;
    mux_d0_51 <= next_mux_d0_51;
    mux_d0_52 <= next_mux_d0_52;
    mux_d0_53 <= next_mux_d0_53;
    mux_d0_54 <= next_mux_d0_54;
    mux_d0_55 <= next_mux_d0_55;
    mux_d0_56 <= next_mux_d0_56;
    mux_d0_57 <= next_mux_d0_57;
    mux_d0_58 <= next_mux_d0_58;
    mux_d0_59 <= next_mux_d0_59;
    mux_d0_60 <= next_mux_d0_60;
    mux_d0_61 <= next_mux_d0_61;
    mux_d0_62 <= next_mux_d0_62;
    mux_d0_63 <= next_mux_d0_63;
    mux_d0_64 <= next_mux_d0_64;
    mux_d0_65 <= next_mux_d0_65;
    mux_d0_66 <= next_mux_d0_66;
    mux_d0_67 <= next_mux_d0_67;
    mux_d0_68 <= next_mux_d0_68;
    mux_d0_69 <= next_mux_d0_69;
    mux_d0_70 <= next_mux_d0_70;
    mux_d0_71 <= next_mux_d0_71;
    mux_d0_72 <= next_mux_d0_72;
    mux_d0_73 <= next_mux_d0_73;
    mux_d0_74 <= next_mux_d0_74;
    mux_d0_75 <= next_mux_d0_75;
    mux_d0_76 <= next_mux_d0_76;
    mux_d0_77 <= next_mux_d0_77;
    mux_d0_78 <= next_mux_d0_78;
    mux_d0_79 <= next_mux_d0_79;
    mux_d0_80 <= next_mux_d0_80;
    mux_d0_81 <= next_mux_d0_81;
    mux_d0_82 <= next_mux_d0_82;
    mux_d0_83 <= next_mux_d0_83;
    mux_d0_84 <= next_mux_d0_84;
    mux_d0_85 <= next_mux_d0_85;
    mux_d0_86 <= next_mux_d0_86;
    mux_d0_87 <= next_mux_d0_87;
    mux_d0_88 <= next_mux_d0_88;
    mux_d0_89 <= next_mux_d0_89;
    mux_d0_90 <= next_mux_d0_90;
    mux_d0_91 <= next_mux_d0_91;
    mux_d0_92 <= next_mux_d0_92;
    mux_d0_93 <= next_mux_d0_93;
    mux_d0_94 <= next_mux_d0_94;
    mux_d0_95 <= next_mux_d0_95;
    mux_d0_96 <= next_mux_d0_96;
    mux_d0_97 <= next_mux_d0_97;
    mux_d0_98 <= next_mux_d0_98;
    mux_d0_99 <= next_mux_d0_99;
    mux_d0_100 <= next_mux_d0_100;
    mux_d0_101 <= next_mux_d0_101;
    mux_d0_102 <= next_mux_d0_102;
    mux_d0_103 <= next_mux_d0_103;
    mux_d0_104 <= next_mux_d0_104;
    mux_d0_105 <= next_mux_d0_105;
    mux_d0_106 <= next_mux_d0_106;
    mux_d0_107 <= next_mux_d0_107;
    mux_d0_108 <= next_mux_d0_108;
    mux_d0_109 <= next_mux_d0_109;
    mux_d0_110 <= next_mux_d0_110;
    mux_d0_111 <= next_mux_d0_111;
    mux_d0_112 <= next_mux_d0_112;
    mux_d0_113 <= next_mux_d0_113;
    mux_d0_114 <= next_mux_d0_114;
    mux_d0_115 <= next_mux_d0_115;
    mux_d0_116 <= next_mux_d0_116;
    mux_d0_117 <= next_mux_d0_117;
    mux_d0_118 <= next_mux_d0_118;
    mux_d0_119 <= next_mux_d0_119;
    mux_d0_120 <= next_mux_d0_120;
    mux_d0_121 <= next_mux_d0_121;
    mux_d0_122 <= next_mux_d0_122;
    mux_d0_123 <= next_mux_d0_123;
    mux_d0_124 <= next_mux_d0_124;
    mux_d0_125 <= next_mux_d0_125;
    mux_d0_126 <= next_mux_d0_126;
    mux_d0_127 <= next_mux_d0_127;
    mux_d0_128 <= next_mux_d0_128;
    mux_d0_129 <= next_mux_d0_129;
    mux_d0_130 <= next_mux_d0_130;
    mux_d0_131 <= next_mux_d0_131;
    mux_d0_132 <= next_mux_d0_132;
    mux_d0_133 <= next_mux_d0_133;
    mux_d0_134 <= next_mux_d0_134;
    mux_d0_135 <= next_mux_d0_135;
    mux_d0_136 <= next_mux_d0_136;
    mux_d0_137 <= next_mux_d0_137;
    mux_d0_138 <= next_mux_d0_138;
    mux_d0_139 <= next_mux_d0_139;
    mux_d0_140 <= next_mux_d0_140;
    mux_d0_141 <= next_mux_d0_141;
    mux_d0_142 <= next_mux_d0_142;
    mux_d0_143 <= next_mux_d0_143;
    mux_d0_144 <= next_mux_d0_144;
    mux_d0_145 <= next_mux_d0_145;
    mux_d0_146 <= next_mux_d0_146;
    mux_d0_147 <= next_mux_d0_147;
    mux_d0_148 <= next_mux_d0_148;
    mux_d0_149 <= next_mux_d0_149;
    mux_d0_150 <= next_mux_d0_150;
    mux_d0_151 <= next_mux_d0_151;
    mux_d0_152 <= next_mux_d0_152;
    mux_d0_153 <= next_mux_d0_153;
    mux_d0_154 <= next_mux_d0_154;
    mux_d0_155 <= next_mux_d0_155;
    mux_d0_156 <= next_mux_d0_156;
    mux_d0_157 <= next_mux_d0_157;
    mux_d0_158 <= next_mux_d0_158;
    mux_d0_159 <= next_mux_d0_159;
    mux_d0_160 <= next_mux_d0_160;
    mux_d0_161 <= next_mux_d0_161;
    mux_d0_162 <= next_mux_d0_162;
    mux_d0_163 <= next_mux_d0_163;
    mux_d0_164 <= next_mux_d0_164;
    mux_d0_165 <= next_mux_d0_165;
    mux_d0_166 <= next_mux_d0_166;
    mux_d0_167 <= next_mux_d0_167;
    mux_d0_168 <= next_mux_d0_168;
    mux_d0_169 <= next_mux_d0_169;
    mux_d0_170 <= next_mux_d0_170;
    mux_d0_171 <= next_mux_d0_171;
    mux_d0_172 <= next_mux_d0_172;
    mux_d0_173 <= next_mux_d0_173;
    mux_d0_174 <= next_mux_d0_174;
    mux_d0_175 <= next_mux_d0_175;
    mux_d0_176 <= next_mux_d0_176;
    mux_d0_177 <= next_mux_d0_177;
    mux_d0_178 <= next_mux_d0_178;
    mux_d0_179 <= next_mux_d0_179;
    mux_d0_180 <= next_mux_d0_180;
    mux_d0_181 <= next_mux_d0_181;
    mux_d0_182 <= next_mux_d0_182;
    mux_d0_183 <= next_mux_d0_183;
    mux_d0_184 <= next_mux_d0_184;
    mux_d0_185 <= next_mux_d0_185;
    mux_d0_186 <= next_mux_d0_186;
    mux_d0_187 <= next_mux_d0_187;
    mux_d0_188 <= next_mux_d0_188;
    mux_d0_189 <= next_mux_d0_189;
    mux_d0_190 <= next_mux_d0_190;
    mux_d0_191 <= next_mux_d0_191;
    mux_d0_192 <= next_mux_d0_192;
    mux_d0_193 <= next_mux_d0_193;
    mux_d0_194 <= next_mux_d0_194;
    mux_d0_195 <= next_mux_d0_195;
    mux_d0_196 <= next_mux_d0_196;
    mux_d0_197 <= next_mux_d0_197;
    mux_d0_198 <= next_mux_d0_198;
    mux_d0_199 <= next_mux_d0_199;
    mux_d0_200 <= next_mux_d0_200;
    mux_d0_201 <= next_mux_d0_201;
    mux_d0_202 <= next_mux_d0_202;
    mux_d0_203 <= next_mux_d0_203;
    mux_d0_204 <= next_mux_d0_204;
    mux_d0_205 <= next_mux_d0_205;
    mux_d0_206 <= next_mux_d0_206;
    mux_d0_207 <= next_mux_d0_207;
    mux_d0_208 <= next_mux_d0_208;
    mux_d0_209 <= next_mux_d0_209;
    mux_d0_210 <= next_mux_d0_210;
    mux_d0_211 <= next_mux_d0_211;
    mux_d0_212 <= next_mux_d0_212;
    mux_d0_213 <= next_mux_d0_213;
    mux_d0_214 <= next_mux_d0_214;
    mux_d0_215 <= next_mux_d0_215;
    mux_d0_216 <= next_mux_d0_216;
    mux_d0_217 <= next_mux_d0_217;
    mux_d0_218 <= next_mux_d0_218;
    mux_d0_219 <= next_mux_d0_219;
    mux_d0_220 <= next_mux_d0_220;
    mux_d0_221 <= next_mux_d0_221;
    mux_d0_222 <= next_mux_d0_222;
    mux_d0_223 <= next_mux_d0_223;
    mux_d0_224 <= next_mux_d0_224;
    mux_d0_225 <= next_mux_d0_225;
    mux_d0_226 <= next_mux_d0_226;
    mux_d0_227 <= next_mux_d0_227;
    mux_d0_228 <= next_mux_d0_228;
    mux_d0_229 <= next_mux_d0_229;
    mux_d0_230 <= next_mux_d0_230;
    mux_d0_231 <= next_mux_d0_231;
    mux_d0_232 <= next_mux_d0_232;
    mux_d0_233 <= next_mux_d0_233;
    mux_d0_234 <= next_mux_d0_234;
    mux_d0_235 <= next_mux_d0_235;
    mux_d0_236 <= next_mux_d0_236;
    mux_d0_237 <= next_mux_d0_237;
    mux_d0_238 <= next_mux_d0_238;
    mux_d0_239 <= next_mux_d0_239;
    mux_d0_240 <= next_mux_d0_240;
    mux_d0_241 <= next_mux_d0_241;
    mux_d0_242 <= next_mux_d0_242;
    mux_d0_243 <= next_mux_d0_243;
    mux_d0_244 <= next_mux_d0_244;
    mux_d0_245 <= next_mux_d0_245;
    mux_d0_246 <= next_mux_d0_246;
    mux_d0_247 <= next_mux_d0_247;
    mux_d0_248 <= next_mux_d0_248;
    mux_d0_249 <= next_mux_d0_249;
    mux_d0_250 <= next_mux_d0_250;
    mux_d0_251 <= next_mux_d0_251;
    mux_d0_252 <= next_mux_d0_252;
    mux_d0_253 <= next_mux_d0_253;
    mux_d0_254 <= next_mux_d0_254;
    mux_d0_255 <= next_mux_d0_255;
    mux_d1_0 <= next_mux_d1_0;
    mux_d1_1 <= next_mux_d1_1;
    mux_d1_2 <= next_mux_d1_2;
    mux_d1_3 <= next_mux_d1_3;
    mux_d1_4 <= next_mux_d1_4;
    mux_d1_5 <= next_mux_d1_5;
    mux_d1_6 <= next_mux_d1_6;
    mux_d1_7 <= next_mux_d1_7;
    mux_d1_8 <= next_mux_d1_8;
    mux_d1_9 <= next_mux_d1_9;
    mux_d1_10 <= next_mux_d1_10;
    mux_d1_11 <= next_mux_d1_11;
    mux_d1_12 <= next_mux_d1_12;
    mux_d1_13 <= next_mux_d1_13;
    mux_d1_14 <= next_mux_d1_14;
    mux_d1_15 <= next_mux_d1_15;
    mux_d1_16 <= next_mux_d1_16;
    mux_d1_17 <= next_mux_d1_17;
    mux_d1_18 <= next_mux_d1_18;
    mux_d1_19 <= next_mux_d1_19;
    mux_d1_20 <= next_mux_d1_20;
    mux_d1_21 <= next_mux_d1_21;
    mux_d1_22 <= next_mux_d1_22;
    mux_d1_23 <= next_mux_d1_23;
    mux_d1_24 <= next_mux_d1_24;
    mux_d1_25 <= next_mux_d1_25;
    mux_d1_26 <= next_mux_d1_26;
    mux_d1_27 <= next_mux_d1_27;
    mux_d1_28 <= next_mux_d1_28;
    mux_d1_29 <= next_mux_d1_29;
    mux_d1_30 <= next_mux_d1_30;
    mux_d1_31 <= next_mux_d1_31;
    mux_d2_0 <= next_mux_d2_0;
    mux_d2_1 <= next_mux_d2_1;
    mux_d2_2 <= next_mux_d2_2;
    mux_d2_3 <= next_mux_d2_3;
    mux_d3_0 <= next_mux_d3_0;
    sel_d0_0 <= sel;
    sel_d0_1 <= sel;
    sel_d0_2 <= sel;
    sel_d0_3 <= sel;
    sel_d0_4 <= sel;
    sel_d0_5 <= sel;
    sel_d0_6 <= sel;
    sel_d0_7 <= sel;
    sel_d0_8 <= sel;
    sel_d0_9 <= sel;
    sel_d0_10 <= sel;
    sel_d0_11 <= sel;
    sel_d0_12 <= sel;
    sel_d0_13 <= sel;
    sel_d0_14 <= sel;
    sel_d0_15 <= sel;
    sel_d0_16 <= sel;
    sel_d0_17 <= sel;
    sel_d0_18 <= sel;
    sel_d0_19 <= sel;
    sel_d0_20 <= sel;
    sel_d0_21 <= sel;
    sel_d0_22 <= sel;
    sel_d0_23 <= sel;
    sel_d0_24 <= sel;
    sel_d0_25 <= sel;
    sel_d0_26 <= sel;
    sel_d0_27 <= sel;
    sel_d0_28 <= sel;
    sel_d0_29 <= sel;
    sel_d0_30 <= sel;
    sel_d0_31 <= sel;
    sel_d0_32 <= sel;
    sel_d0_33 <= sel;
    sel_d0_34 <= sel;
    sel_d0_35 <= sel;
    sel_d0_36 <= sel;
    sel_d0_37 <= sel;
    sel_d0_38 <= sel;
    sel_d0_39 <= sel;
    sel_d0_40 <= sel;
    sel_d0_41 <= sel;
    sel_d0_42 <= sel;
    sel_d0_43 <= sel;
    sel_d0_44 <= sel;
    sel_d0_45 <= sel;
    sel_d0_46 <= sel;
    sel_d0_47 <= sel;
    sel_d0_48 <= sel;
    sel_d0_49 <= sel;
    sel_d0_50 <= sel;
    sel_d0_51 <= sel;
    sel_d0_52 <= sel;
    sel_d0_53 <= sel;
    sel_d0_54 <= sel;
    sel_d0_55 <= sel;
    sel_d0_56 <= sel;
    sel_d0_57 <= sel;
    sel_d0_58 <= sel;
    sel_d0_59 <= sel;
    sel_d0_60 <= sel;
    sel_d0_61 <= sel;
    sel_d0_62 <= sel;
    sel_d0_63 <= sel;
    sel_d0_64 <= sel;
    sel_d0_65 <= sel;
    sel_d0_66 <= sel;
    sel_d0_67 <= sel;
    sel_d0_68 <= sel;
    sel_d0_69 <= sel;
    sel_d0_70 <= sel;
    sel_d0_71 <= sel;
    sel_d0_72 <= sel;
    sel_d0_73 <= sel;
    sel_d0_74 <= sel;
    sel_d0_75 <= sel;
    sel_d0_76 <= sel;
    sel_d0_77 <= sel;
    sel_d0_78 <= sel;
    sel_d0_79 <= sel;
    sel_d0_80 <= sel;
    sel_d0_81 <= sel;
    sel_d0_82 <= sel;
    sel_d0_83 <= sel;
    sel_d0_84 <= sel;
    sel_d0_85 <= sel;
    sel_d0_86 <= sel;
    sel_d0_87 <= sel;
    sel_d0_88 <= sel;
    sel_d0_89 <= sel;
    sel_d0_90 <= sel;
    sel_d0_91 <= sel;
    sel_d0_92 <= sel;
    sel_d0_93 <= sel;
    sel_d0_94 <= sel;
    sel_d0_95 <= sel;
    sel_d0_96 <= sel;
    sel_d0_97 <= sel;
    sel_d0_98 <= sel;
    sel_d0_99 <= sel;
    sel_d0_100 <= sel;
    sel_d0_101 <= sel;
    sel_d0_102 <= sel;
    sel_d0_103 <= sel;
    sel_d0_104 <= sel;
    sel_d0_105 <= sel;
    sel_d0_106 <= sel;
    sel_d0_107 <= sel;
    sel_d0_108 <= sel;
    sel_d0_109 <= sel;
    sel_d0_110 <= sel;
    sel_d0_111 <= sel;
    sel_d0_112 <= sel;
    sel_d0_113 <= sel;
    sel_d0_114 <= sel;
    sel_d0_115 <= sel;
    sel_d0_116 <= sel;
    sel_d0_117 <= sel;
    sel_d0_118 <= sel;
    sel_d0_119 <= sel;
    sel_d0_120 <= sel;
    sel_d0_121 <= sel;
    sel_d0_122 <= sel;
    sel_d0_123 <= sel;
    sel_d0_124 <= sel;
    sel_d0_125 <= sel;
    sel_d0_126 <= sel;
    sel_d0_127 <= sel;
    sel_d0_128 <= sel;
    sel_d0_129 <= sel;
    sel_d0_130 <= sel;
    sel_d0_131 <= sel;
    sel_d0_132 <= sel;
    sel_d0_133 <= sel;
    sel_d0_134 <= sel;
    sel_d0_135 <= sel;
    sel_d0_136 <= sel;
    sel_d0_137 <= sel;
    sel_d0_138 <= sel;
    sel_d0_139 <= sel;
    sel_d0_140 <= sel;
    sel_d0_141 <= sel;
    sel_d0_142 <= sel;
    sel_d0_143 <= sel;
    sel_d0_144 <= sel;
    sel_d0_145 <= sel;
    sel_d0_146 <= sel;
    sel_d0_147 <= sel;
    sel_d0_148 <= sel;
    sel_d0_149 <= sel;
    sel_d0_150 <= sel;
    sel_d0_151 <= sel;
    sel_d0_152 <= sel;
    sel_d0_153 <= sel;
    sel_d0_154 <= sel;
    sel_d0_155 <= sel;
    sel_d0_156 <= sel;
    sel_d0_157 <= sel;
    sel_d0_158 <= sel;
    sel_d0_159 <= sel;
    sel_d0_160 <= sel;
    sel_d0_161 <= sel;
    sel_d0_162 <= sel;
    sel_d0_163 <= sel;
    sel_d0_164 <= sel;
    sel_d0_165 <= sel;
    sel_d0_166 <= sel;
    sel_d0_167 <= sel;
    sel_d0_168 <= sel;
    sel_d0_169 <= sel;
    sel_d0_170 <= sel;
    sel_d0_171 <= sel;
    sel_d0_172 <= sel;
    sel_d0_173 <= sel;
    sel_d0_174 <= sel;
    sel_d0_175 <= sel;
    sel_d0_176 <= sel;
    sel_d0_177 <= sel;
    sel_d0_178 <= sel;
    sel_d0_179 <= sel;
    sel_d0_180 <= sel;
    sel_d0_181 <= sel;
    sel_d0_182 <= sel;
    sel_d0_183 <= sel;
    sel_d0_184 <= sel;
    sel_d0_185 <= sel;
    sel_d0_186 <= sel;
    sel_d0_187 <= sel;
    sel_d0_188 <= sel;
    sel_d0_189 <= sel;
    sel_d0_190 <= sel;
    sel_d0_191 <= sel;
    sel_d0_192 <= sel;
    sel_d0_193 <= sel;
    sel_d0_194 <= sel;
    sel_d0_195 <= sel;
    sel_d0_196 <= sel;
    sel_d0_197 <= sel;
    sel_d0_198 <= sel;
    sel_d0_199 <= sel;
    sel_d0_200 <= sel;
    sel_d0_201 <= sel;
    sel_d0_202 <= sel;
    sel_d0_203 <= sel;
    sel_d0_204 <= sel;
    sel_d0_205 <= sel;
    sel_d0_206 <= sel;
    sel_d0_207 <= sel;
    sel_d0_208 <= sel;
    sel_d0_209 <= sel;
    sel_d0_210 <= sel;
    sel_d0_211 <= sel;
    sel_d0_212 <= sel;
    sel_d0_213 <= sel;
    sel_d0_214 <= sel;
    sel_d0_215 <= sel;
    sel_d0_216 <= sel;
    sel_d0_217 <= sel;
    sel_d0_218 <= sel;
    sel_d0_219 <= sel;
    sel_d0_220 <= sel;
    sel_d0_221 <= sel;
    sel_d0_222 <= sel;
    sel_d0_223 <= sel;
    sel_d0_224 <= sel;
    sel_d0_225 <= sel;
    sel_d0_226 <= sel;
    sel_d0_227 <= sel;
    sel_d0_228 <= sel;
    sel_d0_229 <= sel;
    sel_d0_230 <= sel;
    sel_d0_231 <= sel;
    sel_d0_232 <= sel;
    sel_d0_233 <= sel;
    sel_d0_234 <= sel;
    sel_d0_235 <= sel;
    sel_d0_236 <= sel;
    sel_d0_237 <= sel;
    sel_d0_238 <= sel;
    sel_d0_239 <= sel;
    sel_d0_240 <= sel;
    sel_d0_241 <= sel;
    sel_d0_242 <= sel;
    sel_d0_243 <= sel;
    sel_d0_244 <= sel;
    sel_d0_245 <= sel;
    sel_d0_246 <= sel;
    sel_d0_247 <= sel;
    sel_d0_248 <= sel;
    sel_d0_249 <= sel;
    sel_d0_250 <= sel;
    sel_d0_251 <= sel;
    sel_d0_252 <= sel;
    sel_d0_253 <= sel;
    sel_d0_254 <= sel;
    sel_d0_255 <= sel;
    sel_d1_0 <= sel_d0_255;
    sel_d1_1 <= sel_d0_255;
    sel_d1_2 <= sel_d0_255;
    sel_d1_3 <= sel_d0_255;
    sel_d1_4 <= sel_d0_255;
    sel_d1_5 <= sel_d0_255;
    sel_d1_6 <= sel_d0_255;
    sel_d1_7 <= sel_d0_255;
    sel_d1_8 <= sel_d0_255;
    sel_d1_9 <= sel_d0_255;
    sel_d1_10 <= sel_d0_255;
    sel_d1_11 <= sel_d0_255;
    sel_d1_12 <= sel_d0_255;
    sel_d1_13 <= sel_d0_255;
    sel_d1_14 <= sel_d0_255;
    sel_d1_15 <= sel_d0_255;
    sel_d1_16 <= sel_d0_255;
    sel_d1_17 <= sel_d0_255;
    sel_d1_18 <= sel_d0_255;
    sel_d1_19 <= sel_d0_255;
    sel_d1_20 <= sel_d0_255;
    sel_d1_21 <= sel_d0_255;
    sel_d1_22 <= sel_d0_255;
    sel_d1_23 <= sel_d0_255;
    sel_d1_24 <= sel_d0_255;
    sel_d1_25 <= sel_d0_255;
    sel_d1_26 <= sel_d0_255;
    sel_d1_27 <= sel_d0_255;
    sel_d1_28 <= sel_d0_255;
    sel_d1_29 <= sel_d0_255;
    sel_d1_30 <= sel_d0_255;
    sel_d1_31 <= sel_d0_255;
    sel_d2_0 <= sel_d1_31;
    sel_d2_1 <= sel_d1_31;
    sel_d2_2 <= sel_d1_31;
    sel_d2_3 <= sel_d1_31;
    sel_d3_0 <= sel_d2_3;
    sel_d4 <= sel_d3_0;
end


always @*
begin
    next_mux_d0_0 = mux_d0_0;
    next_mux_d0_1 = mux_d0_1;
    next_mux_d0_2 = mux_d0_2;
    next_mux_d0_3 = mux_d0_3;
    next_mux_d0_4 = mux_d0_4;
    next_mux_d0_5 = mux_d0_5;
    next_mux_d0_6 = mux_d0_6;
    next_mux_d0_7 = mux_d0_7;
    next_mux_d0_8 = mux_d0_8;
    next_mux_d0_9 = mux_d0_9;
    next_mux_d0_10 = mux_d0_10;
    next_mux_d0_11 = mux_d0_11;
    next_mux_d0_12 = mux_d0_12;
    next_mux_d0_13 = mux_d0_13;
    next_mux_d0_14 = mux_d0_14;
    next_mux_d0_15 = mux_d0_15;
    next_mux_d0_16 = mux_d0_16;
    next_mux_d0_17 = mux_d0_17;
    next_mux_d0_18 = mux_d0_18;
    next_mux_d0_19 = mux_d0_19;
    next_mux_d0_20 = mux_d0_20;
    next_mux_d0_21 = mux_d0_21;
    next_mux_d0_22 = mux_d0_22;
    next_mux_d0_23 = mux_d0_23;
    next_mux_d0_24 = mux_d0_24;
    next_mux_d0_25 = mux_d0_25;
    next_mux_d0_26 = mux_d0_26;
    next_mux_d0_27 = mux_d0_27;
    next_mux_d0_28 = mux_d0_28;
    next_mux_d0_29 = mux_d0_29;
    next_mux_d0_30 = mux_d0_30;
    next_mux_d0_31 = mux_d0_31;
    next_mux_d0_32 = mux_d0_32;
    next_mux_d0_33 = mux_d0_33;
    next_mux_d0_34 = mux_d0_34;
    next_mux_d0_35 = mux_d0_35;
    next_mux_d0_36 = mux_d0_36;
    next_mux_d0_37 = mux_d0_37;
    next_mux_d0_38 = mux_d0_38;
    next_mux_d0_39 = mux_d0_39;
    next_mux_d0_40 = mux_d0_40;
    next_mux_d0_41 = mux_d0_41;
    next_mux_d0_42 = mux_d0_42;
    next_mux_d0_43 = mux_d0_43;
    next_mux_d0_44 = mux_d0_44;
    next_mux_d0_45 = mux_d0_45;
    next_mux_d0_46 = mux_d0_46;
    next_mux_d0_47 = mux_d0_47;
    next_mux_d0_48 = mux_d0_48;
    next_mux_d0_49 = mux_d0_49;
    next_mux_d0_50 = mux_d0_50;
    next_mux_d0_51 = mux_d0_51;
    next_mux_d0_52 = mux_d0_52;
    next_mux_d0_53 = mux_d0_53;
    next_mux_d0_54 = mux_d0_54;
    next_mux_d0_55 = mux_d0_55;
    next_mux_d0_56 = mux_d0_56;
    next_mux_d0_57 = mux_d0_57;
    next_mux_d0_58 = mux_d0_58;
    next_mux_d0_59 = mux_d0_59;
    next_mux_d0_60 = mux_d0_60;
    next_mux_d0_61 = mux_d0_61;
    next_mux_d0_62 = mux_d0_62;
    next_mux_d0_63 = mux_d0_63;
    next_mux_d0_64 = mux_d0_64;
    next_mux_d0_65 = mux_d0_65;
    next_mux_d0_66 = mux_d0_66;
    next_mux_d0_67 = mux_d0_67;
    next_mux_d0_68 = mux_d0_68;
    next_mux_d0_69 = mux_d0_69;
    next_mux_d0_70 = mux_d0_70;
    next_mux_d0_71 = mux_d0_71;
    next_mux_d0_72 = mux_d0_72;
    next_mux_d0_73 = mux_d0_73;
    next_mux_d0_74 = mux_d0_74;
    next_mux_d0_75 = mux_d0_75;
    next_mux_d0_76 = mux_d0_76;
    next_mux_d0_77 = mux_d0_77;
    next_mux_d0_78 = mux_d0_78;
    next_mux_d0_79 = mux_d0_79;
    next_mux_d0_80 = mux_d0_80;
    next_mux_d0_81 = mux_d0_81;
    next_mux_d0_82 = mux_d0_82;
    next_mux_d0_83 = mux_d0_83;
    next_mux_d0_84 = mux_d0_84;
    next_mux_d0_85 = mux_d0_85;
    next_mux_d0_86 = mux_d0_86;
    next_mux_d0_87 = mux_d0_87;
    next_mux_d0_88 = mux_d0_88;
    next_mux_d0_89 = mux_d0_89;
    next_mux_d0_90 = mux_d0_90;
    next_mux_d0_91 = mux_d0_91;
    next_mux_d0_92 = mux_d0_92;
    next_mux_d0_93 = mux_d0_93;
    next_mux_d0_94 = mux_d0_94;
    next_mux_d0_95 = mux_d0_95;
    next_mux_d0_96 = mux_d0_96;
    next_mux_d0_97 = mux_d0_97;
    next_mux_d0_98 = mux_d0_98;
    next_mux_d0_99 = mux_d0_99;
    next_mux_d0_100 = mux_d0_100;
    next_mux_d0_101 = mux_d0_101;
    next_mux_d0_102 = mux_d0_102;
    next_mux_d0_103 = mux_d0_103;
    next_mux_d0_104 = mux_d0_104;
    next_mux_d0_105 = mux_d0_105;
    next_mux_d0_106 = mux_d0_106;
    next_mux_d0_107 = mux_d0_107;
    next_mux_d0_108 = mux_d0_108;
    next_mux_d0_109 = mux_d0_109;
    next_mux_d0_110 = mux_d0_110;
    next_mux_d0_111 = mux_d0_111;
    next_mux_d0_112 = mux_d0_112;
    next_mux_d0_113 = mux_d0_113;
    next_mux_d0_114 = mux_d0_114;
    next_mux_d0_115 = mux_d0_115;
    next_mux_d0_116 = mux_d0_116;
    next_mux_d0_117 = mux_d0_117;
    next_mux_d0_118 = mux_d0_118;
    next_mux_d0_119 = mux_d0_119;
    next_mux_d0_120 = mux_d0_120;
    next_mux_d0_121 = mux_d0_121;
    next_mux_d0_122 = mux_d0_122;
    next_mux_d0_123 = mux_d0_123;
    next_mux_d0_124 = mux_d0_124;
    next_mux_d0_125 = mux_d0_125;
    next_mux_d0_126 = mux_d0_126;
    next_mux_d0_127 = mux_d0_127;
    next_mux_d0_128 = mux_d0_128;
    next_mux_d0_129 = mux_d0_129;
    next_mux_d0_130 = mux_d0_130;
    next_mux_d0_131 = mux_d0_131;
    next_mux_d0_132 = mux_d0_132;
    next_mux_d0_133 = mux_d0_133;
    next_mux_d0_134 = mux_d0_134;
    next_mux_d0_135 = mux_d0_135;
    next_mux_d0_136 = mux_d0_136;
    next_mux_d0_137 = mux_d0_137;
    next_mux_d0_138 = mux_d0_138;
    next_mux_d0_139 = mux_d0_139;
    next_mux_d0_140 = mux_d0_140;
    next_mux_d0_141 = mux_d0_141;
    next_mux_d0_142 = mux_d0_142;
    next_mux_d0_143 = mux_d0_143;
    next_mux_d0_144 = mux_d0_144;
    next_mux_d0_145 = mux_d0_145;
    next_mux_d0_146 = mux_d0_146;
    next_mux_d0_147 = mux_d0_147;
    next_mux_d0_148 = mux_d0_148;
    next_mux_d0_149 = mux_d0_149;
    next_mux_d0_150 = mux_d0_150;
    next_mux_d0_151 = mux_d0_151;
    next_mux_d0_152 = mux_d0_152;
    next_mux_d0_153 = mux_d0_153;
    next_mux_d0_154 = mux_d0_154;
    next_mux_d0_155 = mux_d0_155;
    next_mux_d0_156 = mux_d0_156;
    next_mux_d0_157 = mux_d0_157;
    next_mux_d0_158 = mux_d0_158;
    next_mux_d0_159 = mux_d0_159;
    next_mux_d0_160 = mux_d0_160;
    next_mux_d0_161 = mux_d0_161;
    next_mux_d0_162 = mux_d0_162;
    next_mux_d0_163 = mux_d0_163;
    next_mux_d0_164 = mux_d0_164;
    next_mux_d0_165 = mux_d0_165;
    next_mux_d0_166 = mux_d0_166;
    next_mux_d0_167 = mux_d0_167;
    next_mux_d0_168 = mux_d0_168;
    next_mux_d0_169 = mux_d0_169;
    next_mux_d0_170 = mux_d0_170;
    next_mux_d0_171 = mux_d0_171;
    next_mux_d0_172 = mux_d0_172;
    next_mux_d0_173 = mux_d0_173;
    next_mux_d0_174 = mux_d0_174;
    next_mux_d0_175 = mux_d0_175;
    next_mux_d0_176 = mux_d0_176;
    next_mux_d0_177 = mux_d0_177;
    next_mux_d0_178 = mux_d0_178;
    next_mux_d0_179 = mux_d0_179;
    next_mux_d0_180 = mux_d0_180;
    next_mux_d0_181 = mux_d0_181;
    next_mux_d0_182 = mux_d0_182;
    next_mux_d0_183 = mux_d0_183;
    next_mux_d0_184 = mux_d0_184;
    next_mux_d0_185 = mux_d0_185;
    next_mux_d0_186 = mux_d0_186;
    next_mux_d0_187 = mux_d0_187;
    next_mux_d0_188 = mux_d0_188;
    next_mux_d0_189 = mux_d0_189;
    next_mux_d0_190 = mux_d0_190;
    next_mux_d0_191 = mux_d0_191;
    next_mux_d0_192 = mux_d0_192;
    next_mux_d0_193 = mux_d0_193;
    next_mux_d0_194 = mux_d0_194;
    next_mux_d0_195 = mux_d0_195;
    next_mux_d0_196 = mux_d0_196;
    next_mux_d0_197 = mux_d0_197;
    next_mux_d0_198 = mux_d0_198;
    next_mux_d0_199 = mux_d0_199;
    next_mux_d0_200 = mux_d0_200;
    next_mux_d0_201 = mux_d0_201;
    next_mux_d0_202 = mux_d0_202;
    next_mux_d0_203 = mux_d0_203;
    next_mux_d0_204 = mux_d0_204;
    next_mux_d0_205 = mux_d0_205;
    next_mux_d0_206 = mux_d0_206;
    next_mux_d0_207 = mux_d0_207;
    next_mux_d0_208 = mux_d0_208;
    next_mux_d0_209 = mux_d0_209;
    next_mux_d0_210 = mux_d0_210;
    next_mux_d0_211 = mux_d0_211;
    next_mux_d0_212 = mux_d0_212;
    next_mux_d0_213 = mux_d0_213;
    next_mux_d0_214 = mux_d0_214;
    next_mux_d0_215 = mux_d0_215;
    next_mux_d0_216 = mux_d0_216;
    next_mux_d0_217 = mux_d0_217;
    next_mux_d0_218 = mux_d0_218;
    next_mux_d0_219 = mux_d0_219;
    next_mux_d0_220 = mux_d0_220;
    next_mux_d0_221 = mux_d0_221;
    next_mux_d0_222 = mux_d0_222;
    next_mux_d0_223 = mux_d0_223;
    next_mux_d0_224 = mux_d0_224;
    next_mux_d0_225 = mux_d0_225;
    next_mux_d0_226 = mux_d0_226;
    next_mux_d0_227 = mux_d0_227;
    next_mux_d0_228 = mux_d0_228;
    next_mux_d0_229 = mux_d0_229;
    next_mux_d0_230 = mux_d0_230;
    next_mux_d0_231 = mux_d0_231;
    next_mux_d0_232 = mux_d0_232;
    next_mux_d0_233 = mux_d0_233;
    next_mux_d0_234 = mux_d0_234;
    next_mux_d0_235 = mux_d0_235;
    next_mux_d0_236 = mux_d0_236;
    next_mux_d0_237 = mux_d0_237;
    next_mux_d0_238 = mux_d0_238;
    next_mux_d0_239 = mux_d0_239;
    next_mux_d0_240 = mux_d0_240;
    next_mux_d0_241 = mux_d0_241;
    next_mux_d0_242 = mux_d0_242;
    next_mux_d0_243 = mux_d0_243;
    next_mux_d0_244 = mux_d0_244;
    next_mux_d0_245 = mux_d0_245;
    next_mux_d0_246 = mux_d0_246;
    next_mux_d0_247 = mux_d0_247;
    next_mux_d0_248 = mux_d0_248;
    next_mux_d0_249 = mux_d0_249;
    next_mux_d0_250 = mux_d0_250;
    next_mux_d0_251 = mux_d0_251;
    next_mux_d0_252 = mux_d0_252;
    next_mux_d0_253 = mux_d0_253;
    next_mux_d0_254 = mux_d0_254;
    next_mux_d0_255 = mux_d0_255;
    next_mux_d1_0 = mux_d1_0;
    next_mux_d1_1 = mux_d1_1;
    next_mux_d1_2 = mux_d1_2;
    next_mux_d1_3 = mux_d1_3;
    next_mux_d1_4 = mux_d1_4;
    next_mux_d1_5 = mux_d1_5;
    next_mux_d1_6 = mux_d1_6;
    next_mux_d1_7 = mux_d1_7;
    next_mux_d1_8 = mux_d1_8;
    next_mux_d1_9 = mux_d1_9;
    next_mux_d1_10 = mux_d1_10;
    next_mux_d1_11 = mux_d1_11;
    next_mux_d1_12 = mux_d1_12;
    next_mux_d1_13 = mux_d1_13;
    next_mux_d1_14 = mux_d1_14;
    next_mux_d1_15 = mux_d1_15;
    next_mux_d1_16 = mux_d1_16;
    next_mux_d1_17 = mux_d1_17;
    next_mux_d1_18 = mux_d1_18;
    next_mux_d1_19 = mux_d1_19;
    next_mux_d1_20 = mux_d1_20;
    next_mux_d1_21 = mux_d1_21;
    next_mux_d1_22 = mux_d1_22;
    next_mux_d1_23 = mux_d1_23;
    next_mux_d1_24 = mux_d1_24;
    next_mux_d1_25 = mux_d1_25;
    next_mux_d1_26 = mux_d1_26;
    next_mux_d1_27 = mux_d1_27;
    next_mux_d1_28 = mux_d1_28;
    next_mux_d1_29 = mux_d1_29;
    next_mux_d1_30 = mux_d1_30;
    next_mux_d1_31 = mux_d1_31;
    next_mux_d2_0 = mux_d2_0;
    next_mux_d2_1 = mux_d2_1;
    next_mux_d2_2 = mux_d2_2;
    next_mux_d2_3 = mux_d2_3;
    next_mux_d3_0 = mux_d3_0;

    if (sel_d0_0[2:0] == 0) begin
        next_mux_d0_0 = input_word_d[0];
    end else if (sel_d0_0[2:0] == 1) begin
        next_mux_d0_0 = input_word_d[1];
    end else if (sel_d0_0[2:0] == 2) begin
        next_mux_d0_0 = input_word_d[2];
    end else if (sel_d0_0[2:0] == 3) begin
        next_mux_d0_0 = input_word_d[3];
    end else if (sel_d0_0[2:0] == 4) begin
        next_mux_d0_0 = input_word_d[4];
    end else if (sel_d0_0[2:0] == 5) begin
        next_mux_d0_0 = input_word_d[5];
    end else if (sel_d0_0[2:0] == 6) begin
        next_mux_d0_0 = input_word_d[6];
    end else begin
        next_mux_d0_0 = input_word_d[7];
    end

    if (sel_d0_1[2:0] == 0) begin
        next_mux_d0_1 = input_word_d[8];
    end else if (sel_d0_1[2:0] == 1) begin
        next_mux_d0_1 = input_word_d[9];
    end else if (sel_d0_1[2:0] == 2) begin
        next_mux_d0_1 = input_word_d[10];
    end else if (sel_d0_1[2:0] == 3) begin
        next_mux_d0_1 = input_word_d[11];
    end else if (sel_d0_1[2:0] == 4) begin
        next_mux_d0_1 = input_word_d[12];
    end else if (sel_d0_1[2:0] == 5) begin
        next_mux_d0_1 = input_word_d[13];
    end else if (sel_d0_1[2:0] == 6) begin
        next_mux_d0_1 = input_word_d[14];
    end else begin
        next_mux_d0_1 = input_word_d[15];
    end

    if (sel_d0_2[2:0] == 0) begin
        next_mux_d0_2 = input_word_d[16];
    end else if (sel_d0_2[2:0] == 1) begin
        next_mux_d0_2 = input_word_d[17];
    end else if (sel_d0_2[2:0] == 2) begin
        next_mux_d0_2 = input_word_d[18];
    end else if (sel_d0_2[2:0] == 3) begin
        next_mux_d0_2 = input_word_d[19];
    end else if (sel_d0_2[2:0] == 4) begin
        next_mux_d0_2 = input_word_d[20];
    end else if (sel_d0_2[2:0] == 5) begin
        next_mux_d0_2 = input_word_d[21];
    end else if (sel_d0_2[2:0] == 6) begin
        next_mux_d0_2 = input_word_d[22];
    end else begin
        next_mux_d0_2 = input_word_d[23];
    end

    if (sel_d0_3[2:0] == 0) begin
        next_mux_d0_3 = input_word_d[24];
    end else if (sel_d0_3[2:0] == 1) begin
        next_mux_d0_3 = input_word_d[25];
    end else if (sel_d0_3[2:0] == 2) begin
        next_mux_d0_3 = input_word_d[26];
    end else if (sel_d0_3[2:0] == 3) begin
        next_mux_d0_3 = input_word_d[27];
    end else if (sel_d0_3[2:0] == 4) begin
        next_mux_d0_3 = input_word_d[28];
    end else if (sel_d0_3[2:0] == 5) begin
        next_mux_d0_3 = input_word_d[29];
    end else if (sel_d0_3[2:0] == 6) begin
        next_mux_d0_3 = input_word_d[30];
    end else begin
        next_mux_d0_3 = input_word_d[31];
    end

    if (sel_d0_4[2:0] == 0) begin
        next_mux_d0_4 = input_word_d[32];
    end else if (sel_d0_4[2:0] == 1) begin
        next_mux_d0_4 = input_word_d[33];
    end else if (sel_d0_4[2:0] == 2) begin
        next_mux_d0_4 = input_word_d[34];
    end else if (sel_d0_4[2:0] == 3) begin
        next_mux_d0_4 = input_word_d[35];
    end else if (sel_d0_4[2:0] == 4) begin
        next_mux_d0_4 = input_word_d[36];
    end else if (sel_d0_4[2:0] == 5) begin
        next_mux_d0_4 = input_word_d[37];
    end else if (sel_d0_4[2:0] == 6) begin
        next_mux_d0_4 = input_word_d[38];
    end else begin
        next_mux_d0_4 = input_word_d[39];
    end

    if (sel_d0_5[2:0] == 0) begin
        next_mux_d0_5 = input_word_d[40];
    end else if (sel_d0_5[2:0] == 1) begin
        next_mux_d0_5 = input_word_d[41];
    end else if (sel_d0_5[2:0] == 2) begin
        next_mux_d0_5 = input_word_d[42];
    end else if (sel_d0_5[2:0] == 3) begin
        next_mux_d0_5 = input_word_d[43];
    end else if (sel_d0_5[2:0] == 4) begin
        next_mux_d0_5 = input_word_d[44];
    end else if (sel_d0_5[2:0] == 5) begin
        next_mux_d0_5 = input_word_d[45];
    end else if (sel_d0_5[2:0] == 6) begin
        next_mux_d0_5 = input_word_d[46];
    end else begin
        next_mux_d0_5 = input_word_d[47];
    end

    if (sel_d0_6[2:0] == 0) begin
        next_mux_d0_6 = input_word_d[48];
    end else if (sel_d0_6[2:0] == 1) begin
        next_mux_d0_6 = input_word_d[49];
    end else if (sel_d0_6[2:0] == 2) begin
        next_mux_d0_6 = input_word_d[50];
    end else if (sel_d0_6[2:0] == 3) begin
        next_mux_d0_6 = input_word_d[51];
    end else if (sel_d0_6[2:0] == 4) begin
        next_mux_d0_6 = input_word_d[52];
    end else if (sel_d0_6[2:0] == 5) begin
        next_mux_d0_6 = input_word_d[53];
    end else if (sel_d0_6[2:0] == 6) begin
        next_mux_d0_6 = input_word_d[54];
    end else begin
        next_mux_d0_6 = input_word_d[55];
    end

    if (sel_d0_7[2:0] == 0) begin
        next_mux_d0_7 = input_word_d[56];
    end else if (sel_d0_7[2:0] == 1) begin
        next_mux_d0_7 = input_word_d[57];
    end else if (sel_d0_7[2:0] == 2) begin
        next_mux_d0_7 = input_word_d[58];
    end else if (sel_d0_7[2:0] == 3) begin
        next_mux_d0_7 = input_word_d[59];
    end else if (sel_d0_7[2:0] == 4) begin
        next_mux_d0_7 = input_word_d[60];
    end else if (sel_d0_7[2:0] == 5) begin
        next_mux_d0_7 = input_word_d[61];
    end else if (sel_d0_7[2:0] == 6) begin
        next_mux_d0_7 = input_word_d[62];
    end else begin
        next_mux_d0_7 = input_word_d[63];
    end

    if (sel_d0_8[2:0] == 0) begin
        next_mux_d0_8 = input_word_d[64];
    end else if (sel_d0_8[2:0] == 1) begin
        next_mux_d0_8 = input_word_d[65];
    end else if (sel_d0_8[2:0] == 2) begin
        next_mux_d0_8 = input_word_d[66];
    end else if (sel_d0_8[2:0] == 3) begin
        next_mux_d0_8 = input_word_d[67];
    end else if (sel_d0_8[2:0] == 4) begin
        next_mux_d0_8 = input_word_d[68];
    end else if (sel_d0_8[2:0] == 5) begin
        next_mux_d0_8 = input_word_d[69];
    end else if (sel_d0_8[2:0] == 6) begin
        next_mux_d0_8 = input_word_d[70];
    end else begin
        next_mux_d0_8 = input_word_d[71];
    end

    if (sel_d0_9[2:0] == 0) begin
        next_mux_d0_9 = input_word_d[72];
    end else if (sel_d0_9[2:0] == 1) begin
        next_mux_d0_9 = input_word_d[73];
    end else if (sel_d0_9[2:0] == 2) begin
        next_mux_d0_9 = input_word_d[74];
    end else if (sel_d0_9[2:0] == 3) begin
        next_mux_d0_9 = input_word_d[75];
    end else if (sel_d0_9[2:0] == 4) begin
        next_mux_d0_9 = input_word_d[76];
    end else if (sel_d0_9[2:0] == 5) begin
        next_mux_d0_9 = input_word_d[77];
    end else if (sel_d0_9[2:0] == 6) begin
        next_mux_d0_9 = input_word_d[78];
    end else begin
        next_mux_d0_9 = input_word_d[79];
    end

    if (sel_d0_10[2:0] == 0) begin
        next_mux_d0_10 = input_word_d[80];
    end else if (sel_d0_10[2:0] == 1) begin
        next_mux_d0_10 = input_word_d[81];
    end else if (sel_d0_10[2:0] == 2) begin
        next_mux_d0_10 = input_word_d[82];
    end else if (sel_d0_10[2:0] == 3) begin
        next_mux_d0_10 = input_word_d[83];
    end else if (sel_d0_10[2:0] == 4) begin
        next_mux_d0_10 = input_word_d[84];
    end else if (sel_d0_10[2:0] == 5) begin
        next_mux_d0_10 = input_word_d[85];
    end else if (sel_d0_10[2:0] == 6) begin
        next_mux_d0_10 = input_word_d[86];
    end else begin
        next_mux_d0_10 = input_word_d[87];
    end

    if (sel_d0_11[2:0] == 0) begin
        next_mux_d0_11 = input_word_d[88];
    end else if (sel_d0_11[2:0] == 1) begin
        next_mux_d0_11 = input_word_d[89];
    end else if (sel_d0_11[2:0] == 2) begin
        next_mux_d0_11 = input_word_d[90];
    end else if (sel_d0_11[2:0] == 3) begin
        next_mux_d0_11 = input_word_d[91];
    end else if (sel_d0_11[2:0] == 4) begin
        next_mux_d0_11 = input_word_d[92];
    end else if (sel_d0_11[2:0] == 5) begin
        next_mux_d0_11 = input_word_d[93];
    end else if (sel_d0_11[2:0] == 6) begin
        next_mux_d0_11 = input_word_d[94];
    end else begin
        next_mux_d0_11 = input_word_d[95];
    end

    if (sel_d0_12[2:0] == 0) begin
        next_mux_d0_12 = input_word_d[96];
    end else if (sel_d0_12[2:0] == 1) begin
        next_mux_d0_12 = input_word_d[97];
    end else if (sel_d0_12[2:0] == 2) begin
        next_mux_d0_12 = input_word_d[98];
    end else if (sel_d0_12[2:0] == 3) begin
        next_mux_d0_12 = input_word_d[99];
    end else if (sel_d0_12[2:0] == 4) begin
        next_mux_d0_12 = input_word_d[100];
    end else if (sel_d0_12[2:0] == 5) begin
        next_mux_d0_12 = input_word_d[101];
    end else if (sel_d0_12[2:0] == 6) begin
        next_mux_d0_12 = input_word_d[102];
    end else begin
        next_mux_d0_12 = input_word_d[103];
    end

    if (sel_d0_13[2:0] == 0) begin
        next_mux_d0_13 = input_word_d[104];
    end else if (sel_d0_13[2:0] == 1) begin
        next_mux_d0_13 = input_word_d[105];
    end else if (sel_d0_13[2:0] == 2) begin
        next_mux_d0_13 = input_word_d[106];
    end else if (sel_d0_13[2:0] == 3) begin
        next_mux_d0_13 = input_word_d[107];
    end else if (sel_d0_13[2:0] == 4) begin
        next_mux_d0_13 = input_word_d[108];
    end else if (sel_d0_13[2:0] == 5) begin
        next_mux_d0_13 = input_word_d[109];
    end else if (sel_d0_13[2:0] == 6) begin
        next_mux_d0_13 = input_word_d[110];
    end else begin
        next_mux_d0_13 = input_word_d[111];
    end

    if (sel_d0_14[2:0] == 0) begin
        next_mux_d0_14 = input_word_d[112];
    end else if (sel_d0_14[2:0] == 1) begin
        next_mux_d0_14 = input_word_d[113];
    end else if (sel_d0_14[2:0] == 2) begin
        next_mux_d0_14 = input_word_d[114];
    end else if (sel_d0_14[2:0] == 3) begin
        next_mux_d0_14 = input_word_d[115];
    end else if (sel_d0_14[2:0] == 4) begin
        next_mux_d0_14 = input_word_d[116];
    end else if (sel_d0_14[2:0] == 5) begin
        next_mux_d0_14 = input_word_d[117];
    end else if (sel_d0_14[2:0] == 6) begin
        next_mux_d0_14 = input_word_d[118];
    end else begin
        next_mux_d0_14 = input_word_d[119];
    end

    if (sel_d0_15[2:0] == 0) begin
        next_mux_d0_15 = input_word_d[120];
    end else if (sel_d0_15[2:0] == 1) begin
        next_mux_d0_15 = input_word_d[121];
    end else if (sel_d0_15[2:0] == 2) begin
        next_mux_d0_15 = input_word_d[122];
    end else if (sel_d0_15[2:0] == 3) begin
        next_mux_d0_15 = input_word_d[123];
    end else if (sel_d0_15[2:0] == 4) begin
        next_mux_d0_15 = input_word_d[124];
    end else if (sel_d0_15[2:0] == 5) begin
        next_mux_d0_15 = input_word_d[125];
    end else if (sel_d0_15[2:0] == 6) begin
        next_mux_d0_15 = input_word_d[126];
    end else begin
        next_mux_d0_15 = input_word_d[127];
    end

    if (sel_d0_16[2:0] == 0) begin
        next_mux_d0_16 = input_word_d[128];
    end else if (sel_d0_16[2:0] == 1) begin
        next_mux_d0_16 = input_word_d[129];
    end else if (sel_d0_16[2:0] == 2) begin
        next_mux_d0_16 = input_word_d[130];
    end else if (sel_d0_16[2:0] == 3) begin
        next_mux_d0_16 = input_word_d[131];
    end else if (sel_d0_16[2:0] == 4) begin
        next_mux_d0_16 = input_word_d[132];
    end else if (sel_d0_16[2:0] == 5) begin
        next_mux_d0_16 = input_word_d[133];
    end else if (sel_d0_16[2:0] == 6) begin
        next_mux_d0_16 = input_word_d[134];
    end else begin
        next_mux_d0_16 = input_word_d[135];
    end

    if (sel_d0_17[2:0] == 0) begin
        next_mux_d0_17 = input_word_d[136];
    end else if (sel_d0_17[2:0] == 1) begin
        next_mux_d0_17 = input_word_d[137];
    end else if (sel_d0_17[2:0] == 2) begin
        next_mux_d0_17 = input_word_d[138];
    end else if (sel_d0_17[2:0] == 3) begin
        next_mux_d0_17 = input_word_d[139];
    end else if (sel_d0_17[2:0] == 4) begin
        next_mux_d0_17 = input_word_d[140];
    end else if (sel_d0_17[2:0] == 5) begin
        next_mux_d0_17 = input_word_d[141];
    end else if (sel_d0_17[2:0] == 6) begin
        next_mux_d0_17 = input_word_d[142];
    end else begin
        next_mux_d0_17 = input_word_d[143];
    end

    if (sel_d0_18[2:0] == 0) begin
        next_mux_d0_18 = input_word_d[144];
    end else if (sel_d0_18[2:0] == 1) begin
        next_mux_d0_18 = input_word_d[145];
    end else if (sel_d0_18[2:0] == 2) begin
        next_mux_d0_18 = input_word_d[146];
    end else if (sel_d0_18[2:0] == 3) begin
        next_mux_d0_18 = input_word_d[147];
    end else if (sel_d0_18[2:0] == 4) begin
        next_mux_d0_18 = input_word_d[148];
    end else if (sel_d0_18[2:0] == 5) begin
        next_mux_d0_18 = input_word_d[149];
    end else if (sel_d0_18[2:0] == 6) begin
        next_mux_d0_18 = input_word_d[150];
    end else begin
        next_mux_d0_18 = input_word_d[151];
    end

    if (sel_d0_19[2:0] == 0) begin
        next_mux_d0_19 = input_word_d[152];
    end else if (sel_d0_19[2:0] == 1) begin
        next_mux_d0_19 = input_word_d[153];
    end else if (sel_d0_19[2:0] == 2) begin
        next_mux_d0_19 = input_word_d[154];
    end else if (sel_d0_19[2:0] == 3) begin
        next_mux_d0_19 = input_word_d[155];
    end else if (sel_d0_19[2:0] == 4) begin
        next_mux_d0_19 = input_word_d[156];
    end else if (sel_d0_19[2:0] == 5) begin
        next_mux_d0_19 = input_word_d[157];
    end else if (sel_d0_19[2:0] == 6) begin
        next_mux_d0_19 = input_word_d[158];
    end else begin
        next_mux_d0_19 = input_word_d[159];
    end

    if (sel_d0_20[2:0] == 0) begin
        next_mux_d0_20 = input_word_d[160];
    end else if (sel_d0_20[2:0] == 1) begin
        next_mux_d0_20 = input_word_d[161];
    end else if (sel_d0_20[2:0] == 2) begin
        next_mux_d0_20 = input_word_d[162];
    end else if (sel_d0_20[2:0] == 3) begin
        next_mux_d0_20 = input_word_d[163];
    end else if (sel_d0_20[2:0] == 4) begin
        next_mux_d0_20 = input_word_d[164];
    end else if (sel_d0_20[2:0] == 5) begin
        next_mux_d0_20 = input_word_d[165];
    end else if (sel_d0_20[2:0] == 6) begin
        next_mux_d0_20 = input_word_d[166];
    end else begin
        next_mux_d0_20 = input_word_d[167];
    end

    if (sel_d0_21[2:0] == 0) begin
        next_mux_d0_21 = input_word_d[168];
    end else if (sel_d0_21[2:0] == 1) begin
        next_mux_d0_21 = input_word_d[169];
    end else if (sel_d0_21[2:0] == 2) begin
        next_mux_d0_21 = input_word_d[170];
    end else if (sel_d0_21[2:0] == 3) begin
        next_mux_d0_21 = input_word_d[171];
    end else if (sel_d0_21[2:0] == 4) begin
        next_mux_d0_21 = input_word_d[172];
    end else if (sel_d0_21[2:0] == 5) begin
        next_mux_d0_21 = input_word_d[173];
    end else if (sel_d0_21[2:0] == 6) begin
        next_mux_d0_21 = input_word_d[174];
    end else begin
        next_mux_d0_21 = input_word_d[175];
    end

    if (sel_d0_22[2:0] == 0) begin
        next_mux_d0_22 = input_word_d[176];
    end else if (sel_d0_22[2:0] == 1) begin
        next_mux_d0_22 = input_word_d[177];
    end else if (sel_d0_22[2:0] == 2) begin
        next_mux_d0_22 = input_word_d[178];
    end else if (sel_d0_22[2:0] == 3) begin
        next_mux_d0_22 = input_word_d[179];
    end else if (sel_d0_22[2:0] == 4) begin
        next_mux_d0_22 = input_word_d[180];
    end else if (sel_d0_22[2:0] == 5) begin
        next_mux_d0_22 = input_word_d[181];
    end else if (sel_d0_22[2:0] == 6) begin
        next_mux_d0_22 = input_word_d[182];
    end else begin
        next_mux_d0_22 = input_word_d[183];
    end

    if (sel_d0_23[2:0] == 0) begin
        next_mux_d0_23 = input_word_d[184];
    end else if (sel_d0_23[2:0] == 1) begin
        next_mux_d0_23 = input_word_d[185];
    end else if (sel_d0_23[2:0] == 2) begin
        next_mux_d0_23 = input_word_d[186];
    end else if (sel_d0_23[2:0] == 3) begin
        next_mux_d0_23 = input_word_d[187];
    end else if (sel_d0_23[2:0] == 4) begin
        next_mux_d0_23 = input_word_d[188];
    end else if (sel_d0_23[2:0] == 5) begin
        next_mux_d0_23 = input_word_d[189];
    end else if (sel_d0_23[2:0] == 6) begin
        next_mux_d0_23 = input_word_d[190];
    end else begin
        next_mux_d0_23 = input_word_d[191];
    end

    if (sel_d0_24[2:0] == 0) begin
        next_mux_d0_24 = input_word_d[192];
    end else if (sel_d0_24[2:0] == 1) begin
        next_mux_d0_24 = input_word_d[193];
    end else if (sel_d0_24[2:0] == 2) begin
        next_mux_d0_24 = input_word_d[194];
    end else if (sel_d0_24[2:0] == 3) begin
        next_mux_d0_24 = input_word_d[195];
    end else if (sel_d0_24[2:0] == 4) begin
        next_mux_d0_24 = input_word_d[196];
    end else if (sel_d0_24[2:0] == 5) begin
        next_mux_d0_24 = input_word_d[197];
    end else if (sel_d0_24[2:0] == 6) begin
        next_mux_d0_24 = input_word_d[198];
    end else begin
        next_mux_d0_24 = input_word_d[199];
    end

    if (sel_d0_25[2:0] == 0) begin
        next_mux_d0_25 = input_word_d[200];
    end else if (sel_d0_25[2:0] == 1) begin
        next_mux_d0_25 = input_word_d[201];
    end else if (sel_d0_25[2:0] == 2) begin
        next_mux_d0_25 = input_word_d[202];
    end else if (sel_d0_25[2:0] == 3) begin
        next_mux_d0_25 = input_word_d[203];
    end else if (sel_d0_25[2:0] == 4) begin
        next_mux_d0_25 = input_word_d[204];
    end else if (sel_d0_25[2:0] == 5) begin
        next_mux_d0_25 = input_word_d[205];
    end else if (sel_d0_25[2:0] == 6) begin
        next_mux_d0_25 = input_word_d[206];
    end else begin
        next_mux_d0_25 = input_word_d[207];
    end

    if (sel_d0_26[2:0] == 0) begin
        next_mux_d0_26 = input_word_d[208];
    end else if (sel_d0_26[2:0] == 1) begin
        next_mux_d0_26 = input_word_d[209];
    end else if (sel_d0_26[2:0] == 2) begin
        next_mux_d0_26 = input_word_d[210];
    end else if (sel_d0_26[2:0] == 3) begin
        next_mux_d0_26 = input_word_d[211];
    end else if (sel_d0_26[2:0] == 4) begin
        next_mux_d0_26 = input_word_d[212];
    end else if (sel_d0_26[2:0] == 5) begin
        next_mux_d0_26 = input_word_d[213];
    end else if (sel_d0_26[2:0] == 6) begin
        next_mux_d0_26 = input_word_d[214];
    end else begin
        next_mux_d0_26 = input_word_d[215];
    end

    if (sel_d0_27[2:0] == 0) begin
        next_mux_d0_27 = input_word_d[216];
    end else if (sel_d0_27[2:0] == 1) begin
        next_mux_d0_27 = input_word_d[217];
    end else if (sel_d0_27[2:0] == 2) begin
        next_mux_d0_27 = input_word_d[218];
    end else if (sel_d0_27[2:0] == 3) begin
        next_mux_d0_27 = input_word_d[219];
    end else if (sel_d0_27[2:0] == 4) begin
        next_mux_d0_27 = input_word_d[220];
    end else if (sel_d0_27[2:0] == 5) begin
        next_mux_d0_27 = input_word_d[221];
    end else if (sel_d0_27[2:0] == 6) begin
        next_mux_d0_27 = input_word_d[222];
    end else begin
        next_mux_d0_27 = input_word_d[223];
    end

    if (sel_d0_28[2:0] == 0) begin
        next_mux_d0_28 = input_word_d[224];
    end else if (sel_d0_28[2:0] == 1) begin
        next_mux_d0_28 = input_word_d[225];
    end else if (sel_d0_28[2:0] == 2) begin
        next_mux_d0_28 = input_word_d[226];
    end else if (sel_d0_28[2:0] == 3) begin
        next_mux_d0_28 = input_word_d[227];
    end else if (sel_d0_28[2:0] == 4) begin
        next_mux_d0_28 = input_word_d[228];
    end else if (sel_d0_28[2:0] == 5) begin
        next_mux_d0_28 = input_word_d[229];
    end else if (sel_d0_28[2:0] == 6) begin
        next_mux_d0_28 = input_word_d[230];
    end else begin
        next_mux_d0_28 = input_word_d[231];
    end

    if (sel_d0_29[2:0] == 0) begin
        next_mux_d0_29 = input_word_d[232];
    end else if (sel_d0_29[2:0] == 1) begin
        next_mux_d0_29 = input_word_d[233];
    end else if (sel_d0_29[2:0] == 2) begin
        next_mux_d0_29 = input_word_d[234];
    end else if (sel_d0_29[2:0] == 3) begin
        next_mux_d0_29 = input_word_d[235];
    end else if (sel_d0_29[2:0] == 4) begin
        next_mux_d0_29 = input_word_d[236];
    end else if (sel_d0_29[2:0] == 5) begin
        next_mux_d0_29 = input_word_d[237];
    end else if (sel_d0_29[2:0] == 6) begin
        next_mux_d0_29 = input_word_d[238];
    end else begin
        next_mux_d0_29 = input_word_d[239];
    end

    if (sel_d0_30[2:0] == 0) begin
        next_mux_d0_30 = input_word_d[240];
    end else if (sel_d0_30[2:0] == 1) begin
        next_mux_d0_30 = input_word_d[241];
    end else if (sel_d0_30[2:0] == 2) begin
        next_mux_d0_30 = input_word_d[242];
    end else if (sel_d0_30[2:0] == 3) begin
        next_mux_d0_30 = input_word_d[243];
    end else if (sel_d0_30[2:0] == 4) begin
        next_mux_d0_30 = input_word_d[244];
    end else if (sel_d0_30[2:0] == 5) begin
        next_mux_d0_30 = input_word_d[245];
    end else if (sel_d0_30[2:0] == 6) begin
        next_mux_d0_30 = input_word_d[246];
    end else begin
        next_mux_d0_30 = input_word_d[247];
    end

    if (sel_d0_31[2:0] == 0) begin
        next_mux_d0_31 = input_word_d[248];
    end else if (sel_d0_31[2:0] == 1) begin
        next_mux_d0_31 = input_word_d[249];
    end else if (sel_d0_31[2:0] == 2) begin
        next_mux_d0_31 = input_word_d[250];
    end else if (sel_d0_31[2:0] == 3) begin
        next_mux_d0_31 = input_word_d[251];
    end else if (sel_d0_31[2:0] == 4) begin
        next_mux_d0_31 = input_word_d[252];
    end else if (sel_d0_31[2:0] == 5) begin
        next_mux_d0_31 = input_word_d[253];
    end else if (sel_d0_31[2:0] == 6) begin
        next_mux_d0_31 = input_word_d[254];
    end else begin
        next_mux_d0_31 = input_word_d[255];
    end

    if (sel_d0_32[2:0] == 0) begin
        next_mux_d0_32 = input_word_d[256];
    end else if (sel_d0_32[2:0] == 1) begin
        next_mux_d0_32 = input_word_d[257];
    end else if (sel_d0_32[2:0] == 2) begin
        next_mux_d0_32 = input_word_d[258];
    end else if (sel_d0_32[2:0] == 3) begin
        next_mux_d0_32 = input_word_d[259];
    end else if (sel_d0_32[2:0] == 4) begin
        next_mux_d0_32 = input_word_d[260];
    end else if (sel_d0_32[2:0] == 5) begin
        next_mux_d0_32 = input_word_d[261];
    end else if (sel_d0_32[2:0] == 6) begin
        next_mux_d0_32 = input_word_d[262];
    end else begin
        next_mux_d0_32 = input_word_d[263];
    end

    if (sel_d0_33[2:0] == 0) begin
        next_mux_d0_33 = input_word_d[264];
    end else if (sel_d0_33[2:0] == 1) begin
        next_mux_d0_33 = input_word_d[265];
    end else if (sel_d0_33[2:0] == 2) begin
        next_mux_d0_33 = input_word_d[266];
    end else if (sel_d0_33[2:0] == 3) begin
        next_mux_d0_33 = input_word_d[267];
    end else if (sel_d0_33[2:0] == 4) begin
        next_mux_d0_33 = input_word_d[268];
    end else if (sel_d0_33[2:0] == 5) begin
        next_mux_d0_33 = input_word_d[269];
    end else if (sel_d0_33[2:0] == 6) begin
        next_mux_d0_33 = input_word_d[270];
    end else begin
        next_mux_d0_33 = input_word_d[271];
    end

    if (sel_d0_34[2:0] == 0) begin
        next_mux_d0_34 = input_word_d[272];
    end else if (sel_d0_34[2:0] == 1) begin
        next_mux_d0_34 = input_word_d[273];
    end else if (sel_d0_34[2:0] == 2) begin
        next_mux_d0_34 = input_word_d[274];
    end else if (sel_d0_34[2:0] == 3) begin
        next_mux_d0_34 = input_word_d[275];
    end else if (sel_d0_34[2:0] == 4) begin
        next_mux_d0_34 = input_word_d[276];
    end else if (sel_d0_34[2:0] == 5) begin
        next_mux_d0_34 = input_word_d[277];
    end else if (sel_d0_34[2:0] == 6) begin
        next_mux_d0_34 = input_word_d[278];
    end else begin
        next_mux_d0_34 = input_word_d[279];
    end

    if (sel_d0_35[2:0] == 0) begin
        next_mux_d0_35 = input_word_d[280];
    end else if (sel_d0_35[2:0] == 1) begin
        next_mux_d0_35 = input_word_d[281];
    end else if (sel_d0_35[2:0] == 2) begin
        next_mux_d0_35 = input_word_d[282];
    end else if (sel_d0_35[2:0] == 3) begin
        next_mux_d0_35 = input_word_d[283];
    end else if (sel_d0_35[2:0] == 4) begin
        next_mux_d0_35 = input_word_d[284];
    end else if (sel_d0_35[2:0] == 5) begin
        next_mux_d0_35 = input_word_d[285];
    end else if (sel_d0_35[2:0] == 6) begin
        next_mux_d0_35 = input_word_d[286];
    end else begin
        next_mux_d0_35 = input_word_d[287];
    end

    if (sel_d0_36[2:0] == 0) begin
        next_mux_d0_36 = input_word_d[288];
    end else if (sel_d0_36[2:0] == 1) begin
        next_mux_d0_36 = input_word_d[289];
    end else if (sel_d0_36[2:0] == 2) begin
        next_mux_d0_36 = input_word_d[290];
    end else if (sel_d0_36[2:0] == 3) begin
        next_mux_d0_36 = input_word_d[291];
    end else if (sel_d0_36[2:0] == 4) begin
        next_mux_d0_36 = input_word_d[292];
    end else if (sel_d0_36[2:0] == 5) begin
        next_mux_d0_36 = input_word_d[293];
    end else if (sel_d0_36[2:0] == 6) begin
        next_mux_d0_36 = input_word_d[294];
    end else begin
        next_mux_d0_36 = input_word_d[295];
    end

    if (sel_d0_37[2:0] == 0) begin
        next_mux_d0_37 = input_word_d[296];
    end else if (sel_d0_37[2:0] == 1) begin
        next_mux_d0_37 = input_word_d[297];
    end else if (sel_d0_37[2:0] == 2) begin
        next_mux_d0_37 = input_word_d[298];
    end else if (sel_d0_37[2:0] == 3) begin
        next_mux_d0_37 = input_word_d[299];
    end else if (sel_d0_37[2:0] == 4) begin
        next_mux_d0_37 = input_word_d[300];
    end else if (sel_d0_37[2:0] == 5) begin
        next_mux_d0_37 = input_word_d[301];
    end else if (sel_d0_37[2:0] == 6) begin
        next_mux_d0_37 = input_word_d[302];
    end else begin
        next_mux_d0_37 = input_word_d[303];
    end

    if (sel_d0_38[2:0] == 0) begin
        next_mux_d0_38 = input_word_d[304];
    end else if (sel_d0_38[2:0] == 1) begin
        next_mux_d0_38 = input_word_d[305];
    end else if (sel_d0_38[2:0] == 2) begin
        next_mux_d0_38 = input_word_d[306];
    end else if (sel_d0_38[2:0] == 3) begin
        next_mux_d0_38 = input_word_d[307];
    end else if (sel_d0_38[2:0] == 4) begin
        next_mux_d0_38 = input_word_d[308];
    end else if (sel_d0_38[2:0] == 5) begin
        next_mux_d0_38 = input_word_d[309];
    end else if (sel_d0_38[2:0] == 6) begin
        next_mux_d0_38 = input_word_d[310];
    end else begin
        next_mux_d0_38 = input_word_d[311];
    end

    if (sel_d0_39[2:0] == 0) begin
        next_mux_d0_39 = input_word_d[312];
    end else if (sel_d0_39[2:0] == 1) begin
        next_mux_d0_39 = input_word_d[313];
    end else if (sel_d0_39[2:0] == 2) begin
        next_mux_d0_39 = input_word_d[314];
    end else if (sel_d0_39[2:0] == 3) begin
        next_mux_d0_39 = input_word_d[315];
    end else if (sel_d0_39[2:0] == 4) begin
        next_mux_d0_39 = input_word_d[316];
    end else if (sel_d0_39[2:0] == 5) begin
        next_mux_d0_39 = input_word_d[317];
    end else if (sel_d0_39[2:0] == 6) begin
        next_mux_d0_39 = input_word_d[318];
    end else begin
        next_mux_d0_39 = input_word_d[319];
    end

    if (sel_d0_40[2:0] == 0) begin
        next_mux_d0_40 = input_word_d[320];
    end else if (sel_d0_40[2:0] == 1) begin
        next_mux_d0_40 = input_word_d[321];
    end else if (sel_d0_40[2:0] == 2) begin
        next_mux_d0_40 = input_word_d[322];
    end else if (sel_d0_40[2:0] == 3) begin
        next_mux_d0_40 = input_word_d[323];
    end else if (sel_d0_40[2:0] == 4) begin
        next_mux_d0_40 = input_word_d[324];
    end else if (sel_d0_40[2:0] == 5) begin
        next_mux_d0_40 = input_word_d[325];
    end else if (sel_d0_40[2:0] == 6) begin
        next_mux_d0_40 = input_word_d[326];
    end else begin
        next_mux_d0_40 = input_word_d[327];
    end

    if (sel_d0_41[2:0] == 0) begin
        next_mux_d0_41 = input_word_d[328];
    end else if (sel_d0_41[2:0] == 1) begin
        next_mux_d0_41 = input_word_d[329];
    end else if (sel_d0_41[2:0] == 2) begin
        next_mux_d0_41 = input_word_d[330];
    end else if (sel_d0_41[2:0] == 3) begin
        next_mux_d0_41 = input_word_d[331];
    end else if (sel_d0_41[2:0] == 4) begin
        next_mux_d0_41 = input_word_d[332];
    end else if (sel_d0_41[2:0] == 5) begin
        next_mux_d0_41 = input_word_d[333];
    end else if (sel_d0_41[2:0] == 6) begin
        next_mux_d0_41 = input_word_d[334];
    end else begin
        next_mux_d0_41 = input_word_d[335];
    end

    if (sel_d0_42[2:0] == 0) begin
        next_mux_d0_42 = input_word_d[336];
    end else if (sel_d0_42[2:0] == 1) begin
        next_mux_d0_42 = input_word_d[337];
    end else if (sel_d0_42[2:0] == 2) begin
        next_mux_d0_42 = input_word_d[338];
    end else if (sel_d0_42[2:0] == 3) begin
        next_mux_d0_42 = input_word_d[339];
    end else if (sel_d0_42[2:0] == 4) begin
        next_mux_d0_42 = input_word_d[340];
    end else if (sel_d0_42[2:0] == 5) begin
        next_mux_d0_42 = input_word_d[341];
    end else if (sel_d0_42[2:0] == 6) begin
        next_mux_d0_42 = input_word_d[342];
    end else begin
        next_mux_d0_42 = input_word_d[343];
    end

    if (sel_d0_43[2:0] == 0) begin
        next_mux_d0_43 = input_word_d[344];
    end else if (sel_d0_43[2:0] == 1) begin
        next_mux_d0_43 = input_word_d[345];
    end else if (sel_d0_43[2:0] == 2) begin
        next_mux_d0_43 = input_word_d[346];
    end else if (sel_d0_43[2:0] == 3) begin
        next_mux_d0_43 = input_word_d[347];
    end else if (sel_d0_43[2:0] == 4) begin
        next_mux_d0_43 = input_word_d[348];
    end else if (sel_d0_43[2:0] == 5) begin
        next_mux_d0_43 = input_word_d[349];
    end else if (sel_d0_43[2:0] == 6) begin
        next_mux_d0_43 = input_word_d[350];
    end else begin
        next_mux_d0_43 = input_word_d[351];
    end

    if (sel_d0_44[2:0] == 0) begin
        next_mux_d0_44 = input_word_d[352];
    end else if (sel_d0_44[2:0] == 1) begin
        next_mux_d0_44 = input_word_d[353];
    end else if (sel_d0_44[2:0] == 2) begin
        next_mux_d0_44 = input_word_d[354];
    end else if (sel_d0_44[2:0] == 3) begin
        next_mux_d0_44 = input_word_d[355];
    end else if (sel_d0_44[2:0] == 4) begin
        next_mux_d0_44 = input_word_d[356];
    end else if (sel_d0_44[2:0] == 5) begin
        next_mux_d0_44 = input_word_d[357];
    end else if (sel_d0_44[2:0] == 6) begin
        next_mux_d0_44 = input_word_d[358];
    end else begin
        next_mux_d0_44 = input_word_d[359];
    end

    if (sel_d0_45[2:0] == 0) begin
        next_mux_d0_45 = input_word_d[360];
    end else if (sel_d0_45[2:0] == 1) begin
        next_mux_d0_45 = input_word_d[361];
    end else if (sel_d0_45[2:0] == 2) begin
        next_mux_d0_45 = input_word_d[362];
    end else if (sel_d0_45[2:0] == 3) begin
        next_mux_d0_45 = input_word_d[363];
    end else if (sel_d0_45[2:0] == 4) begin
        next_mux_d0_45 = input_word_d[364];
    end else if (sel_d0_45[2:0] == 5) begin
        next_mux_d0_45 = input_word_d[365];
    end else if (sel_d0_45[2:0] == 6) begin
        next_mux_d0_45 = input_word_d[366];
    end else begin
        next_mux_d0_45 = input_word_d[367];
    end

    if (sel_d0_46[2:0] == 0) begin
        next_mux_d0_46 = input_word_d[368];
    end else if (sel_d0_46[2:0] == 1) begin
        next_mux_d0_46 = input_word_d[369];
    end else if (sel_d0_46[2:0] == 2) begin
        next_mux_d0_46 = input_word_d[370];
    end else if (sel_d0_46[2:0] == 3) begin
        next_mux_d0_46 = input_word_d[371];
    end else if (sel_d0_46[2:0] == 4) begin
        next_mux_d0_46 = input_word_d[372];
    end else if (sel_d0_46[2:0] == 5) begin
        next_mux_d0_46 = input_word_d[373];
    end else if (sel_d0_46[2:0] == 6) begin
        next_mux_d0_46 = input_word_d[374];
    end else begin
        next_mux_d0_46 = input_word_d[375];
    end

    if (sel_d0_47[2:0] == 0) begin
        next_mux_d0_47 = input_word_d[376];
    end else if (sel_d0_47[2:0] == 1) begin
        next_mux_d0_47 = input_word_d[377];
    end else if (sel_d0_47[2:0] == 2) begin
        next_mux_d0_47 = input_word_d[378];
    end else if (sel_d0_47[2:0] == 3) begin
        next_mux_d0_47 = input_word_d[379];
    end else if (sel_d0_47[2:0] == 4) begin
        next_mux_d0_47 = input_word_d[380];
    end else if (sel_d0_47[2:0] == 5) begin
        next_mux_d0_47 = input_word_d[381];
    end else if (sel_d0_47[2:0] == 6) begin
        next_mux_d0_47 = input_word_d[382];
    end else begin
        next_mux_d0_47 = input_word_d[383];
    end

    if (sel_d0_48[2:0] == 0) begin
        next_mux_d0_48 = input_word_d[384];
    end else if (sel_d0_48[2:0] == 1) begin
        next_mux_d0_48 = input_word_d[385];
    end else if (sel_d0_48[2:0] == 2) begin
        next_mux_d0_48 = input_word_d[386];
    end else if (sel_d0_48[2:0] == 3) begin
        next_mux_d0_48 = input_word_d[387];
    end else if (sel_d0_48[2:0] == 4) begin
        next_mux_d0_48 = input_word_d[388];
    end else if (sel_d0_48[2:0] == 5) begin
        next_mux_d0_48 = input_word_d[389];
    end else if (sel_d0_48[2:0] == 6) begin
        next_mux_d0_48 = input_word_d[390];
    end else begin
        next_mux_d0_48 = input_word_d[391];
    end

    if (sel_d0_49[2:0] == 0) begin
        next_mux_d0_49 = input_word_d[392];
    end else if (sel_d0_49[2:0] == 1) begin
        next_mux_d0_49 = input_word_d[393];
    end else if (sel_d0_49[2:0] == 2) begin
        next_mux_d0_49 = input_word_d[394];
    end else if (sel_d0_49[2:0] == 3) begin
        next_mux_d0_49 = input_word_d[395];
    end else if (sel_d0_49[2:0] == 4) begin
        next_mux_d0_49 = input_word_d[396];
    end else if (sel_d0_49[2:0] == 5) begin
        next_mux_d0_49 = input_word_d[397];
    end else if (sel_d0_49[2:0] == 6) begin
        next_mux_d0_49 = input_word_d[398];
    end else begin
        next_mux_d0_49 = input_word_d[399];
    end

    if (sel_d0_50[2:0] == 0) begin
        next_mux_d0_50 = input_word_d[400];
    end else if (sel_d0_50[2:0] == 1) begin
        next_mux_d0_50 = input_word_d[401];
    end else if (sel_d0_50[2:0] == 2) begin
        next_mux_d0_50 = input_word_d[402];
    end else if (sel_d0_50[2:0] == 3) begin
        next_mux_d0_50 = input_word_d[403];
    end else if (sel_d0_50[2:0] == 4) begin
        next_mux_d0_50 = input_word_d[404];
    end else if (sel_d0_50[2:0] == 5) begin
        next_mux_d0_50 = input_word_d[405];
    end else if (sel_d0_50[2:0] == 6) begin
        next_mux_d0_50 = input_word_d[406];
    end else begin
        next_mux_d0_50 = input_word_d[407];
    end

    if (sel_d0_51[2:0] == 0) begin
        next_mux_d0_51 = input_word_d[408];
    end else if (sel_d0_51[2:0] == 1) begin
        next_mux_d0_51 = input_word_d[409];
    end else if (sel_d0_51[2:0] == 2) begin
        next_mux_d0_51 = input_word_d[410];
    end else if (sel_d0_51[2:0] == 3) begin
        next_mux_d0_51 = input_word_d[411];
    end else if (sel_d0_51[2:0] == 4) begin
        next_mux_d0_51 = input_word_d[412];
    end else if (sel_d0_51[2:0] == 5) begin
        next_mux_d0_51 = input_word_d[413];
    end else if (sel_d0_51[2:0] == 6) begin
        next_mux_d0_51 = input_word_d[414];
    end else begin
        next_mux_d0_51 = input_word_d[415];
    end

    if (sel_d0_52[2:0] == 0) begin
        next_mux_d0_52 = input_word_d[416];
    end else if (sel_d0_52[2:0] == 1) begin
        next_mux_d0_52 = input_word_d[417];
    end else if (sel_d0_52[2:0] == 2) begin
        next_mux_d0_52 = input_word_d[418];
    end else if (sel_d0_52[2:0] == 3) begin
        next_mux_d0_52 = input_word_d[419];
    end else if (sel_d0_52[2:0] == 4) begin
        next_mux_d0_52 = input_word_d[420];
    end else if (sel_d0_52[2:0] == 5) begin
        next_mux_d0_52 = input_word_d[421];
    end else if (sel_d0_52[2:0] == 6) begin
        next_mux_d0_52 = input_word_d[422];
    end else begin
        next_mux_d0_52 = input_word_d[423];
    end

    if (sel_d0_53[2:0] == 0) begin
        next_mux_d0_53 = input_word_d[424];
    end else if (sel_d0_53[2:0] == 1) begin
        next_mux_d0_53 = input_word_d[425];
    end else if (sel_d0_53[2:0] == 2) begin
        next_mux_d0_53 = input_word_d[426];
    end else if (sel_d0_53[2:0] == 3) begin
        next_mux_d0_53 = input_word_d[427];
    end else if (sel_d0_53[2:0] == 4) begin
        next_mux_d0_53 = input_word_d[428];
    end else if (sel_d0_53[2:0] == 5) begin
        next_mux_d0_53 = input_word_d[429];
    end else if (sel_d0_53[2:0] == 6) begin
        next_mux_d0_53 = input_word_d[430];
    end else begin
        next_mux_d0_53 = input_word_d[431];
    end

    if (sel_d0_54[2:0] == 0) begin
        next_mux_d0_54 = input_word_d[432];
    end else if (sel_d0_54[2:0] == 1) begin
        next_mux_d0_54 = input_word_d[433];
    end else if (sel_d0_54[2:0] == 2) begin
        next_mux_d0_54 = input_word_d[434];
    end else if (sel_d0_54[2:0] == 3) begin
        next_mux_d0_54 = input_word_d[435];
    end else if (sel_d0_54[2:0] == 4) begin
        next_mux_d0_54 = input_word_d[436];
    end else if (sel_d0_54[2:0] == 5) begin
        next_mux_d0_54 = input_word_d[437];
    end else if (sel_d0_54[2:0] == 6) begin
        next_mux_d0_54 = input_word_d[438];
    end else begin
        next_mux_d0_54 = input_word_d[439];
    end

    if (sel_d0_55[2:0] == 0) begin
        next_mux_d0_55 = input_word_d[440];
    end else if (sel_d0_55[2:0] == 1) begin
        next_mux_d0_55 = input_word_d[441];
    end else if (sel_d0_55[2:0] == 2) begin
        next_mux_d0_55 = input_word_d[442];
    end else if (sel_d0_55[2:0] == 3) begin
        next_mux_d0_55 = input_word_d[443];
    end else if (sel_d0_55[2:0] == 4) begin
        next_mux_d0_55 = input_word_d[444];
    end else if (sel_d0_55[2:0] == 5) begin
        next_mux_d0_55 = input_word_d[445];
    end else if (sel_d0_55[2:0] == 6) begin
        next_mux_d0_55 = input_word_d[446];
    end else begin
        next_mux_d0_55 = input_word_d[447];
    end

    if (sel_d0_56[2:0] == 0) begin
        next_mux_d0_56 = input_word_d[448];
    end else if (sel_d0_56[2:0] == 1) begin
        next_mux_d0_56 = input_word_d[449];
    end else if (sel_d0_56[2:0] == 2) begin
        next_mux_d0_56 = input_word_d[450];
    end else if (sel_d0_56[2:0] == 3) begin
        next_mux_d0_56 = input_word_d[451];
    end else if (sel_d0_56[2:0] == 4) begin
        next_mux_d0_56 = input_word_d[452];
    end else if (sel_d0_56[2:0] == 5) begin
        next_mux_d0_56 = input_word_d[453];
    end else if (sel_d0_56[2:0] == 6) begin
        next_mux_d0_56 = input_word_d[454];
    end else begin
        next_mux_d0_56 = input_word_d[455];
    end

    if (sel_d0_57[2:0] == 0) begin
        next_mux_d0_57 = input_word_d[456];
    end else if (sel_d0_57[2:0] == 1) begin
        next_mux_d0_57 = input_word_d[457];
    end else if (sel_d0_57[2:0] == 2) begin
        next_mux_d0_57 = input_word_d[458];
    end else if (sel_d0_57[2:0] == 3) begin
        next_mux_d0_57 = input_word_d[459];
    end else if (sel_d0_57[2:0] == 4) begin
        next_mux_d0_57 = input_word_d[460];
    end else if (sel_d0_57[2:0] == 5) begin
        next_mux_d0_57 = input_word_d[461];
    end else if (sel_d0_57[2:0] == 6) begin
        next_mux_d0_57 = input_word_d[462];
    end else begin
        next_mux_d0_57 = input_word_d[463];
    end

    if (sel_d0_58[2:0] == 0) begin
        next_mux_d0_58 = input_word_d[464];
    end else if (sel_d0_58[2:0] == 1) begin
        next_mux_d0_58 = input_word_d[465];
    end else if (sel_d0_58[2:0] == 2) begin
        next_mux_d0_58 = input_word_d[466];
    end else if (sel_d0_58[2:0] == 3) begin
        next_mux_d0_58 = input_word_d[467];
    end else if (sel_d0_58[2:0] == 4) begin
        next_mux_d0_58 = input_word_d[468];
    end else if (sel_d0_58[2:0] == 5) begin
        next_mux_d0_58 = input_word_d[469];
    end else if (sel_d0_58[2:0] == 6) begin
        next_mux_d0_58 = input_word_d[470];
    end else begin
        next_mux_d0_58 = input_word_d[471];
    end

    if (sel_d0_59[2:0] == 0) begin
        next_mux_d0_59 = input_word_d[472];
    end else if (sel_d0_59[2:0] == 1) begin
        next_mux_d0_59 = input_word_d[473];
    end else if (sel_d0_59[2:0] == 2) begin
        next_mux_d0_59 = input_word_d[474];
    end else if (sel_d0_59[2:0] == 3) begin
        next_mux_d0_59 = input_word_d[475];
    end else if (sel_d0_59[2:0] == 4) begin
        next_mux_d0_59 = input_word_d[476];
    end else if (sel_d0_59[2:0] == 5) begin
        next_mux_d0_59 = input_word_d[477];
    end else if (sel_d0_59[2:0] == 6) begin
        next_mux_d0_59 = input_word_d[478];
    end else begin
        next_mux_d0_59 = input_word_d[479];
    end

    if (sel_d0_60[2:0] == 0) begin
        next_mux_d0_60 = input_word_d[480];
    end else if (sel_d0_60[2:0] == 1) begin
        next_mux_d0_60 = input_word_d[481];
    end else if (sel_d0_60[2:0] == 2) begin
        next_mux_d0_60 = input_word_d[482];
    end else if (sel_d0_60[2:0] == 3) begin
        next_mux_d0_60 = input_word_d[483];
    end else if (sel_d0_60[2:0] == 4) begin
        next_mux_d0_60 = input_word_d[484];
    end else if (sel_d0_60[2:0] == 5) begin
        next_mux_d0_60 = input_word_d[485];
    end else if (sel_d0_60[2:0] == 6) begin
        next_mux_d0_60 = input_word_d[486];
    end else begin
        next_mux_d0_60 = input_word_d[487];
    end

    if (sel_d0_61[2:0] == 0) begin
        next_mux_d0_61 = input_word_d[488];
    end else if (sel_d0_61[2:0] == 1) begin
        next_mux_d0_61 = input_word_d[489];
    end else if (sel_d0_61[2:0] == 2) begin
        next_mux_d0_61 = input_word_d[490];
    end else if (sel_d0_61[2:0] == 3) begin
        next_mux_d0_61 = input_word_d[491];
    end else if (sel_d0_61[2:0] == 4) begin
        next_mux_d0_61 = input_word_d[492];
    end else if (sel_d0_61[2:0] == 5) begin
        next_mux_d0_61 = input_word_d[493];
    end else if (sel_d0_61[2:0] == 6) begin
        next_mux_d0_61 = input_word_d[494];
    end else begin
        next_mux_d0_61 = input_word_d[495];
    end

    if (sel_d0_62[2:0] == 0) begin
        next_mux_d0_62 = input_word_d[496];
    end else if (sel_d0_62[2:0] == 1) begin
        next_mux_d0_62 = input_word_d[497];
    end else if (sel_d0_62[2:0] == 2) begin
        next_mux_d0_62 = input_word_d[498];
    end else if (sel_d0_62[2:0] == 3) begin
        next_mux_d0_62 = input_word_d[499];
    end else if (sel_d0_62[2:0] == 4) begin
        next_mux_d0_62 = input_word_d[500];
    end else if (sel_d0_62[2:0] == 5) begin
        next_mux_d0_62 = input_word_d[501];
    end else if (sel_d0_62[2:0] == 6) begin
        next_mux_d0_62 = input_word_d[502];
    end else begin
        next_mux_d0_62 = input_word_d[503];
    end

    if (sel_d0_63[2:0] == 0) begin
        next_mux_d0_63 = input_word_d[504];
    end else if (sel_d0_63[2:0] == 1) begin
        next_mux_d0_63 = input_word_d[505];
    end else if (sel_d0_63[2:0] == 2) begin
        next_mux_d0_63 = input_word_d[506];
    end else if (sel_d0_63[2:0] == 3) begin
        next_mux_d0_63 = input_word_d[507];
    end else if (sel_d0_63[2:0] == 4) begin
        next_mux_d0_63 = input_word_d[508];
    end else if (sel_d0_63[2:0] == 5) begin
        next_mux_d0_63 = input_word_d[509];
    end else if (sel_d0_63[2:0] == 6) begin
        next_mux_d0_63 = input_word_d[510];
    end else begin
        next_mux_d0_63 = input_word_d[511];
    end

    if (sel_d0_64[2:0] == 0) begin
        next_mux_d0_64 = input_word_d[512];
    end else if (sel_d0_64[2:0] == 1) begin
        next_mux_d0_64 = input_word_d[513];
    end else if (sel_d0_64[2:0] == 2) begin
        next_mux_d0_64 = input_word_d[514];
    end else if (sel_d0_64[2:0] == 3) begin
        next_mux_d0_64 = input_word_d[515];
    end else if (sel_d0_64[2:0] == 4) begin
        next_mux_d0_64 = input_word_d[516];
    end else if (sel_d0_64[2:0] == 5) begin
        next_mux_d0_64 = input_word_d[517];
    end else if (sel_d0_64[2:0] == 6) begin
        next_mux_d0_64 = input_word_d[518];
    end else begin
        next_mux_d0_64 = input_word_d[519];
    end

    if (sel_d0_65[2:0] == 0) begin
        next_mux_d0_65 = input_word_d[520];
    end else if (sel_d0_65[2:0] == 1) begin
        next_mux_d0_65 = input_word_d[521];
    end else if (sel_d0_65[2:0] == 2) begin
        next_mux_d0_65 = input_word_d[522];
    end else if (sel_d0_65[2:0] == 3) begin
        next_mux_d0_65 = input_word_d[523];
    end else if (sel_d0_65[2:0] == 4) begin
        next_mux_d0_65 = input_word_d[524];
    end else if (sel_d0_65[2:0] == 5) begin
        next_mux_d0_65 = input_word_d[525];
    end else if (sel_d0_65[2:0] == 6) begin
        next_mux_d0_65 = input_word_d[526];
    end else begin
        next_mux_d0_65 = input_word_d[527];
    end

    if (sel_d0_66[2:0] == 0) begin
        next_mux_d0_66 = input_word_d[528];
    end else if (sel_d0_66[2:0] == 1) begin
        next_mux_d0_66 = input_word_d[529];
    end else if (sel_d0_66[2:0] == 2) begin
        next_mux_d0_66 = input_word_d[530];
    end else if (sel_d0_66[2:0] == 3) begin
        next_mux_d0_66 = input_word_d[531];
    end else if (sel_d0_66[2:0] == 4) begin
        next_mux_d0_66 = input_word_d[532];
    end else if (sel_d0_66[2:0] == 5) begin
        next_mux_d0_66 = input_word_d[533];
    end else if (sel_d0_66[2:0] == 6) begin
        next_mux_d0_66 = input_word_d[534];
    end else begin
        next_mux_d0_66 = input_word_d[535];
    end

    if (sel_d0_67[2:0] == 0) begin
        next_mux_d0_67 = input_word_d[536];
    end else if (sel_d0_67[2:0] == 1) begin
        next_mux_d0_67 = input_word_d[537];
    end else if (sel_d0_67[2:0] == 2) begin
        next_mux_d0_67 = input_word_d[538];
    end else if (sel_d0_67[2:0] == 3) begin
        next_mux_d0_67 = input_word_d[539];
    end else if (sel_d0_67[2:0] == 4) begin
        next_mux_d0_67 = input_word_d[540];
    end else if (sel_d0_67[2:0] == 5) begin
        next_mux_d0_67 = input_word_d[541];
    end else if (sel_d0_67[2:0] == 6) begin
        next_mux_d0_67 = input_word_d[542];
    end else begin
        next_mux_d0_67 = input_word_d[543];
    end

    if (sel_d0_68[2:0] == 0) begin
        next_mux_d0_68 = input_word_d[544];
    end else if (sel_d0_68[2:0] == 1) begin
        next_mux_d0_68 = input_word_d[545];
    end else if (sel_d0_68[2:0] == 2) begin
        next_mux_d0_68 = input_word_d[546];
    end else if (sel_d0_68[2:0] == 3) begin
        next_mux_d0_68 = input_word_d[547];
    end else if (sel_d0_68[2:0] == 4) begin
        next_mux_d0_68 = input_word_d[548];
    end else if (sel_d0_68[2:0] == 5) begin
        next_mux_d0_68 = input_word_d[549];
    end else if (sel_d0_68[2:0] == 6) begin
        next_mux_d0_68 = input_word_d[550];
    end else begin
        next_mux_d0_68 = input_word_d[551];
    end

    if (sel_d0_69[2:0] == 0) begin
        next_mux_d0_69 = input_word_d[552];
    end else if (sel_d0_69[2:0] == 1) begin
        next_mux_d0_69 = input_word_d[553];
    end else if (sel_d0_69[2:0] == 2) begin
        next_mux_d0_69 = input_word_d[554];
    end else if (sel_d0_69[2:0] == 3) begin
        next_mux_d0_69 = input_word_d[555];
    end else if (sel_d0_69[2:0] == 4) begin
        next_mux_d0_69 = input_word_d[556];
    end else if (sel_d0_69[2:0] == 5) begin
        next_mux_d0_69 = input_word_d[557];
    end else if (sel_d0_69[2:0] == 6) begin
        next_mux_d0_69 = input_word_d[558];
    end else begin
        next_mux_d0_69 = input_word_d[559];
    end

    if (sel_d0_70[2:0] == 0) begin
        next_mux_d0_70 = input_word_d[560];
    end else if (sel_d0_70[2:0] == 1) begin
        next_mux_d0_70 = input_word_d[561];
    end else if (sel_d0_70[2:0] == 2) begin
        next_mux_d0_70 = input_word_d[562];
    end else if (sel_d0_70[2:0] == 3) begin
        next_mux_d0_70 = input_word_d[563];
    end else if (sel_d0_70[2:0] == 4) begin
        next_mux_d0_70 = input_word_d[564];
    end else if (sel_d0_70[2:0] == 5) begin
        next_mux_d0_70 = input_word_d[565];
    end else if (sel_d0_70[2:0] == 6) begin
        next_mux_d0_70 = input_word_d[566];
    end else begin
        next_mux_d0_70 = input_word_d[567];
    end

    if (sel_d0_71[2:0] == 0) begin
        next_mux_d0_71 = input_word_d[568];
    end else if (sel_d0_71[2:0] == 1) begin
        next_mux_d0_71 = input_word_d[569];
    end else if (sel_d0_71[2:0] == 2) begin
        next_mux_d0_71 = input_word_d[570];
    end else if (sel_d0_71[2:0] == 3) begin
        next_mux_d0_71 = input_word_d[571];
    end else if (sel_d0_71[2:0] == 4) begin
        next_mux_d0_71 = input_word_d[572];
    end else if (sel_d0_71[2:0] == 5) begin
        next_mux_d0_71 = input_word_d[573];
    end else if (sel_d0_71[2:0] == 6) begin
        next_mux_d0_71 = input_word_d[574];
    end else begin
        next_mux_d0_71 = input_word_d[575];
    end

    if (sel_d0_72[2:0] == 0) begin
        next_mux_d0_72 = input_word_d[576];
    end else if (sel_d0_72[2:0] == 1) begin
        next_mux_d0_72 = input_word_d[577];
    end else if (sel_d0_72[2:0] == 2) begin
        next_mux_d0_72 = input_word_d[578];
    end else if (sel_d0_72[2:0] == 3) begin
        next_mux_d0_72 = input_word_d[579];
    end else if (sel_d0_72[2:0] == 4) begin
        next_mux_d0_72 = input_word_d[580];
    end else if (sel_d0_72[2:0] == 5) begin
        next_mux_d0_72 = input_word_d[581];
    end else if (sel_d0_72[2:0] == 6) begin
        next_mux_d0_72 = input_word_d[582];
    end else begin
        next_mux_d0_72 = input_word_d[583];
    end

    if (sel_d0_73[2:0] == 0) begin
        next_mux_d0_73 = input_word_d[584];
    end else if (sel_d0_73[2:0] == 1) begin
        next_mux_d0_73 = input_word_d[585];
    end else if (sel_d0_73[2:0] == 2) begin
        next_mux_d0_73 = input_word_d[586];
    end else if (sel_d0_73[2:0] == 3) begin
        next_mux_d0_73 = input_word_d[587];
    end else if (sel_d0_73[2:0] == 4) begin
        next_mux_d0_73 = input_word_d[588];
    end else if (sel_d0_73[2:0] == 5) begin
        next_mux_d0_73 = input_word_d[589];
    end else if (sel_d0_73[2:0] == 6) begin
        next_mux_d0_73 = input_word_d[590];
    end else begin
        next_mux_d0_73 = input_word_d[591];
    end

    if (sel_d0_74[2:0] == 0) begin
        next_mux_d0_74 = input_word_d[592];
    end else if (sel_d0_74[2:0] == 1) begin
        next_mux_d0_74 = input_word_d[593];
    end else if (sel_d0_74[2:0] == 2) begin
        next_mux_d0_74 = input_word_d[594];
    end else if (sel_d0_74[2:0] == 3) begin
        next_mux_d0_74 = input_word_d[595];
    end else if (sel_d0_74[2:0] == 4) begin
        next_mux_d0_74 = input_word_d[596];
    end else if (sel_d0_74[2:0] == 5) begin
        next_mux_d0_74 = input_word_d[597];
    end else if (sel_d0_74[2:0] == 6) begin
        next_mux_d0_74 = input_word_d[598];
    end else begin
        next_mux_d0_74 = input_word_d[599];
    end

    if (sel_d0_75[2:0] == 0) begin
        next_mux_d0_75 = input_word_d[600];
    end else if (sel_d0_75[2:0] == 1) begin
        next_mux_d0_75 = input_word_d[601];
    end else if (sel_d0_75[2:0] == 2) begin
        next_mux_d0_75 = input_word_d[602];
    end else if (sel_d0_75[2:0] == 3) begin
        next_mux_d0_75 = input_word_d[603];
    end else if (sel_d0_75[2:0] == 4) begin
        next_mux_d0_75 = input_word_d[604];
    end else if (sel_d0_75[2:0] == 5) begin
        next_mux_d0_75 = input_word_d[605];
    end else if (sel_d0_75[2:0] == 6) begin
        next_mux_d0_75 = input_word_d[606];
    end else begin
        next_mux_d0_75 = input_word_d[607];
    end

    if (sel_d0_76[2:0] == 0) begin
        next_mux_d0_76 = input_word_d[608];
    end else if (sel_d0_76[2:0] == 1) begin
        next_mux_d0_76 = input_word_d[609];
    end else if (sel_d0_76[2:0] == 2) begin
        next_mux_d0_76 = input_word_d[610];
    end else if (sel_d0_76[2:0] == 3) begin
        next_mux_d0_76 = input_word_d[611];
    end else if (sel_d0_76[2:0] == 4) begin
        next_mux_d0_76 = input_word_d[612];
    end else if (sel_d0_76[2:0] == 5) begin
        next_mux_d0_76 = input_word_d[613];
    end else if (sel_d0_76[2:0] == 6) begin
        next_mux_d0_76 = input_word_d[614];
    end else begin
        next_mux_d0_76 = input_word_d[615];
    end

    if (sel_d0_77[2:0] == 0) begin
        next_mux_d0_77 = input_word_d[616];
    end else if (sel_d0_77[2:0] == 1) begin
        next_mux_d0_77 = input_word_d[617];
    end else if (sel_d0_77[2:0] == 2) begin
        next_mux_d0_77 = input_word_d[618];
    end else if (sel_d0_77[2:0] == 3) begin
        next_mux_d0_77 = input_word_d[619];
    end else if (sel_d0_77[2:0] == 4) begin
        next_mux_d0_77 = input_word_d[620];
    end else if (sel_d0_77[2:0] == 5) begin
        next_mux_d0_77 = input_word_d[621];
    end else if (sel_d0_77[2:0] == 6) begin
        next_mux_d0_77 = input_word_d[622];
    end else begin
        next_mux_d0_77 = input_word_d[623];
    end

    if (sel_d0_78[2:0] == 0) begin
        next_mux_d0_78 = input_word_d[624];
    end else if (sel_d0_78[2:0] == 1) begin
        next_mux_d0_78 = input_word_d[625];
    end else if (sel_d0_78[2:0] == 2) begin
        next_mux_d0_78 = input_word_d[626];
    end else if (sel_d0_78[2:0] == 3) begin
        next_mux_d0_78 = input_word_d[627];
    end else if (sel_d0_78[2:0] == 4) begin
        next_mux_d0_78 = input_word_d[628];
    end else if (sel_d0_78[2:0] == 5) begin
        next_mux_d0_78 = input_word_d[629];
    end else if (sel_d0_78[2:0] == 6) begin
        next_mux_d0_78 = input_word_d[630];
    end else begin
        next_mux_d0_78 = input_word_d[631];
    end

    if (sel_d0_79[2:0] == 0) begin
        next_mux_d0_79 = input_word_d[632];
    end else if (sel_d0_79[2:0] == 1) begin
        next_mux_d0_79 = input_word_d[633];
    end else if (sel_d0_79[2:0] == 2) begin
        next_mux_d0_79 = input_word_d[634];
    end else if (sel_d0_79[2:0] == 3) begin
        next_mux_d0_79 = input_word_d[635];
    end else if (sel_d0_79[2:0] == 4) begin
        next_mux_d0_79 = input_word_d[636];
    end else if (sel_d0_79[2:0] == 5) begin
        next_mux_d0_79 = input_word_d[637];
    end else if (sel_d0_79[2:0] == 6) begin
        next_mux_d0_79 = input_word_d[638];
    end else begin
        next_mux_d0_79 = input_word_d[639];
    end

    if (sel_d0_80[2:0] == 0) begin
        next_mux_d0_80 = input_word_d[640];
    end else if (sel_d0_80[2:0] == 1) begin
        next_mux_d0_80 = input_word_d[641];
    end else if (sel_d0_80[2:0] == 2) begin
        next_mux_d0_80 = input_word_d[642];
    end else if (sel_d0_80[2:0] == 3) begin
        next_mux_d0_80 = input_word_d[643];
    end else if (sel_d0_80[2:0] == 4) begin
        next_mux_d0_80 = input_word_d[644];
    end else if (sel_d0_80[2:0] == 5) begin
        next_mux_d0_80 = input_word_d[645];
    end else if (sel_d0_80[2:0] == 6) begin
        next_mux_d0_80 = input_word_d[646];
    end else begin
        next_mux_d0_80 = input_word_d[647];
    end

    if (sel_d0_81[2:0] == 0) begin
        next_mux_d0_81 = input_word_d[648];
    end else if (sel_d0_81[2:0] == 1) begin
        next_mux_d0_81 = input_word_d[649];
    end else if (sel_d0_81[2:0] == 2) begin
        next_mux_d0_81 = input_word_d[650];
    end else if (sel_d0_81[2:0] == 3) begin
        next_mux_d0_81 = input_word_d[651];
    end else if (sel_d0_81[2:0] == 4) begin
        next_mux_d0_81 = input_word_d[652];
    end else if (sel_d0_81[2:0] == 5) begin
        next_mux_d0_81 = input_word_d[653];
    end else if (sel_d0_81[2:0] == 6) begin
        next_mux_d0_81 = input_word_d[654];
    end else begin
        next_mux_d0_81 = input_word_d[655];
    end

    if (sel_d0_82[2:0] == 0) begin
        next_mux_d0_82 = input_word_d[656];
    end else if (sel_d0_82[2:0] == 1) begin
        next_mux_d0_82 = input_word_d[657];
    end else if (sel_d0_82[2:0] == 2) begin
        next_mux_d0_82 = input_word_d[658];
    end else if (sel_d0_82[2:0] == 3) begin
        next_mux_d0_82 = input_word_d[659];
    end else if (sel_d0_82[2:0] == 4) begin
        next_mux_d0_82 = input_word_d[660];
    end else if (sel_d0_82[2:0] == 5) begin
        next_mux_d0_82 = input_word_d[661];
    end else if (sel_d0_82[2:0] == 6) begin
        next_mux_d0_82 = input_word_d[662];
    end else begin
        next_mux_d0_82 = input_word_d[663];
    end

    if (sel_d0_83[2:0] == 0) begin
        next_mux_d0_83 = input_word_d[664];
    end else if (sel_d0_83[2:0] == 1) begin
        next_mux_d0_83 = input_word_d[665];
    end else if (sel_d0_83[2:0] == 2) begin
        next_mux_d0_83 = input_word_d[666];
    end else if (sel_d0_83[2:0] == 3) begin
        next_mux_d0_83 = input_word_d[667];
    end else if (sel_d0_83[2:0] == 4) begin
        next_mux_d0_83 = input_word_d[668];
    end else if (sel_d0_83[2:0] == 5) begin
        next_mux_d0_83 = input_word_d[669];
    end else if (sel_d0_83[2:0] == 6) begin
        next_mux_d0_83 = input_word_d[670];
    end else begin
        next_mux_d0_83 = input_word_d[671];
    end

    if (sel_d0_84[2:0] == 0) begin
        next_mux_d0_84 = input_word_d[672];
    end else if (sel_d0_84[2:0] == 1) begin
        next_mux_d0_84 = input_word_d[673];
    end else if (sel_d0_84[2:0] == 2) begin
        next_mux_d0_84 = input_word_d[674];
    end else if (sel_d0_84[2:0] == 3) begin
        next_mux_d0_84 = input_word_d[675];
    end else if (sel_d0_84[2:0] == 4) begin
        next_mux_d0_84 = input_word_d[676];
    end else if (sel_d0_84[2:0] == 5) begin
        next_mux_d0_84 = input_word_d[677];
    end else if (sel_d0_84[2:0] == 6) begin
        next_mux_d0_84 = input_word_d[678];
    end else begin
        next_mux_d0_84 = input_word_d[679];
    end

    if (sel_d0_85[2:0] == 0) begin
        next_mux_d0_85 = input_word_d[680];
    end else if (sel_d0_85[2:0] == 1) begin
        next_mux_d0_85 = input_word_d[681];
    end else if (sel_d0_85[2:0] == 2) begin
        next_mux_d0_85 = input_word_d[682];
    end else if (sel_d0_85[2:0] == 3) begin
        next_mux_d0_85 = input_word_d[683];
    end else if (sel_d0_85[2:0] == 4) begin
        next_mux_d0_85 = input_word_d[684];
    end else if (sel_d0_85[2:0] == 5) begin
        next_mux_d0_85 = input_word_d[685];
    end else if (sel_d0_85[2:0] == 6) begin
        next_mux_d0_85 = input_word_d[686];
    end else begin
        next_mux_d0_85 = input_word_d[687];
    end

    if (sel_d0_86[2:0] == 0) begin
        next_mux_d0_86 = input_word_d[688];
    end else if (sel_d0_86[2:0] == 1) begin
        next_mux_d0_86 = input_word_d[689];
    end else if (sel_d0_86[2:0] == 2) begin
        next_mux_d0_86 = input_word_d[690];
    end else if (sel_d0_86[2:0] == 3) begin
        next_mux_d0_86 = input_word_d[691];
    end else if (sel_d0_86[2:0] == 4) begin
        next_mux_d0_86 = input_word_d[692];
    end else if (sel_d0_86[2:0] == 5) begin
        next_mux_d0_86 = input_word_d[693];
    end else if (sel_d0_86[2:0] == 6) begin
        next_mux_d0_86 = input_word_d[694];
    end else begin
        next_mux_d0_86 = input_word_d[695];
    end

    if (sel_d0_87[2:0] == 0) begin
        next_mux_d0_87 = input_word_d[696];
    end else if (sel_d0_87[2:0] == 1) begin
        next_mux_d0_87 = input_word_d[697];
    end else if (sel_d0_87[2:0] == 2) begin
        next_mux_d0_87 = input_word_d[698];
    end else if (sel_d0_87[2:0] == 3) begin
        next_mux_d0_87 = input_word_d[699];
    end else if (sel_d0_87[2:0] == 4) begin
        next_mux_d0_87 = input_word_d[700];
    end else if (sel_d0_87[2:0] == 5) begin
        next_mux_d0_87 = input_word_d[701];
    end else if (sel_d0_87[2:0] == 6) begin
        next_mux_d0_87 = input_word_d[702];
    end else begin
        next_mux_d0_87 = input_word_d[703];
    end

    if (sel_d0_88[2:0] == 0) begin
        next_mux_d0_88 = input_word_d[704];
    end else if (sel_d0_88[2:0] == 1) begin
        next_mux_d0_88 = input_word_d[705];
    end else if (sel_d0_88[2:0] == 2) begin
        next_mux_d0_88 = input_word_d[706];
    end else if (sel_d0_88[2:0] == 3) begin
        next_mux_d0_88 = input_word_d[707];
    end else if (sel_d0_88[2:0] == 4) begin
        next_mux_d0_88 = input_word_d[708];
    end else if (sel_d0_88[2:0] == 5) begin
        next_mux_d0_88 = input_word_d[709];
    end else if (sel_d0_88[2:0] == 6) begin
        next_mux_d0_88 = input_word_d[710];
    end else begin
        next_mux_d0_88 = input_word_d[711];
    end

    if (sel_d0_89[2:0] == 0) begin
        next_mux_d0_89 = input_word_d[712];
    end else if (sel_d0_89[2:0] == 1) begin
        next_mux_d0_89 = input_word_d[713];
    end else if (sel_d0_89[2:0] == 2) begin
        next_mux_d0_89 = input_word_d[714];
    end else if (sel_d0_89[2:0] == 3) begin
        next_mux_d0_89 = input_word_d[715];
    end else if (sel_d0_89[2:0] == 4) begin
        next_mux_d0_89 = input_word_d[716];
    end else if (sel_d0_89[2:0] == 5) begin
        next_mux_d0_89 = input_word_d[717];
    end else if (sel_d0_89[2:0] == 6) begin
        next_mux_d0_89 = input_word_d[718];
    end else begin
        next_mux_d0_89 = input_word_d[719];
    end

    if (sel_d0_90[2:0] == 0) begin
        next_mux_d0_90 = input_word_d[720];
    end else if (sel_d0_90[2:0] == 1) begin
        next_mux_d0_90 = input_word_d[721];
    end else if (sel_d0_90[2:0] == 2) begin
        next_mux_d0_90 = input_word_d[722];
    end else if (sel_d0_90[2:0] == 3) begin
        next_mux_d0_90 = input_word_d[723];
    end else if (sel_d0_90[2:0] == 4) begin
        next_mux_d0_90 = input_word_d[724];
    end else if (sel_d0_90[2:0] == 5) begin
        next_mux_d0_90 = input_word_d[725];
    end else if (sel_d0_90[2:0] == 6) begin
        next_mux_d0_90 = input_word_d[726];
    end else begin
        next_mux_d0_90 = input_word_d[727];
    end

    if (sel_d0_91[2:0] == 0) begin
        next_mux_d0_91 = input_word_d[728];
    end else if (sel_d0_91[2:0] == 1) begin
        next_mux_d0_91 = input_word_d[729];
    end else if (sel_d0_91[2:0] == 2) begin
        next_mux_d0_91 = input_word_d[730];
    end else if (sel_d0_91[2:0] == 3) begin
        next_mux_d0_91 = input_word_d[731];
    end else if (sel_d0_91[2:0] == 4) begin
        next_mux_d0_91 = input_word_d[732];
    end else if (sel_d0_91[2:0] == 5) begin
        next_mux_d0_91 = input_word_d[733];
    end else if (sel_d0_91[2:0] == 6) begin
        next_mux_d0_91 = input_word_d[734];
    end else begin
        next_mux_d0_91 = input_word_d[735];
    end

    if (sel_d0_92[2:0] == 0) begin
        next_mux_d0_92 = input_word_d[736];
    end else if (sel_d0_92[2:0] == 1) begin
        next_mux_d0_92 = input_word_d[737];
    end else if (sel_d0_92[2:0] == 2) begin
        next_mux_d0_92 = input_word_d[738];
    end else if (sel_d0_92[2:0] == 3) begin
        next_mux_d0_92 = input_word_d[739];
    end else if (sel_d0_92[2:0] == 4) begin
        next_mux_d0_92 = input_word_d[740];
    end else if (sel_d0_92[2:0] == 5) begin
        next_mux_d0_92 = input_word_d[741];
    end else if (sel_d0_92[2:0] == 6) begin
        next_mux_d0_92 = input_word_d[742];
    end else begin
        next_mux_d0_92 = input_word_d[743];
    end

    if (sel_d0_93[2:0] == 0) begin
        next_mux_d0_93 = input_word_d[744];
    end else if (sel_d0_93[2:0] == 1) begin
        next_mux_d0_93 = input_word_d[745];
    end else if (sel_d0_93[2:0] == 2) begin
        next_mux_d0_93 = input_word_d[746];
    end else if (sel_d0_93[2:0] == 3) begin
        next_mux_d0_93 = input_word_d[747];
    end else if (sel_d0_93[2:0] == 4) begin
        next_mux_d0_93 = input_word_d[748];
    end else if (sel_d0_93[2:0] == 5) begin
        next_mux_d0_93 = input_word_d[749];
    end else if (sel_d0_93[2:0] == 6) begin
        next_mux_d0_93 = input_word_d[750];
    end else begin
        next_mux_d0_93 = input_word_d[751];
    end

    if (sel_d0_94[2:0] == 0) begin
        next_mux_d0_94 = input_word_d[752];
    end else if (sel_d0_94[2:0] == 1) begin
        next_mux_d0_94 = input_word_d[753];
    end else if (sel_d0_94[2:0] == 2) begin
        next_mux_d0_94 = input_word_d[754];
    end else if (sel_d0_94[2:0] == 3) begin
        next_mux_d0_94 = input_word_d[755];
    end else if (sel_d0_94[2:0] == 4) begin
        next_mux_d0_94 = input_word_d[756];
    end else if (sel_d0_94[2:0] == 5) begin
        next_mux_d0_94 = input_word_d[757];
    end else if (sel_d0_94[2:0] == 6) begin
        next_mux_d0_94 = input_word_d[758];
    end else begin
        next_mux_d0_94 = input_word_d[759];
    end

    if (sel_d0_95[2:0] == 0) begin
        next_mux_d0_95 = input_word_d[760];
    end else if (sel_d0_95[2:0] == 1) begin
        next_mux_d0_95 = input_word_d[761];
    end else if (sel_d0_95[2:0] == 2) begin
        next_mux_d0_95 = input_word_d[762];
    end else if (sel_d0_95[2:0] == 3) begin
        next_mux_d0_95 = input_word_d[763];
    end else if (sel_d0_95[2:0] == 4) begin
        next_mux_d0_95 = input_word_d[764];
    end else if (sel_d0_95[2:0] == 5) begin
        next_mux_d0_95 = input_word_d[765];
    end else if (sel_d0_95[2:0] == 6) begin
        next_mux_d0_95 = input_word_d[766];
    end else begin
        next_mux_d0_95 = input_word_d[767];
    end

    if (sel_d0_96[2:0] == 0) begin
        next_mux_d0_96 = input_word_d[768];
    end else if (sel_d0_96[2:0] == 1) begin
        next_mux_d0_96 = input_word_d[769];
    end else if (sel_d0_96[2:0] == 2) begin
        next_mux_d0_96 = input_word_d[770];
    end else if (sel_d0_96[2:0] == 3) begin
        next_mux_d0_96 = input_word_d[771];
    end else if (sel_d0_96[2:0] == 4) begin
        next_mux_d0_96 = input_word_d[772];
    end else if (sel_d0_96[2:0] == 5) begin
        next_mux_d0_96 = input_word_d[773];
    end else if (sel_d0_96[2:0] == 6) begin
        next_mux_d0_96 = input_word_d[774];
    end else begin
        next_mux_d0_96 = input_word_d[775];
    end

    if (sel_d0_97[2:0] == 0) begin
        next_mux_d0_97 = input_word_d[776];
    end else if (sel_d0_97[2:0] == 1) begin
        next_mux_d0_97 = input_word_d[777];
    end else if (sel_d0_97[2:0] == 2) begin
        next_mux_d0_97 = input_word_d[778];
    end else if (sel_d0_97[2:0] == 3) begin
        next_mux_d0_97 = input_word_d[779];
    end else if (sel_d0_97[2:0] == 4) begin
        next_mux_d0_97 = input_word_d[780];
    end else if (sel_d0_97[2:0] == 5) begin
        next_mux_d0_97 = input_word_d[781];
    end else if (sel_d0_97[2:0] == 6) begin
        next_mux_d0_97 = input_word_d[782];
    end else begin
        next_mux_d0_97 = input_word_d[783];
    end

    if (sel_d0_98[2:0] == 0) begin
        next_mux_d0_98 = input_word_d[784];
    end else if (sel_d0_98[2:0] == 1) begin
        next_mux_d0_98 = input_word_d[785];
    end else if (sel_d0_98[2:0] == 2) begin
        next_mux_d0_98 = input_word_d[786];
    end else if (sel_d0_98[2:0] == 3) begin
        next_mux_d0_98 = input_word_d[787];
    end else if (sel_d0_98[2:0] == 4) begin
        next_mux_d0_98 = input_word_d[788];
    end else if (sel_d0_98[2:0] == 5) begin
        next_mux_d0_98 = input_word_d[789];
    end else if (sel_d0_98[2:0] == 6) begin
        next_mux_d0_98 = input_word_d[790];
    end else begin
        next_mux_d0_98 = input_word_d[791];
    end

    if (sel_d0_99[2:0] == 0) begin
        next_mux_d0_99 = input_word_d[792];
    end else if (sel_d0_99[2:0] == 1) begin
        next_mux_d0_99 = input_word_d[793];
    end else if (sel_d0_99[2:0] == 2) begin
        next_mux_d0_99 = input_word_d[794];
    end else if (sel_d0_99[2:0] == 3) begin
        next_mux_d0_99 = input_word_d[795];
    end else if (sel_d0_99[2:0] == 4) begin
        next_mux_d0_99 = input_word_d[796];
    end else if (sel_d0_99[2:0] == 5) begin
        next_mux_d0_99 = input_word_d[797];
    end else if (sel_d0_99[2:0] == 6) begin
        next_mux_d0_99 = input_word_d[798];
    end else begin
        next_mux_d0_99 = input_word_d[799];
    end

    if (sel_d0_100[2:0] == 0) begin
        next_mux_d0_100 = input_word_d[800];
    end else if (sel_d0_100[2:0] == 1) begin
        next_mux_d0_100 = input_word_d[801];
    end else if (sel_d0_100[2:0] == 2) begin
        next_mux_d0_100 = input_word_d[802];
    end else if (sel_d0_100[2:0] == 3) begin
        next_mux_d0_100 = input_word_d[803];
    end else if (sel_d0_100[2:0] == 4) begin
        next_mux_d0_100 = input_word_d[804];
    end else if (sel_d0_100[2:0] == 5) begin
        next_mux_d0_100 = input_word_d[805];
    end else if (sel_d0_100[2:0] == 6) begin
        next_mux_d0_100 = input_word_d[806];
    end else begin
        next_mux_d0_100 = input_word_d[807];
    end

    if (sel_d0_101[2:0] == 0) begin
        next_mux_d0_101 = input_word_d[808];
    end else if (sel_d0_101[2:0] == 1) begin
        next_mux_d0_101 = input_word_d[809];
    end else if (sel_d0_101[2:0] == 2) begin
        next_mux_d0_101 = input_word_d[810];
    end else if (sel_d0_101[2:0] == 3) begin
        next_mux_d0_101 = input_word_d[811];
    end else if (sel_d0_101[2:0] == 4) begin
        next_mux_d0_101 = input_word_d[812];
    end else if (sel_d0_101[2:0] == 5) begin
        next_mux_d0_101 = input_word_d[813];
    end else if (sel_d0_101[2:0] == 6) begin
        next_mux_d0_101 = input_word_d[814];
    end else begin
        next_mux_d0_101 = input_word_d[815];
    end

    if (sel_d0_102[2:0] == 0) begin
        next_mux_d0_102 = input_word_d[816];
    end else if (sel_d0_102[2:0] == 1) begin
        next_mux_d0_102 = input_word_d[817];
    end else if (sel_d0_102[2:0] == 2) begin
        next_mux_d0_102 = input_word_d[818];
    end else if (sel_d0_102[2:0] == 3) begin
        next_mux_d0_102 = input_word_d[819];
    end else if (sel_d0_102[2:0] == 4) begin
        next_mux_d0_102 = input_word_d[820];
    end else if (sel_d0_102[2:0] == 5) begin
        next_mux_d0_102 = input_word_d[821];
    end else if (sel_d0_102[2:0] == 6) begin
        next_mux_d0_102 = input_word_d[822];
    end else begin
        next_mux_d0_102 = input_word_d[823];
    end

    if (sel_d0_103[2:0] == 0) begin
        next_mux_d0_103 = input_word_d[824];
    end else if (sel_d0_103[2:0] == 1) begin
        next_mux_d0_103 = input_word_d[825];
    end else if (sel_d0_103[2:0] == 2) begin
        next_mux_d0_103 = input_word_d[826];
    end else if (sel_d0_103[2:0] == 3) begin
        next_mux_d0_103 = input_word_d[827];
    end else if (sel_d0_103[2:0] == 4) begin
        next_mux_d0_103 = input_word_d[828];
    end else if (sel_d0_103[2:0] == 5) begin
        next_mux_d0_103 = input_word_d[829];
    end else if (sel_d0_103[2:0] == 6) begin
        next_mux_d0_103 = input_word_d[830];
    end else begin
        next_mux_d0_103 = input_word_d[831];
    end

    if (sel_d0_104[2:0] == 0) begin
        next_mux_d0_104 = input_word_d[832];
    end else if (sel_d0_104[2:0] == 1) begin
        next_mux_d0_104 = input_word_d[833];
    end else if (sel_d0_104[2:0] == 2) begin
        next_mux_d0_104 = input_word_d[834];
    end else if (sel_d0_104[2:0] == 3) begin
        next_mux_d0_104 = input_word_d[835];
    end else if (sel_d0_104[2:0] == 4) begin
        next_mux_d0_104 = input_word_d[836];
    end else if (sel_d0_104[2:0] == 5) begin
        next_mux_d0_104 = input_word_d[837];
    end else if (sel_d0_104[2:0] == 6) begin
        next_mux_d0_104 = input_word_d[838];
    end else begin
        next_mux_d0_104 = input_word_d[839];
    end

    if (sel_d0_105[2:0] == 0) begin
        next_mux_d0_105 = input_word_d[840];
    end else if (sel_d0_105[2:0] == 1) begin
        next_mux_d0_105 = input_word_d[841];
    end else if (sel_d0_105[2:0] == 2) begin
        next_mux_d0_105 = input_word_d[842];
    end else if (sel_d0_105[2:0] == 3) begin
        next_mux_d0_105 = input_word_d[843];
    end else if (sel_d0_105[2:0] == 4) begin
        next_mux_d0_105 = input_word_d[844];
    end else if (sel_d0_105[2:0] == 5) begin
        next_mux_d0_105 = input_word_d[845];
    end else if (sel_d0_105[2:0] == 6) begin
        next_mux_d0_105 = input_word_d[846];
    end else begin
        next_mux_d0_105 = input_word_d[847];
    end

    if (sel_d0_106[2:0] == 0) begin
        next_mux_d0_106 = input_word_d[848];
    end else if (sel_d0_106[2:0] == 1) begin
        next_mux_d0_106 = input_word_d[849];
    end else if (sel_d0_106[2:0] == 2) begin
        next_mux_d0_106 = input_word_d[850];
    end else if (sel_d0_106[2:0] == 3) begin
        next_mux_d0_106 = input_word_d[851];
    end else if (sel_d0_106[2:0] == 4) begin
        next_mux_d0_106 = input_word_d[852];
    end else if (sel_d0_106[2:0] == 5) begin
        next_mux_d0_106 = input_word_d[853];
    end else if (sel_d0_106[2:0] == 6) begin
        next_mux_d0_106 = input_word_d[854];
    end else begin
        next_mux_d0_106 = input_word_d[855];
    end

    if (sel_d0_107[2:0] == 0) begin
        next_mux_d0_107 = input_word_d[856];
    end else if (sel_d0_107[2:0] == 1) begin
        next_mux_d0_107 = input_word_d[857];
    end else if (sel_d0_107[2:0] == 2) begin
        next_mux_d0_107 = input_word_d[858];
    end else if (sel_d0_107[2:0] == 3) begin
        next_mux_d0_107 = input_word_d[859];
    end else if (sel_d0_107[2:0] == 4) begin
        next_mux_d0_107 = input_word_d[860];
    end else if (sel_d0_107[2:0] == 5) begin
        next_mux_d0_107 = input_word_d[861];
    end else if (sel_d0_107[2:0] == 6) begin
        next_mux_d0_107 = input_word_d[862];
    end else begin
        next_mux_d0_107 = input_word_d[863];
    end

    if (sel_d0_108[2:0] == 0) begin
        next_mux_d0_108 = input_word_d[864];
    end else if (sel_d0_108[2:0] == 1) begin
        next_mux_d0_108 = input_word_d[865];
    end else if (sel_d0_108[2:0] == 2) begin
        next_mux_d0_108 = input_word_d[866];
    end else if (sel_d0_108[2:0] == 3) begin
        next_mux_d0_108 = input_word_d[867];
    end else if (sel_d0_108[2:0] == 4) begin
        next_mux_d0_108 = input_word_d[868];
    end else if (sel_d0_108[2:0] == 5) begin
        next_mux_d0_108 = input_word_d[869];
    end else if (sel_d0_108[2:0] == 6) begin
        next_mux_d0_108 = input_word_d[870];
    end else begin
        next_mux_d0_108 = input_word_d[871];
    end

    if (sel_d0_109[2:0] == 0) begin
        next_mux_d0_109 = input_word_d[872];
    end else if (sel_d0_109[2:0] == 1) begin
        next_mux_d0_109 = input_word_d[873];
    end else if (sel_d0_109[2:0] == 2) begin
        next_mux_d0_109 = input_word_d[874];
    end else if (sel_d0_109[2:0] == 3) begin
        next_mux_d0_109 = input_word_d[875];
    end else if (sel_d0_109[2:0] == 4) begin
        next_mux_d0_109 = input_word_d[876];
    end else if (sel_d0_109[2:0] == 5) begin
        next_mux_d0_109 = input_word_d[877];
    end else if (sel_d0_109[2:0] == 6) begin
        next_mux_d0_109 = input_word_d[878];
    end else begin
        next_mux_d0_109 = input_word_d[879];
    end

    if (sel_d0_110[2:0] == 0) begin
        next_mux_d0_110 = input_word_d[880];
    end else if (sel_d0_110[2:0] == 1) begin
        next_mux_d0_110 = input_word_d[881];
    end else if (sel_d0_110[2:0] == 2) begin
        next_mux_d0_110 = input_word_d[882];
    end else if (sel_d0_110[2:0] == 3) begin
        next_mux_d0_110 = input_word_d[883];
    end else if (sel_d0_110[2:0] == 4) begin
        next_mux_d0_110 = input_word_d[884];
    end else if (sel_d0_110[2:0] == 5) begin
        next_mux_d0_110 = input_word_d[885];
    end else if (sel_d0_110[2:0] == 6) begin
        next_mux_d0_110 = input_word_d[886];
    end else begin
        next_mux_d0_110 = input_word_d[887];
    end

    if (sel_d0_111[2:0] == 0) begin
        next_mux_d0_111 = input_word_d[888];
    end else if (sel_d0_111[2:0] == 1) begin
        next_mux_d0_111 = input_word_d[889];
    end else if (sel_d0_111[2:0] == 2) begin
        next_mux_d0_111 = input_word_d[890];
    end else if (sel_d0_111[2:0] == 3) begin
        next_mux_d0_111 = input_word_d[891];
    end else if (sel_d0_111[2:0] == 4) begin
        next_mux_d0_111 = input_word_d[892];
    end else if (sel_d0_111[2:0] == 5) begin
        next_mux_d0_111 = input_word_d[893];
    end else if (sel_d0_111[2:0] == 6) begin
        next_mux_d0_111 = input_word_d[894];
    end else begin
        next_mux_d0_111 = input_word_d[895];
    end

    if (sel_d0_112[2:0] == 0) begin
        next_mux_d0_112 = input_word_d[896];
    end else if (sel_d0_112[2:0] == 1) begin
        next_mux_d0_112 = input_word_d[897];
    end else if (sel_d0_112[2:0] == 2) begin
        next_mux_d0_112 = input_word_d[898];
    end else if (sel_d0_112[2:0] == 3) begin
        next_mux_d0_112 = input_word_d[899];
    end else if (sel_d0_112[2:0] == 4) begin
        next_mux_d0_112 = input_word_d[900];
    end else if (sel_d0_112[2:0] == 5) begin
        next_mux_d0_112 = input_word_d[901];
    end else if (sel_d0_112[2:0] == 6) begin
        next_mux_d0_112 = input_word_d[902];
    end else begin
        next_mux_d0_112 = input_word_d[903];
    end

    if (sel_d0_113[2:0] == 0) begin
        next_mux_d0_113 = input_word_d[904];
    end else if (sel_d0_113[2:0] == 1) begin
        next_mux_d0_113 = input_word_d[905];
    end else if (sel_d0_113[2:0] == 2) begin
        next_mux_d0_113 = input_word_d[906];
    end else if (sel_d0_113[2:0] == 3) begin
        next_mux_d0_113 = input_word_d[907];
    end else if (sel_d0_113[2:0] == 4) begin
        next_mux_d0_113 = input_word_d[908];
    end else if (sel_d0_113[2:0] == 5) begin
        next_mux_d0_113 = input_word_d[909];
    end else if (sel_d0_113[2:0] == 6) begin
        next_mux_d0_113 = input_word_d[910];
    end else begin
        next_mux_d0_113 = input_word_d[911];
    end

    if (sel_d0_114[2:0] == 0) begin
        next_mux_d0_114 = input_word_d[912];
    end else if (sel_d0_114[2:0] == 1) begin
        next_mux_d0_114 = input_word_d[913];
    end else if (sel_d0_114[2:0] == 2) begin
        next_mux_d0_114 = input_word_d[914];
    end else if (sel_d0_114[2:0] == 3) begin
        next_mux_d0_114 = input_word_d[915];
    end else if (sel_d0_114[2:0] == 4) begin
        next_mux_d0_114 = input_word_d[916];
    end else if (sel_d0_114[2:0] == 5) begin
        next_mux_d0_114 = input_word_d[917];
    end else if (sel_d0_114[2:0] == 6) begin
        next_mux_d0_114 = input_word_d[918];
    end else begin
        next_mux_d0_114 = input_word_d[919];
    end

    if (sel_d0_115[2:0] == 0) begin
        next_mux_d0_115 = input_word_d[920];
    end else if (sel_d0_115[2:0] == 1) begin
        next_mux_d0_115 = input_word_d[921];
    end else if (sel_d0_115[2:0] == 2) begin
        next_mux_d0_115 = input_word_d[922];
    end else if (sel_d0_115[2:0] == 3) begin
        next_mux_d0_115 = input_word_d[923];
    end else if (sel_d0_115[2:0] == 4) begin
        next_mux_d0_115 = input_word_d[924];
    end else if (sel_d0_115[2:0] == 5) begin
        next_mux_d0_115 = input_word_d[925];
    end else if (sel_d0_115[2:0] == 6) begin
        next_mux_d0_115 = input_word_d[926];
    end else begin
        next_mux_d0_115 = input_word_d[927];
    end

    if (sel_d0_116[2:0] == 0) begin
        next_mux_d0_116 = input_word_d[928];
    end else if (sel_d0_116[2:0] == 1) begin
        next_mux_d0_116 = input_word_d[929];
    end else if (sel_d0_116[2:0] == 2) begin
        next_mux_d0_116 = input_word_d[930];
    end else if (sel_d0_116[2:0] == 3) begin
        next_mux_d0_116 = input_word_d[931];
    end else if (sel_d0_116[2:0] == 4) begin
        next_mux_d0_116 = input_word_d[932];
    end else if (sel_d0_116[2:0] == 5) begin
        next_mux_d0_116 = input_word_d[933];
    end else if (sel_d0_116[2:0] == 6) begin
        next_mux_d0_116 = input_word_d[934];
    end else begin
        next_mux_d0_116 = input_word_d[935];
    end

    if (sel_d0_117[2:0] == 0) begin
        next_mux_d0_117 = input_word_d[936];
    end else if (sel_d0_117[2:0] == 1) begin
        next_mux_d0_117 = input_word_d[937];
    end else if (sel_d0_117[2:0] == 2) begin
        next_mux_d0_117 = input_word_d[938];
    end else if (sel_d0_117[2:0] == 3) begin
        next_mux_d0_117 = input_word_d[939];
    end else if (sel_d0_117[2:0] == 4) begin
        next_mux_d0_117 = input_word_d[940];
    end else if (sel_d0_117[2:0] == 5) begin
        next_mux_d0_117 = input_word_d[941];
    end else if (sel_d0_117[2:0] == 6) begin
        next_mux_d0_117 = input_word_d[942];
    end else begin
        next_mux_d0_117 = input_word_d[943];
    end

    if (sel_d0_118[2:0] == 0) begin
        next_mux_d0_118 = input_word_d[944];
    end else if (sel_d0_118[2:0] == 1) begin
        next_mux_d0_118 = input_word_d[945];
    end else if (sel_d0_118[2:0] == 2) begin
        next_mux_d0_118 = input_word_d[946];
    end else if (sel_d0_118[2:0] == 3) begin
        next_mux_d0_118 = input_word_d[947];
    end else if (sel_d0_118[2:0] == 4) begin
        next_mux_d0_118 = input_word_d[948];
    end else if (sel_d0_118[2:0] == 5) begin
        next_mux_d0_118 = input_word_d[949];
    end else if (sel_d0_118[2:0] == 6) begin
        next_mux_d0_118 = input_word_d[950];
    end else begin
        next_mux_d0_118 = input_word_d[951];
    end

    if (sel_d0_119[2:0] == 0) begin
        next_mux_d0_119 = input_word_d[952];
    end else if (sel_d0_119[2:0] == 1) begin
        next_mux_d0_119 = input_word_d[953];
    end else if (sel_d0_119[2:0] == 2) begin
        next_mux_d0_119 = input_word_d[954];
    end else if (sel_d0_119[2:0] == 3) begin
        next_mux_d0_119 = input_word_d[955];
    end else if (sel_d0_119[2:0] == 4) begin
        next_mux_d0_119 = input_word_d[956];
    end else if (sel_d0_119[2:0] == 5) begin
        next_mux_d0_119 = input_word_d[957];
    end else if (sel_d0_119[2:0] == 6) begin
        next_mux_d0_119 = input_word_d[958];
    end else begin
        next_mux_d0_119 = input_word_d[959];
    end

    if (sel_d0_120[2:0] == 0) begin
        next_mux_d0_120 = input_word_d[960];
    end else if (sel_d0_120[2:0] == 1) begin
        next_mux_d0_120 = input_word_d[961];
    end else if (sel_d0_120[2:0] == 2) begin
        next_mux_d0_120 = input_word_d[962];
    end else if (sel_d0_120[2:0] == 3) begin
        next_mux_d0_120 = input_word_d[963];
    end else if (sel_d0_120[2:0] == 4) begin
        next_mux_d0_120 = input_word_d[964];
    end else if (sel_d0_120[2:0] == 5) begin
        next_mux_d0_120 = input_word_d[965];
    end else if (sel_d0_120[2:0] == 6) begin
        next_mux_d0_120 = input_word_d[966];
    end else begin
        next_mux_d0_120 = input_word_d[967];
    end

    if (sel_d0_121[2:0] == 0) begin
        next_mux_d0_121 = input_word_d[968];
    end else if (sel_d0_121[2:0] == 1) begin
        next_mux_d0_121 = input_word_d[969];
    end else if (sel_d0_121[2:0] == 2) begin
        next_mux_d0_121 = input_word_d[970];
    end else if (sel_d0_121[2:0] == 3) begin
        next_mux_d0_121 = input_word_d[971];
    end else if (sel_d0_121[2:0] == 4) begin
        next_mux_d0_121 = input_word_d[972];
    end else if (sel_d0_121[2:0] == 5) begin
        next_mux_d0_121 = input_word_d[973];
    end else if (sel_d0_121[2:0] == 6) begin
        next_mux_d0_121 = input_word_d[974];
    end else begin
        next_mux_d0_121 = input_word_d[975];
    end

    if (sel_d0_122[2:0] == 0) begin
        next_mux_d0_122 = input_word_d[976];
    end else if (sel_d0_122[2:0] == 1) begin
        next_mux_d0_122 = input_word_d[977];
    end else if (sel_d0_122[2:0] == 2) begin
        next_mux_d0_122 = input_word_d[978];
    end else if (sel_d0_122[2:0] == 3) begin
        next_mux_d0_122 = input_word_d[979];
    end else if (sel_d0_122[2:0] == 4) begin
        next_mux_d0_122 = input_word_d[980];
    end else if (sel_d0_122[2:0] == 5) begin
        next_mux_d0_122 = input_word_d[981];
    end else if (sel_d0_122[2:0] == 6) begin
        next_mux_d0_122 = input_word_d[982];
    end else begin
        next_mux_d0_122 = input_word_d[983];
    end

    if (sel_d0_123[2:0] == 0) begin
        next_mux_d0_123 = input_word_d[984];
    end else if (sel_d0_123[2:0] == 1) begin
        next_mux_d0_123 = input_word_d[985];
    end else if (sel_d0_123[2:0] == 2) begin
        next_mux_d0_123 = input_word_d[986];
    end else if (sel_d0_123[2:0] == 3) begin
        next_mux_d0_123 = input_word_d[987];
    end else if (sel_d0_123[2:0] == 4) begin
        next_mux_d0_123 = input_word_d[988];
    end else if (sel_d0_123[2:0] == 5) begin
        next_mux_d0_123 = input_word_d[989];
    end else if (sel_d0_123[2:0] == 6) begin
        next_mux_d0_123 = input_word_d[990];
    end else begin
        next_mux_d0_123 = input_word_d[991];
    end

    if (sel_d0_124[2:0] == 0) begin
        next_mux_d0_124 = input_word_d[992];
    end else if (sel_d0_124[2:0] == 1) begin
        next_mux_d0_124 = input_word_d[993];
    end else if (sel_d0_124[2:0] == 2) begin
        next_mux_d0_124 = input_word_d[994];
    end else if (sel_d0_124[2:0] == 3) begin
        next_mux_d0_124 = input_word_d[995];
    end else if (sel_d0_124[2:0] == 4) begin
        next_mux_d0_124 = input_word_d[996];
    end else if (sel_d0_124[2:0] == 5) begin
        next_mux_d0_124 = input_word_d[997];
    end else if (sel_d0_124[2:0] == 6) begin
        next_mux_d0_124 = input_word_d[998];
    end else begin
        next_mux_d0_124 = input_word_d[999];
    end

    if (sel_d0_125[2:0] == 0) begin
        next_mux_d0_125 = input_word_d[1000];
    end else if (sel_d0_125[2:0] == 1) begin
        next_mux_d0_125 = input_word_d[1001];
    end else if (sel_d0_125[2:0] == 2) begin
        next_mux_d0_125 = input_word_d[1002];
    end else if (sel_d0_125[2:0] == 3) begin
        next_mux_d0_125 = input_word_d[1003];
    end else if (sel_d0_125[2:0] == 4) begin
        next_mux_d0_125 = input_word_d[1004];
    end else if (sel_d0_125[2:0] == 5) begin
        next_mux_d0_125 = input_word_d[1005];
    end else if (sel_d0_125[2:0] == 6) begin
        next_mux_d0_125 = input_word_d[1006];
    end else begin
        next_mux_d0_125 = input_word_d[1007];
    end

    if (sel_d0_126[2:0] == 0) begin
        next_mux_d0_126 = input_word_d[1008];
    end else if (sel_d0_126[2:0] == 1) begin
        next_mux_d0_126 = input_word_d[1009];
    end else if (sel_d0_126[2:0] == 2) begin
        next_mux_d0_126 = input_word_d[1010];
    end else if (sel_d0_126[2:0] == 3) begin
        next_mux_d0_126 = input_word_d[1011];
    end else if (sel_d0_126[2:0] == 4) begin
        next_mux_d0_126 = input_word_d[1012];
    end else if (sel_d0_126[2:0] == 5) begin
        next_mux_d0_126 = input_word_d[1013];
    end else if (sel_d0_126[2:0] == 6) begin
        next_mux_d0_126 = input_word_d[1014];
    end else begin
        next_mux_d0_126 = input_word_d[1015];
    end

    if (sel_d0_127[2:0] == 0) begin
        next_mux_d0_127 = input_word_d[1016];
    end else if (sel_d0_127[2:0] == 1) begin
        next_mux_d0_127 = input_word_d[1017];
    end else if (sel_d0_127[2:0] == 2) begin
        next_mux_d0_127 = input_word_d[1018];
    end else if (sel_d0_127[2:0] == 3) begin
        next_mux_d0_127 = input_word_d[1019];
    end else if (sel_d0_127[2:0] == 4) begin
        next_mux_d0_127 = input_word_d[1020];
    end else if (sel_d0_127[2:0] == 5) begin
        next_mux_d0_127 = input_word_d[1021];
    end else if (sel_d0_127[2:0] == 6) begin
        next_mux_d0_127 = input_word_d[1022];
    end else begin
        next_mux_d0_127 = input_word_d[1023];
    end

    if (sel_d0_128[2:0] == 0) begin
        next_mux_d0_128 = input_word_d[1024];
    end else if (sel_d0_128[2:0] == 1) begin
        next_mux_d0_128 = input_word_d[1025];
    end else if (sel_d0_128[2:0] == 2) begin
        next_mux_d0_128 = input_word_d[1026];
    end else if (sel_d0_128[2:0] == 3) begin
        next_mux_d0_128 = input_word_d[1027];
    end else if (sel_d0_128[2:0] == 4) begin
        next_mux_d0_128 = input_word_d[1028];
    end else if (sel_d0_128[2:0] == 5) begin
        next_mux_d0_128 = input_word_d[1029];
    end else if (sel_d0_128[2:0] == 6) begin
        next_mux_d0_128 = input_word_d[1030];
    end else begin
        next_mux_d0_128 = input_word_d[1031];
    end

    if (sel_d0_129[2:0] == 0) begin
        next_mux_d0_129 = input_word_d[1032];
    end else if (sel_d0_129[2:0] == 1) begin
        next_mux_d0_129 = input_word_d[1033];
    end else if (sel_d0_129[2:0] == 2) begin
        next_mux_d0_129 = input_word_d[1034];
    end else if (sel_d0_129[2:0] == 3) begin
        next_mux_d0_129 = input_word_d[1035];
    end else if (sel_d0_129[2:0] == 4) begin
        next_mux_d0_129 = input_word_d[1036];
    end else if (sel_d0_129[2:0] == 5) begin
        next_mux_d0_129 = input_word_d[1037];
    end else if (sel_d0_129[2:0] == 6) begin
        next_mux_d0_129 = input_word_d[1038];
    end else begin
        next_mux_d0_129 = input_word_d[1039];
    end

    if (sel_d0_130[2:0] == 0) begin
        next_mux_d0_130 = input_word_d[1040];
    end else if (sel_d0_130[2:0] == 1) begin
        next_mux_d0_130 = input_word_d[1041];
    end else if (sel_d0_130[2:0] == 2) begin
        next_mux_d0_130 = input_word_d[1042];
    end else if (sel_d0_130[2:0] == 3) begin
        next_mux_d0_130 = input_word_d[1043];
    end else if (sel_d0_130[2:0] == 4) begin
        next_mux_d0_130 = input_word_d[1044];
    end else if (sel_d0_130[2:0] == 5) begin
        next_mux_d0_130 = input_word_d[1045];
    end else if (sel_d0_130[2:0] == 6) begin
        next_mux_d0_130 = input_word_d[1046];
    end else begin
        next_mux_d0_130 = input_word_d[1047];
    end

    if (sel_d0_131[2:0] == 0) begin
        next_mux_d0_131 = input_word_d[1048];
    end else if (sel_d0_131[2:0] == 1) begin
        next_mux_d0_131 = input_word_d[1049];
    end else if (sel_d0_131[2:0] == 2) begin
        next_mux_d0_131 = input_word_d[1050];
    end else if (sel_d0_131[2:0] == 3) begin
        next_mux_d0_131 = input_word_d[1051];
    end else if (sel_d0_131[2:0] == 4) begin
        next_mux_d0_131 = input_word_d[1052];
    end else if (sel_d0_131[2:0] == 5) begin
        next_mux_d0_131 = input_word_d[1053];
    end else if (sel_d0_131[2:0] == 6) begin
        next_mux_d0_131 = input_word_d[1054];
    end else begin
        next_mux_d0_131 = input_word_d[1055];
    end

    if (sel_d0_132[2:0] == 0) begin
        next_mux_d0_132 = input_word_d[1056];
    end else if (sel_d0_132[2:0] == 1) begin
        next_mux_d0_132 = input_word_d[1057];
    end else if (sel_d0_132[2:0] == 2) begin
        next_mux_d0_132 = input_word_d[1058];
    end else if (sel_d0_132[2:0] == 3) begin
        next_mux_d0_132 = input_word_d[1059];
    end else if (sel_d0_132[2:0] == 4) begin
        next_mux_d0_132 = input_word_d[1060];
    end else if (sel_d0_132[2:0] == 5) begin
        next_mux_d0_132 = input_word_d[1061];
    end else if (sel_d0_132[2:0] == 6) begin
        next_mux_d0_132 = input_word_d[1062];
    end else begin
        next_mux_d0_132 = input_word_d[1063];
    end

    if (sel_d0_133[2:0] == 0) begin
        next_mux_d0_133 = input_word_d[1064];
    end else if (sel_d0_133[2:0] == 1) begin
        next_mux_d0_133 = input_word_d[1065];
    end else if (sel_d0_133[2:0] == 2) begin
        next_mux_d0_133 = input_word_d[1066];
    end else if (sel_d0_133[2:0] == 3) begin
        next_mux_d0_133 = input_word_d[1067];
    end else if (sel_d0_133[2:0] == 4) begin
        next_mux_d0_133 = input_word_d[1068];
    end else if (sel_d0_133[2:0] == 5) begin
        next_mux_d0_133 = input_word_d[1069];
    end else if (sel_d0_133[2:0] == 6) begin
        next_mux_d0_133 = input_word_d[1070];
    end else begin
        next_mux_d0_133 = input_word_d[1071];
    end

    if (sel_d0_134[2:0] == 0) begin
        next_mux_d0_134 = input_word_d[1072];
    end else if (sel_d0_134[2:0] == 1) begin
        next_mux_d0_134 = input_word_d[1073];
    end else if (sel_d0_134[2:0] == 2) begin
        next_mux_d0_134 = input_word_d[1074];
    end else if (sel_d0_134[2:0] == 3) begin
        next_mux_d0_134 = input_word_d[1075];
    end else if (sel_d0_134[2:0] == 4) begin
        next_mux_d0_134 = input_word_d[1076];
    end else if (sel_d0_134[2:0] == 5) begin
        next_mux_d0_134 = input_word_d[1077];
    end else if (sel_d0_134[2:0] == 6) begin
        next_mux_d0_134 = input_word_d[1078];
    end else begin
        next_mux_d0_134 = input_word_d[1079];
    end

    if (sel_d0_135[2:0] == 0) begin
        next_mux_d0_135 = input_word_d[1080];
    end else if (sel_d0_135[2:0] == 1) begin
        next_mux_d0_135 = input_word_d[1081];
    end else if (sel_d0_135[2:0] == 2) begin
        next_mux_d0_135 = input_word_d[1082];
    end else if (sel_d0_135[2:0] == 3) begin
        next_mux_d0_135 = input_word_d[1083];
    end else if (sel_d0_135[2:0] == 4) begin
        next_mux_d0_135 = input_word_d[1084];
    end else if (sel_d0_135[2:0] == 5) begin
        next_mux_d0_135 = input_word_d[1085];
    end else if (sel_d0_135[2:0] == 6) begin
        next_mux_d0_135 = input_word_d[1086];
    end else begin
        next_mux_d0_135 = input_word_d[1087];
    end

    if (sel_d0_136[2:0] == 0) begin
        next_mux_d0_136 = input_word_d[1088];
    end else if (sel_d0_136[2:0] == 1) begin
        next_mux_d0_136 = input_word_d[1089];
    end else if (sel_d0_136[2:0] == 2) begin
        next_mux_d0_136 = input_word_d[1090];
    end else if (sel_d0_136[2:0] == 3) begin
        next_mux_d0_136 = input_word_d[1091];
    end else if (sel_d0_136[2:0] == 4) begin
        next_mux_d0_136 = input_word_d[1092];
    end else if (sel_d0_136[2:0] == 5) begin
        next_mux_d0_136 = input_word_d[1093];
    end else if (sel_d0_136[2:0] == 6) begin
        next_mux_d0_136 = input_word_d[1094];
    end else begin
        next_mux_d0_136 = input_word_d[1095];
    end

    if (sel_d0_137[2:0] == 0) begin
        next_mux_d0_137 = input_word_d[1096];
    end else if (sel_d0_137[2:0] == 1) begin
        next_mux_d0_137 = input_word_d[1097];
    end else if (sel_d0_137[2:0] == 2) begin
        next_mux_d0_137 = input_word_d[1098];
    end else if (sel_d0_137[2:0] == 3) begin
        next_mux_d0_137 = input_word_d[1099];
    end else if (sel_d0_137[2:0] == 4) begin
        next_mux_d0_137 = input_word_d[1100];
    end else if (sel_d0_137[2:0] == 5) begin
        next_mux_d0_137 = input_word_d[1101];
    end else if (sel_d0_137[2:0] == 6) begin
        next_mux_d0_137 = input_word_d[1102];
    end else begin
        next_mux_d0_137 = input_word_d[1103];
    end

    if (sel_d0_138[2:0] == 0) begin
        next_mux_d0_138 = input_word_d[1104];
    end else if (sel_d0_138[2:0] == 1) begin
        next_mux_d0_138 = input_word_d[1105];
    end else if (sel_d0_138[2:0] == 2) begin
        next_mux_d0_138 = input_word_d[1106];
    end else if (sel_d0_138[2:0] == 3) begin
        next_mux_d0_138 = input_word_d[1107];
    end else if (sel_d0_138[2:0] == 4) begin
        next_mux_d0_138 = input_word_d[1108];
    end else if (sel_d0_138[2:0] == 5) begin
        next_mux_d0_138 = input_word_d[1109];
    end else if (sel_d0_138[2:0] == 6) begin
        next_mux_d0_138 = input_word_d[1110];
    end else begin
        next_mux_d0_138 = input_word_d[1111];
    end

    if (sel_d0_139[2:0] == 0) begin
        next_mux_d0_139 = input_word_d[1112];
    end else if (sel_d0_139[2:0] == 1) begin
        next_mux_d0_139 = input_word_d[1113];
    end else if (sel_d0_139[2:0] == 2) begin
        next_mux_d0_139 = input_word_d[1114];
    end else if (sel_d0_139[2:0] == 3) begin
        next_mux_d0_139 = input_word_d[1115];
    end else if (sel_d0_139[2:0] == 4) begin
        next_mux_d0_139 = input_word_d[1116];
    end else if (sel_d0_139[2:0] == 5) begin
        next_mux_d0_139 = input_word_d[1117];
    end else if (sel_d0_139[2:0] == 6) begin
        next_mux_d0_139 = input_word_d[1118];
    end else begin
        next_mux_d0_139 = input_word_d[1119];
    end

    if (sel_d0_140[2:0] == 0) begin
        next_mux_d0_140 = input_word_d[1120];
    end else if (sel_d0_140[2:0] == 1) begin
        next_mux_d0_140 = input_word_d[1121];
    end else if (sel_d0_140[2:0] == 2) begin
        next_mux_d0_140 = input_word_d[1122];
    end else if (sel_d0_140[2:0] == 3) begin
        next_mux_d0_140 = input_word_d[1123];
    end else if (sel_d0_140[2:0] == 4) begin
        next_mux_d0_140 = input_word_d[1124];
    end else if (sel_d0_140[2:0] == 5) begin
        next_mux_d0_140 = input_word_d[1125];
    end else if (sel_d0_140[2:0] == 6) begin
        next_mux_d0_140 = input_word_d[1126];
    end else begin
        next_mux_d0_140 = input_word_d[1127];
    end

    if (sel_d0_141[2:0] == 0) begin
        next_mux_d0_141 = input_word_d[1128];
    end else if (sel_d0_141[2:0] == 1) begin
        next_mux_d0_141 = input_word_d[1129];
    end else if (sel_d0_141[2:0] == 2) begin
        next_mux_d0_141 = input_word_d[1130];
    end else if (sel_d0_141[2:0] == 3) begin
        next_mux_d0_141 = input_word_d[1131];
    end else if (sel_d0_141[2:0] == 4) begin
        next_mux_d0_141 = input_word_d[1132];
    end else if (sel_d0_141[2:0] == 5) begin
        next_mux_d0_141 = input_word_d[1133];
    end else if (sel_d0_141[2:0] == 6) begin
        next_mux_d0_141 = input_word_d[1134];
    end else begin
        next_mux_d0_141 = input_word_d[1135];
    end

    if (sel_d0_142[2:0] == 0) begin
        next_mux_d0_142 = input_word_d[1136];
    end else if (sel_d0_142[2:0] == 1) begin
        next_mux_d0_142 = input_word_d[1137];
    end else if (sel_d0_142[2:0] == 2) begin
        next_mux_d0_142 = input_word_d[1138];
    end else if (sel_d0_142[2:0] == 3) begin
        next_mux_d0_142 = input_word_d[1139];
    end else if (sel_d0_142[2:0] == 4) begin
        next_mux_d0_142 = input_word_d[1140];
    end else if (sel_d0_142[2:0] == 5) begin
        next_mux_d0_142 = input_word_d[1141];
    end else if (sel_d0_142[2:0] == 6) begin
        next_mux_d0_142 = input_word_d[1142];
    end else begin
        next_mux_d0_142 = input_word_d[1143];
    end

    if (sel_d0_143[2:0] == 0) begin
        next_mux_d0_143 = input_word_d[1144];
    end else if (sel_d0_143[2:0] == 1) begin
        next_mux_d0_143 = input_word_d[1145];
    end else if (sel_d0_143[2:0] == 2) begin
        next_mux_d0_143 = input_word_d[1146];
    end else if (sel_d0_143[2:0] == 3) begin
        next_mux_d0_143 = input_word_d[1147];
    end else if (sel_d0_143[2:0] == 4) begin
        next_mux_d0_143 = input_word_d[1148];
    end else if (sel_d0_143[2:0] == 5) begin
        next_mux_d0_143 = input_word_d[1149];
    end else if (sel_d0_143[2:0] == 6) begin
        next_mux_d0_143 = input_word_d[1150];
    end else begin
        next_mux_d0_143 = input_word_d[1151];
    end

    if (sel_d0_144[2:0] == 0) begin
        next_mux_d0_144 = input_word_d[1152];
    end else if (sel_d0_144[2:0] == 1) begin
        next_mux_d0_144 = input_word_d[1153];
    end else if (sel_d0_144[2:0] == 2) begin
        next_mux_d0_144 = input_word_d[1154];
    end else if (sel_d0_144[2:0] == 3) begin
        next_mux_d0_144 = input_word_d[1155];
    end else if (sel_d0_144[2:0] == 4) begin
        next_mux_d0_144 = input_word_d[1156];
    end else if (sel_d0_144[2:0] == 5) begin
        next_mux_d0_144 = input_word_d[1157];
    end else if (sel_d0_144[2:0] == 6) begin
        next_mux_d0_144 = input_word_d[1158];
    end else begin
        next_mux_d0_144 = input_word_d[1159];
    end

    if (sel_d0_145[2:0] == 0) begin
        next_mux_d0_145 = input_word_d[1160];
    end else if (sel_d0_145[2:0] == 1) begin
        next_mux_d0_145 = input_word_d[1161];
    end else if (sel_d0_145[2:0] == 2) begin
        next_mux_d0_145 = input_word_d[1162];
    end else if (sel_d0_145[2:0] == 3) begin
        next_mux_d0_145 = input_word_d[1163];
    end else if (sel_d0_145[2:0] == 4) begin
        next_mux_d0_145 = input_word_d[1164];
    end else if (sel_d0_145[2:0] == 5) begin
        next_mux_d0_145 = input_word_d[1165];
    end else if (sel_d0_145[2:0] == 6) begin
        next_mux_d0_145 = input_word_d[1166];
    end else begin
        next_mux_d0_145 = input_word_d[1167];
    end

    if (sel_d0_146[2:0] == 0) begin
        next_mux_d0_146 = input_word_d[1168];
    end else if (sel_d0_146[2:0] == 1) begin
        next_mux_d0_146 = input_word_d[1169];
    end else if (sel_d0_146[2:0] == 2) begin
        next_mux_d0_146 = input_word_d[1170];
    end else if (sel_d0_146[2:0] == 3) begin
        next_mux_d0_146 = input_word_d[1171];
    end else if (sel_d0_146[2:0] == 4) begin
        next_mux_d0_146 = input_word_d[1172];
    end else if (sel_d0_146[2:0] == 5) begin
        next_mux_d0_146 = input_word_d[1173];
    end else if (sel_d0_146[2:0] == 6) begin
        next_mux_d0_146 = input_word_d[1174];
    end else begin
        next_mux_d0_146 = input_word_d[1175];
    end

    if (sel_d0_147[2:0] == 0) begin
        next_mux_d0_147 = input_word_d[1176];
    end else if (sel_d0_147[2:0] == 1) begin
        next_mux_d0_147 = input_word_d[1177];
    end else if (sel_d0_147[2:0] == 2) begin
        next_mux_d0_147 = input_word_d[1178];
    end else if (sel_d0_147[2:0] == 3) begin
        next_mux_d0_147 = input_word_d[1179];
    end else if (sel_d0_147[2:0] == 4) begin
        next_mux_d0_147 = input_word_d[1180];
    end else if (sel_d0_147[2:0] == 5) begin
        next_mux_d0_147 = input_word_d[1181];
    end else if (sel_d0_147[2:0] == 6) begin
        next_mux_d0_147 = input_word_d[1182];
    end else begin
        next_mux_d0_147 = input_word_d[1183];
    end

    if (sel_d0_148[2:0] == 0) begin
        next_mux_d0_148 = input_word_d[1184];
    end else if (sel_d0_148[2:0] == 1) begin
        next_mux_d0_148 = input_word_d[1185];
    end else if (sel_d0_148[2:0] == 2) begin
        next_mux_d0_148 = input_word_d[1186];
    end else if (sel_d0_148[2:0] == 3) begin
        next_mux_d0_148 = input_word_d[1187];
    end else if (sel_d0_148[2:0] == 4) begin
        next_mux_d0_148 = input_word_d[1188];
    end else if (sel_d0_148[2:0] == 5) begin
        next_mux_d0_148 = input_word_d[1189];
    end else if (sel_d0_148[2:0] == 6) begin
        next_mux_d0_148 = input_word_d[1190];
    end else begin
        next_mux_d0_148 = input_word_d[1191];
    end

    if (sel_d0_149[2:0] == 0) begin
        next_mux_d0_149 = input_word_d[1192];
    end else if (sel_d0_149[2:0] == 1) begin
        next_mux_d0_149 = input_word_d[1193];
    end else if (sel_d0_149[2:0] == 2) begin
        next_mux_d0_149 = input_word_d[1194];
    end else if (sel_d0_149[2:0] == 3) begin
        next_mux_d0_149 = input_word_d[1195];
    end else if (sel_d0_149[2:0] == 4) begin
        next_mux_d0_149 = input_word_d[1196];
    end else if (sel_d0_149[2:0] == 5) begin
        next_mux_d0_149 = input_word_d[1197];
    end else if (sel_d0_149[2:0] == 6) begin
        next_mux_d0_149 = input_word_d[1198];
    end else begin
        next_mux_d0_149 = input_word_d[1199];
    end

    if (sel_d0_150[2:0] == 0) begin
        next_mux_d0_150 = input_word_d[1200];
    end else if (sel_d0_150[2:0] == 1) begin
        next_mux_d0_150 = input_word_d[1201];
    end else if (sel_d0_150[2:0] == 2) begin
        next_mux_d0_150 = input_word_d[1202];
    end else if (sel_d0_150[2:0] == 3) begin
        next_mux_d0_150 = input_word_d[1203];
    end else if (sel_d0_150[2:0] == 4) begin
        next_mux_d0_150 = input_word_d[1204];
    end else if (sel_d0_150[2:0] == 5) begin
        next_mux_d0_150 = input_word_d[1205];
    end else if (sel_d0_150[2:0] == 6) begin
        next_mux_d0_150 = input_word_d[1206];
    end else begin
        next_mux_d0_150 = input_word_d[1207];
    end

    if (sel_d0_151[2:0] == 0) begin
        next_mux_d0_151 = input_word_d[1208];
    end else if (sel_d0_151[2:0] == 1) begin
        next_mux_d0_151 = input_word_d[1209];
    end else if (sel_d0_151[2:0] == 2) begin
        next_mux_d0_151 = input_word_d[1210];
    end else if (sel_d0_151[2:0] == 3) begin
        next_mux_d0_151 = input_word_d[1211];
    end else if (sel_d0_151[2:0] == 4) begin
        next_mux_d0_151 = input_word_d[1212];
    end else if (sel_d0_151[2:0] == 5) begin
        next_mux_d0_151 = input_word_d[1213];
    end else if (sel_d0_151[2:0] == 6) begin
        next_mux_d0_151 = input_word_d[1214];
    end else begin
        next_mux_d0_151 = input_word_d[1215];
    end

    if (sel_d0_152[2:0] == 0) begin
        next_mux_d0_152 = input_word_d[1216];
    end else if (sel_d0_152[2:0] == 1) begin
        next_mux_d0_152 = input_word_d[1217];
    end else if (sel_d0_152[2:0] == 2) begin
        next_mux_d0_152 = input_word_d[1218];
    end else if (sel_d0_152[2:0] == 3) begin
        next_mux_d0_152 = input_word_d[1219];
    end else if (sel_d0_152[2:0] == 4) begin
        next_mux_d0_152 = input_word_d[1220];
    end else if (sel_d0_152[2:0] == 5) begin
        next_mux_d0_152 = input_word_d[1221];
    end else if (sel_d0_152[2:0] == 6) begin
        next_mux_d0_152 = input_word_d[1222];
    end else begin
        next_mux_d0_152 = input_word_d[1223];
    end

    if (sel_d0_153[2:0] == 0) begin
        next_mux_d0_153 = input_word_d[1224];
    end else if (sel_d0_153[2:0] == 1) begin
        next_mux_d0_153 = input_word_d[1225];
    end else if (sel_d0_153[2:0] == 2) begin
        next_mux_d0_153 = input_word_d[1226];
    end else if (sel_d0_153[2:0] == 3) begin
        next_mux_d0_153 = input_word_d[1227];
    end else if (sel_d0_153[2:0] == 4) begin
        next_mux_d0_153 = input_word_d[1228];
    end else if (sel_d0_153[2:0] == 5) begin
        next_mux_d0_153 = input_word_d[1229];
    end else if (sel_d0_153[2:0] == 6) begin
        next_mux_d0_153 = input_word_d[1230];
    end else begin
        next_mux_d0_153 = input_word_d[1231];
    end

    if (sel_d0_154[2:0] == 0) begin
        next_mux_d0_154 = input_word_d[1232];
    end else if (sel_d0_154[2:0] == 1) begin
        next_mux_d0_154 = input_word_d[1233];
    end else if (sel_d0_154[2:0] == 2) begin
        next_mux_d0_154 = input_word_d[1234];
    end else if (sel_d0_154[2:0] == 3) begin
        next_mux_d0_154 = input_word_d[1235];
    end else if (sel_d0_154[2:0] == 4) begin
        next_mux_d0_154 = input_word_d[1236];
    end else if (sel_d0_154[2:0] == 5) begin
        next_mux_d0_154 = input_word_d[1237];
    end else if (sel_d0_154[2:0] == 6) begin
        next_mux_d0_154 = input_word_d[1238];
    end else begin
        next_mux_d0_154 = input_word_d[1239];
    end

    if (sel_d0_155[2:0] == 0) begin
        next_mux_d0_155 = input_word_d[1240];
    end else if (sel_d0_155[2:0] == 1) begin
        next_mux_d0_155 = input_word_d[1241];
    end else if (sel_d0_155[2:0] == 2) begin
        next_mux_d0_155 = input_word_d[1242];
    end else if (sel_d0_155[2:0] == 3) begin
        next_mux_d0_155 = input_word_d[1243];
    end else if (sel_d0_155[2:0] == 4) begin
        next_mux_d0_155 = input_word_d[1244];
    end else if (sel_d0_155[2:0] == 5) begin
        next_mux_d0_155 = input_word_d[1245];
    end else if (sel_d0_155[2:0] == 6) begin
        next_mux_d0_155 = input_word_d[1246];
    end else begin
        next_mux_d0_155 = input_word_d[1247];
    end

    if (sel_d0_156[2:0] == 0) begin
        next_mux_d0_156 = input_word_d[1248];
    end else if (sel_d0_156[2:0] == 1) begin
        next_mux_d0_156 = input_word_d[1249];
    end else if (sel_d0_156[2:0] == 2) begin
        next_mux_d0_156 = input_word_d[1250];
    end else if (sel_d0_156[2:0] == 3) begin
        next_mux_d0_156 = input_word_d[1251];
    end else if (sel_d0_156[2:0] == 4) begin
        next_mux_d0_156 = input_word_d[1252];
    end else if (sel_d0_156[2:0] == 5) begin
        next_mux_d0_156 = input_word_d[1253];
    end else if (sel_d0_156[2:0] == 6) begin
        next_mux_d0_156 = input_word_d[1254];
    end else begin
        next_mux_d0_156 = input_word_d[1255];
    end

    if (sel_d0_157[2:0] == 0) begin
        next_mux_d0_157 = input_word_d[1256];
    end else if (sel_d0_157[2:0] == 1) begin
        next_mux_d0_157 = input_word_d[1257];
    end else if (sel_d0_157[2:0] == 2) begin
        next_mux_d0_157 = input_word_d[1258];
    end else if (sel_d0_157[2:0] == 3) begin
        next_mux_d0_157 = input_word_d[1259];
    end else if (sel_d0_157[2:0] == 4) begin
        next_mux_d0_157 = input_word_d[1260];
    end else if (sel_d0_157[2:0] == 5) begin
        next_mux_d0_157 = input_word_d[1261];
    end else if (sel_d0_157[2:0] == 6) begin
        next_mux_d0_157 = input_word_d[1262];
    end else begin
        next_mux_d0_157 = input_word_d[1263];
    end

    if (sel_d0_158[2:0] == 0) begin
        next_mux_d0_158 = input_word_d[1264];
    end else if (sel_d0_158[2:0] == 1) begin
        next_mux_d0_158 = input_word_d[1265];
    end else if (sel_d0_158[2:0] == 2) begin
        next_mux_d0_158 = input_word_d[1266];
    end else if (sel_d0_158[2:0] == 3) begin
        next_mux_d0_158 = input_word_d[1267];
    end else if (sel_d0_158[2:0] == 4) begin
        next_mux_d0_158 = input_word_d[1268];
    end else if (sel_d0_158[2:0] == 5) begin
        next_mux_d0_158 = input_word_d[1269];
    end else if (sel_d0_158[2:0] == 6) begin
        next_mux_d0_158 = input_word_d[1270];
    end else begin
        next_mux_d0_158 = input_word_d[1271];
    end

    if (sel_d0_159[2:0] == 0) begin
        next_mux_d0_159 = input_word_d[1272];
    end else if (sel_d0_159[2:0] == 1) begin
        next_mux_d0_159 = input_word_d[1273];
    end else if (sel_d0_159[2:0] == 2) begin
        next_mux_d0_159 = input_word_d[1274];
    end else if (sel_d0_159[2:0] == 3) begin
        next_mux_d0_159 = input_word_d[1275];
    end else if (sel_d0_159[2:0] == 4) begin
        next_mux_d0_159 = input_word_d[1276];
    end else if (sel_d0_159[2:0] == 5) begin
        next_mux_d0_159 = input_word_d[1277];
    end else if (sel_d0_159[2:0] == 6) begin
        next_mux_d0_159 = input_word_d[1278];
    end else begin
        next_mux_d0_159 = input_word_d[1279];
    end

    if (sel_d0_160[2:0] == 0) begin
        next_mux_d0_160 = input_word_d[1280];
    end else if (sel_d0_160[2:0] == 1) begin
        next_mux_d0_160 = input_word_d[1281];
    end else if (sel_d0_160[2:0] == 2) begin
        next_mux_d0_160 = input_word_d[1282];
    end else if (sel_d0_160[2:0] == 3) begin
        next_mux_d0_160 = input_word_d[1283];
    end else if (sel_d0_160[2:0] == 4) begin
        next_mux_d0_160 = input_word_d[1284];
    end else if (sel_d0_160[2:0] == 5) begin
        next_mux_d0_160 = input_word_d[1285];
    end else if (sel_d0_160[2:0] == 6) begin
        next_mux_d0_160 = input_word_d[1286];
    end else begin
        next_mux_d0_160 = input_word_d[1287];
    end

    if (sel_d0_161[2:0] == 0) begin
        next_mux_d0_161 = input_word_d[1288];
    end else if (sel_d0_161[2:0] == 1) begin
        next_mux_d0_161 = input_word_d[1289];
    end else if (sel_d0_161[2:0] == 2) begin
        next_mux_d0_161 = input_word_d[1290];
    end else if (sel_d0_161[2:0] == 3) begin
        next_mux_d0_161 = input_word_d[1291];
    end else if (sel_d0_161[2:0] == 4) begin
        next_mux_d0_161 = input_word_d[1292];
    end else if (sel_d0_161[2:0] == 5) begin
        next_mux_d0_161 = input_word_d[1293];
    end else if (sel_d0_161[2:0] == 6) begin
        next_mux_d0_161 = input_word_d[1294];
    end else begin
        next_mux_d0_161 = input_word_d[1295];
    end

    if (sel_d0_162[2:0] == 0) begin
        next_mux_d0_162 = input_word_d[1296];
    end else if (sel_d0_162[2:0] == 1) begin
        next_mux_d0_162 = input_word_d[1297];
    end else if (sel_d0_162[2:0] == 2) begin
        next_mux_d0_162 = input_word_d[1298];
    end else if (sel_d0_162[2:0] == 3) begin
        next_mux_d0_162 = input_word_d[1299];
    end else if (sel_d0_162[2:0] == 4) begin
        next_mux_d0_162 = input_word_d[1300];
    end else if (sel_d0_162[2:0] == 5) begin
        next_mux_d0_162 = input_word_d[1301];
    end else if (sel_d0_162[2:0] == 6) begin
        next_mux_d0_162 = input_word_d[1302];
    end else begin
        next_mux_d0_162 = input_word_d[1303];
    end

    if (sel_d0_163[2:0] == 0) begin
        next_mux_d0_163 = input_word_d[1304];
    end else if (sel_d0_163[2:0] == 1) begin
        next_mux_d0_163 = input_word_d[1305];
    end else if (sel_d0_163[2:0] == 2) begin
        next_mux_d0_163 = input_word_d[1306];
    end else if (sel_d0_163[2:0] == 3) begin
        next_mux_d0_163 = input_word_d[1307];
    end else if (sel_d0_163[2:0] == 4) begin
        next_mux_d0_163 = input_word_d[1308];
    end else if (sel_d0_163[2:0] == 5) begin
        next_mux_d0_163 = input_word_d[1309];
    end else if (sel_d0_163[2:0] == 6) begin
        next_mux_d0_163 = input_word_d[1310];
    end else begin
        next_mux_d0_163 = input_word_d[1311];
    end

    if (sel_d0_164[2:0] == 0) begin
        next_mux_d0_164 = input_word_d[1312];
    end else if (sel_d0_164[2:0] == 1) begin
        next_mux_d0_164 = input_word_d[1313];
    end else if (sel_d0_164[2:0] == 2) begin
        next_mux_d0_164 = input_word_d[1314];
    end else if (sel_d0_164[2:0] == 3) begin
        next_mux_d0_164 = input_word_d[1315];
    end else if (sel_d0_164[2:0] == 4) begin
        next_mux_d0_164 = input_word_d[1316];
    end else if (sel_d0_164[2:0] == 5) begin
        next_mux_d0_164 = input_word_d[1317];
    end else if (sel_d0_164[2:0] == 6) begin
        next_mux_d0_164 = input_word_d[1318];
    end else begin
        next_mux_d0_164 = input_word_d[1319];
    end

    if (sel_d0_165[2:0] == 0) begin
        next_mux_d0_165 = input_word_d[1320];
    end else if (sel_d0_165[2:0] == 1) begin
        next_mux_d0_165 = input_word_d[1321];
    end else if (sel_d0_165[2:0] == 2) begin
        next_mux_d0_165 = input_word_d[1322];
    end else if (sel_d0_165[2:0] == 3) begin
        next_mux_d0_165 = input_word_d[1323];
    end else if (sel_d0_165[2:0] == 4) begin
        next_mux_d0_165 = input_word_d[1324];
    end else if (sel_d0_165[2:0] == 5) begin
        next_mux_d0_165 = input_word_d[1325];
    end else if (sel_d0_165[2:0] == 6) begin
        next_mux_d0_165 = input_word_d[1326];
    end else begin
        next_mux_d0_165 = input_word_d[1327];
    end

    if (sel_d0_166[2:0] == 0) begin
        next_mux_d0_166 = input_word_d[1328];
    end else if (sel_d0_166[2:0] == 1) begin
        next_mux_d0_166 = input_word_d[1329];
    end else if (sel_d0_166[2:0] == 2) begin
        next_mux_d0_166 = input_word_d[1330];
    end else if (sel_d0_166[2:0] == 3) begin
        next_mux_d0_166 = input_word_d[1331];
    end else if (sel_d0_166[2:0] == 4) begin
        next_mux_d0_166 = input_word_d[1332];
    end else if (sel_d0_166[2:0] == 5) begin
        next_mux_d0_166 = input_word_d[1333];
    end else if (sel_d0_166[2:0] == 6) begin
        next_mux_d0_166 = input_word_d[1334];
    end else begin
        next_mux_d0_166 = input_word_d[1335];
    end

    if (sel_d0_167[2:0] == 0) begin
        next_mux_d0_167 = input_word_d[1336];
    end else if (sel_d0_167[2:0] == 1) begin
        next_mux_d0_167 = input_word_d[1337];
    end else if (sel_d0_167[2:0] == 2) begin
        next_mux_d0_167 = input_word_d[1338];
    end else if (sel_d0_167[2:0] == 3) begin
        next_mux_d0_167 = input_word_d[1339];
    end else if (sel_d0_167[2:0] == 4) begin
        next_mux_d0_167 = input_word_d[1340];
    end else if (sel_d0_167[2:0] == 5) begin
        next_mux_d0_167 = input_word_d[1341];
    end else if (sel_d0_167[2:0] == 6) begin
        next_mux_d0_167 = input_word_d[1342];
    end else begin
        next_mux_d0_167 = input_word_d[1343];
    end

    if (sel_d0_168[2:0] == 0) begin
        next_mux_d0_168 = input_word_d[1344];
    end else if (sel_d0_168[2:0] == 1) begin
        next_mux_d0_168 = input_word_d[1345];
    end else if (sel_d0_168[2:0] == 2) begin
        next_mux_d0_168 = input_word_d[1346];
    end else if (sel_d0_168[2:0] == 3) begin
        next_mux_d0_168 = input_word_d[1347];
    end else if (sel_d0_168[2:0] == 4) begin
        next_mux_d0_168 = input_word_d[1348];
    end else if (sel_d0_168[2:0] == 5) begin
        next_mux_d0_168 = input_word_d[1349];
    end else if (sel_d0_168[2:0] == 6) begin
        next_mux_d0_168 = input_word_d[1350];
    end else begin
        next_mux_d0_168 = input_word_d[1351];
    end

    if (sel_d0_169[2:0] == 0) begin
        next_mux_d0_169 = input_word_d[1352];
    end else if (sel_d0_169[2:0] == 1) begin
        next_mux_d0_169 = input_word_d[1353];
    end else if (sel_d0_169[2:0] == 2) begin
        next_mux_d0_169 = input_word_d[1354];
    end else if (sel_d0_169[2:0] == 3) begin
        next_mux_d0_169 = input_word_d[1355];
    end else if (sel_d0_169[2:0] == 4) begin
        next_mux_d0_169 = input_word_d[1356];
    end else if (sel_d0_169[2:0] == 5) begin
        next_mux_d0_169 = input_word_d[1357];
    end else if (sel_d0_169[2:0] == 6) begin
        next_mux_d0_169 = input_word_d[1358];
    end else begin
        next_mux_d0_169 = input_word_d[1359];
    end

    if (sel_d0_170[2:0] == 0) begin
        next_mux_d0_170 = input_word_d[1360];
    end else if (sel_d0_170[2:0] == 1) begin
        next_mux_d0_170 = input_word_d[1361];
    end else if (sel_d0_170[2:0] == 2) begin
        next_mux_d0_170 = input_word_d[1362];
    end else if (sel_d0_170[2:0] == 3) begin
        next_mux_d0_170 = input_word_d[1363];
    end else if (sel_d0_170[2:0] == 4) begin
        next_mux_d0_170 = input_word_d[1364];
    end else if (sel_d0_170[2:0] == 5) begin
        next_mux_d0_170 = input_word_d[1365];
    end else if (sel_d0_170[2:0] == 6) begin
        next_mux_d0_170 = input_word_d[1366];
    end else begin
        next_mux_d0_170 = input_word_d[1367];
    end

    if (sel_d0_171[2:0] == 0) begin
        next_mux_d0_171 = input_word_d[1368];
    end else if (sel_d0_171[2:0] == 1) begin
        next_mux_d0_171 = input_word_d[1369];
    end else if (sel_d0_171[2:0] == 2) begin
        next_mux_d0_171 = input_word_d[1370];
    end else if (sel_d0_171[2:0] == 3) begin
        next_mux_d0_171 = input_word_d[1371];
    end else if (sel_d0_171[2:0] == 4) begin
        next_mux_d0_171 = input_word_d[1372];
    end else if (sel_d0_171[2:0] == 5) begin
        next_mux_d0_171 = input_word_d[1373];
    end else if (sel_d0_171[2:0] == 6) begin
        next_mux_d0_171 = input_word_d[1374];
    end else begin
        next_mux_d0_171 = input_word_d[1375];
    end

    if (sel_d0_172[2:0] == 0) begin
        next_mux_d0_172 = input_word_d[1376];
    end else if (sel_d0_172[2:0] == 1) begin
        next_mux_d0_172 = input_word_d[1377];
    end else if (sel_d0_172[2:0] == 2) begin
        next_mux_d0_172 = input_word_d[1378];
    end else if (sel_d0_172[2:0] == 3) begin
        next_mux_d0_172 = input_word_d[1379];
    end else if (sel_d0_172[2:0] == 4) begin
        next_mux_d0_172 = input_word_d[1380];
    end else if (sel_d0_172[2:0] == 5) begin
        next_mux_d0_172 = input_word_d[1381];
    end else if (sel_d0_172[2:0] == 6) begin
        next_mux_d0_172 = input_word_d[1382];
    end else begin
        next_mux_d0_172 = input_word_d[1383];
    end

    if (sel_d0_173[2:0] == 0) begin
        next_mux_d0_173 = input_word_d[1384];
    end else if (sel_d0_173[2:0] == 1) begin
        next_mux_d0_173 = input_word_d[1385];
    end else if (sel_d0_173[2:0] == 2) begin
        next_mux_d0_173 = input_word_d[1386];
    end else if (sel_d0_173[2:0] == 3) begin
        next_mux_d0_173 = input_word_d[1387];
    end else if (sel_d0_173[2:0] == 4) begin
        next_mux_d0_173 = input_word_d[1388];
    end else if (sel_d0_173[2:0] == 5) begin
        next_mux_d0_173 = input_word_d[1389];
    end else if (sel_d0_173[2:0] == 6) begin
        next_mux_d0_173 = input_word_d[1390];
    end else begin
        next_mux_d0_173 = input_word_d[1391];
    end

    if (sel_d0_174[2:0] == 0) begin
        next_mux_d0_174 = input_word_d[1392];
    end else if (sel_d0_174[2:0] == 1) begin
        next_mux_d0_174 = input_word_d[1393];
    end else if (sel_d0_174[2:0] == 2) begin
        next_mux_d0_174 = input_word_d[1394];
    end else if (sel_d0_174[2:0] == 3) begin
        next_mux_d0_174 = input_word_d[1395];
    end else if (sel_d0_174[2:0] == 4) begin
        next_mux_d0_174 = input_word_d[1396];
    end else if (sel_d0_174[2:0] == 5) begin
        next_mux_d0_174 = input_word_d[1397];
    end else if (sel_d0_174[2:0] == 6) begin
        next_mux_d0_174 = input_word_d[1398];
    end else begin
        next_mux_d0_174 = input_word_d[1399];
    end

    if (sel_d0_175[2:0] == 0) begin
        next_mux_d0_175 = input_word_d[1400];
    end else if (sel_d0_175[2:0] == 1) begin
        next_mux_d0_175 = input_word_d[1401];
    end else if (sel_d0_175[2:0] == 2) begin
        next_mux_d0_175 = input_word_d[1402];
    end else if (sel_d0_175[2:0] == 3) begin
        next_mux_d0_175 = input_word_d[1403];
    end else if (sel_d0_175[2:0] == 4) begin
        next_mux_d0_175 = input_word_d[1404];
    end else if (sel_d0_175[2:0] == 5) begin
        next_mux_d0_175 = input_word_d[1405];
    end else if (sel_d0_175[2:0] == 6) begin
        next_mux_d0_175 = input_word_d[1406];
    end else begin
        next_mux_d0_175 = input_word_d[1407];
    end

    if (sel_d0_176[2:0] == 0) begin
        next_mux_d0_176 = input_word_d[1408];
    end else if (sel_d0_176[2:0] == 1) begin
        next_mux_d0_176 = input_word_d[1409];
    end else if (sel_d0_176[2:0] == 2) begin
        next_mux_d0_176 = input_word_d[1410];
    end else if (sel_d0_176[2:0] == 3) begin
        next_mux_d0_176 = input_word_d[1411];
    end else if (sel_d0_176[2:0] == 4) begin
        next_mux_d0_176 = input_word_d[1412];
    end else if (sel_d0_176[2:0] == 5) begin
        next_mux_d0_176 = input_word_d[1413];
    end else if (sel_d0_176[2:0] == 6) begin
        next_mux_d0_176 = input_word_d[1414];
    end else begin
        next_mux_d0_176 = input_word_d[1415];
    end

    if (sel_d0_177[2:0] == 0) begin
        next_mux_d0_177 = input_word_d[1416];
    end else if (sel_d0_177[2:0] == 1) begin
        next_mux_d0_177 = input_word_d[1417];
    end else if (sel_d0_177[2:0] == 2) begin
        next_mux_d0_177 = input_word_d[1418];
    end else if (sel_d0_177[2:0] == 3) begin
        next_mux_d0_177 = input_word_d[1419];
    end else if (sel_d0_177[2:0] == 4) begin
        next_mux_d0_177 = input_word_d[1420];
    end else if (sel_d0_177[2:0] == 5) begin
        next_mux_d0_177 = input_word_d[1421];
    end else if (sel_d0_177[2:0] == 6) begin
        next_mux_d0_177 = input_word_d[1422];
    end else begin
        next_mux_d0_177 = input_word_d[1423];
    end

    if (sel_d0_178[2:0] == 0) begin
        next_mux_d0_178 = input_word_d[1424];
    end else if (sel_d0_178[2:0] == 1) begin
        next_mux_d0_178 = input_word_d[1425];
    end else if (sel_d0_178[2:0] == 2) begin
        next_mux_d0_178 = input_word_d[1426];
    end else if (sel_d0_178[2:0] == 3) begin
        next_mux_d0_178 = input_word_d[1427];
    end else if (sel_d0_178[2:0] == 4) begin
        next_mux_d0_178 = input_word_d[1428];
    end else if (sel_d0_178[2:0] == 5) begin
        next_mux_d0_178 = input_word_d[1429];
    end else if (sel_d0_178[2:0] == 6) begin
        next_mux_d0_178 = input_word_d[1430];
    end else begin
        next_mux_d0_178 = input_word_d[1431];
    end

    if (sel_d0_179[2:0] == 0) begin
        next_mux_d0_179 = input_word_d[1432];
    end else if (sel_d0_179[2:0] == 1) begin
        next_mux_d0_179 = input_word_d[1433];
    end else if (sel_d0_179[2:0] == 2) begin
        next_mux_d0_179 = input_word_d[1434];
    end else if (sel_d0_179[2:0] == 3) begin
        next_mux_d0_179 = input_word_d[1435];
    end else if (sel_d0_179[2:0] == 4) begin
        next_mux_d0_179 = input_word_d[1436];
    end else if (sel_d0_179[2:0] == 5) begin
        next_mux_d0_179 = input_word_d[1437];
    end else if (sel_d0_179[2:0] == 6) begin
        next_mux_d0_179 = input_word_d[1438];
    end else begin
        next_mux_d0_179 = input_word_d[1439];
    end

    if (sel_d0_180[2:0] == 0) begin
        next_mux_d0_180 = input_word_d[1440];
    end else if (sel_d0_180[2:0] == 1) begin
        next_mux_d0_180 = input_word_d[1441];
    end else if (sel_d0_180[2:0] == 2) begin
        next_mux_d0_180 = input_word_d[1442];
    end else if (sel_d0_180[2:0] == 3) begin
        next_mux_d0_180 = input_word_d[1443];
    end else if (sel_d0_180[2:0] == 4) begin
        next_mux_d0_180 = input_word_d[1444];
    end else if (sel_d0_180[2:0] == 5) begin
        next_mux_d0_180 = input_word_d[1445];
    end else if (sel_d0_180[2:0] == 6) begin
        next_mux_d0_180 = input_word_d[1446];
    end else begin
        next_mux_d0_180 = input_word_d[1447];
    end

    if (sel_d0_181[2:0] == 0) begin
        next_mux_d0_181 = input_word_d[1448];
    end else if (sel_d0_181[2:0] == 1) begin
        next_mux_d0_181 = input_word_d[1449];
    end else if (sel_d0_181[2:0] == 2) begin
        next_mux_d0_181 = input_word_d[1450];
    end else if (sel_d0_181[2:0] == 3) begin
        next_mux_d0_181 = input_word_d[1451];
    end else if (sel_d0_181[2:0] == 4) begin
        next_mux_d0_181 = input_word_d[1452];
    end else if (sel_d0_181[2:0] == 5) begin
        next_mux_d0_181 = input_word_d[1453];
    end else if (sel_d0_181[2:0] == 6) begin
        next_mux_d0_181 = input_word_d[1454];
    end else begin
        next_mux_d0_181 = input_word_d[1455];
    end

    if (sel_d0_182[2:0] == 0) begin
        next_mux_d0_182 = input_word_d[1456];
    end else if (sel_d0_182[2:0] == 1) begin
        next_mux_d0_182 = input_word_d[1457];
    end else if (sel_d0_182[2:0] == 2) begin
        next_mux_d0_182 = input_word_d[1458];
    end else if (sel_d0_182[2:0] == 3) begin
        next_mux_d0_182 = input_word_d[1459];
    end else if (sel_d0_182[2:0] == 4) begin
        next_mux_d0_182 = input_word_d[1460];
    end else if (sel_d0_182[2:0] == 5) begin
        next_mux_d0_182 = input_word_d[1461];
    end else if (sel_d0_182[2:0] == 6) begin
        next_mux_d0_182 = input_word_d[1462];
    end else begin
        next_mux_d0_182 = input_word_d[1463];
    end

    if (sel_d0_183[2:0] == 0) begin
        next_mux_d0_183 = input_word_d[1464];
    end else if (sel_d0_183[2:0] == 1) begin
        next_mux_d0_183 = input_word_d[1465];
    end else if (sel_d0_183[2:0] == 2) begin
        next_mux_d0_183 = input_word_d[1466];
    end else if (sel_d0_183[2:0] == 3) begin
        next_mux_d0_183 = input_word_d[1467];
    end else if (sel_d0_183[2:0] == 4) begin
        next_mux_d0_183 = input_word_d[1468];
    end else if (sel_d0_183[2:0] == 5) begin
        next_mux_d0_183 = input_word_d[1469];
    end else if (sel_d0_183[2:0] == 6) begin
        next_mux_d0_183 = input_word_d[1470];
    end else begin
        next_mux_d0_183 = input_word_d[1471];
    end

    if (sel_d0_184[2:0] == 0) begin
        next_mux_d0_184 = input_word_d[1472];
    end else if (sel_d0_184[2:0] == 1) begin
        next_mux_d0_184 = input_word_d[1473];
    end else if (sel_d0_184[2:0] == 2) begin
        next_mux_d0_184 = input_word_d[1474];
    end else if (sel_d0_184[2:0] == 3) begin
        next_mux_d0_184 = input_word_d[1475];
    end else if (sel_d0_184[2:0] == 4) begin
        next_mux_d0_184 = input_word_d[1476];
    end else if (sel_d0_184[2:0] == 5) begin
        next_mux_d0_184 = input_word_d[1477];
    end else if (sel_d0_184[2:0] == 6) begin
        next_mux_d0_184 = input_word_d[1478];
    end else begin
        next_mux_d0_184 = input_word_d[1479];
    end

    if (sel_d0_185[2:0] == 0) begin
        next_mux_d0_185 = input_word_d[1480];
    end else if (sel_d0_185[2:0] == 1) begin
        next_mux_d0_185 = input_word_d[1481];
    end else if (sel_d0_185[2:0] == 2) begin
        next_mux_d0_185 = input_word_d[1482];
    end else if (sel_d0_185[2:0] == 3) begin
        next_mux_d0_185 = input_word_d[1483];
    end else if (sel_d0_185[2:0] == 4) begin
        next_mux_d0_185 = input_word_d[1484];
    end else if (sel_d0_185[2:0] == 5) begin
        next_mux_d0_185 = input_word_d[1485];
    end else if (sel_d0_185[2:0] == 6) begin
        next_mux_d0_185 = input_word_d[1486];
    end else begin
        next_mux_d0_185 = input_word_d[1487];
    end

    if (sel_d0_186[2:0] == 0) begin
        next_mux_d0_186 = input_word_d[1488];
    end else if (sel_d0_186[2:0] == 1) begin
        next_mux_d0_186 = input_word_d[1489];
    end else if (sel_d0_186[2:0] == 2) begin
        next_mux_d0_186 = input_word_d[1490];
    end else if (sel_d0_186[2:0] == 3) begin
        next_mux_d0_186 = input_word_d[1491];
    end else if (sel_d0_186[2:0] == 4) begin
        next_mux_d0_186 = input_word_d[1492];
    end else if (sel_d0_186[2:0] == 5) begin
        next_mux_d0_186 = input_word_d[1493];
    end else if (sel_d0_186[2:0] == 6) begin
        next_mux_d0_186 = input_word_d[1494];
    end else begin
        next_mux_d0_186 = input_word_d[1495];
    end

    if (sel_d0_187[2:0] == 0) begin
        next_mux_d0_187 = input_word_d[1496];
    end else if (sel_d0_187[2:0] == 1) begin
        next_mux_d0_187 = input_word_d[1497];
    end else if (sel_d0_187[2:0] == 2) begin
        next_mux_d0_187 = input_word_d[1498];
    end else if (sel_d0_187[2:0] == 3) begin
        next_mux_d0_187 = input_word_d[1499];
    end else if (sel_d0_187[2:0] == 4) begin
        next_mux_d0_187 = input_word_d[1500];
    end else if (sel_d0_187[2:0] == 5) begin
        next_mux_d0_187 = input_word_d[1501];
    end else if (sel_d0_187[2:0] == 6) begin
        next_mux_d0_187 = input_word_d[1502];
    end else begin
        next_mux_d0_187 = input_word_d[1503];
    end

    if (sel_d0_188[2:0] == 0) begin
        next_mux_d0_188 = input_word_d[1504];
    end else if (sel_d0_188[2:0] == 1) begin
        next_mux_d0_188 = input_word_d[1505];
    end else if (sel_d0_188[2:0] == 2) begin
        next_mux_d0_188 = input_word_d[1506];
    end else if (sel_d0_188[2:0] == 3) begin
        next_mux_d0_188 = input_word_d[1507];
    end else if (sel_d0_188[2:0] == 4) begin
        next_mux_d0_188 = input_word_d[1508];
    end else if (sel_d0_188[2:0] == 5) begin
        next_mux_d0_188 = input_word_d[1509];
    end else if (sel_d0_188[2:0] == 6) begin
        next_mux_d0_188 = input_word_d[1510];
    end else begin
        next_mux_d0_188 = input_word_d[1511];
    end

    if (sel_d0_189[2:0] == 0) begin
        next_mux_d0_189 = input_word_d[1512];
    end else if (sel_d0_189[2:0] == 1) begin
        next_mux_d0_189 = input_word_d[1513];
    end else if (sel_d0_189[2:0] == 2) begin
        next_mux_d0_189 = input_word_d[1514];
    end else if (sel_d0_189[2:0] == 3) begin
        next_mux_d0_189 = input_word_d[1515];
    end else if (sel_d0_189[2:0] == 4) begin
        next_mux_d0_189 = input_word_d[1516];
    end else if (sel_d0_189[2:0] == 5) begin
        next_mux_d0_189 = input_word_d[1517];
    end else if (sel_d0_189[2:0] == 6) begin
        next_mux_d0_189 = input_word_d[1518];
    end else begin
        next_mux_d0_189 = input_word_d[1519];
    end

    if (sel_d0_190[2:0] == 0) begin
        next_mux_d0_190 = input_word_d[1520];
    end else if (sel_d0_190[2:0] == 1) begin
        next_mux_d0_190 = input_word_d[1521];
    end else if (sel_d0_190[2:0] == 2) begin
        next_mux_d0_190 = input_word_d[1522];
    end else if (sel_d0_190[2:0] == 3) begin
        next_mux_d0_190 = input_word_d[1523];
    end else if (sel_d0_190[2:0] == 4) begin
        next_mux_d0_190 = input_word_d[1524];
    end else if (sel_d0_190[2:0] == 5) begin
        next_mux_d0_190 = input_word_d[1525];
    end else if (sel_d0_190[2:0] == 6) begin
        next_mux_d0_190 = input_word_d[1526];
    end else begin
        next_mux_d0_190 = input_word_d[1527];
    end

    if (sel_d0_191[2:0] == 0) begin
        next_mux_d0_191 = input_word_d[1528];
    end else if (sel_d0_191[2:0] == 1) begin
        next_mux_d0_191 = input_word_d[1529];
    end else if (sel_d0_191[2:0] == 2) begin
        next_mux_d0_191 = input_word_d[1530];
    end else if (sel_d0_191[2:0] == 3) begin
        next_mux_d0_191 = input_word_d[1531];
    end else if (sel_d0_191[2:0] == 4) begin
        next_mux_d0_191 = input_word_d[1532];
    end else if (sel_d0_191[2:0] == 5) begin
        next_mux_d0_191 = input_word_d[1533];
    end else if (sel_d0_191[2:0] == 6) begin
        next_mux_d0_191 = input_word_d[1534];
    end else begin
        next_mux_d0_191 = input_word_d[1535];
    end

    if (sel_d0_192[2:0] == 0) begin
        next_mux_d0_192 = input_word_d[1536];
    end else if (sel_d0_192[2:0] == 1) begin
        next_mux_d0_192 = input_word_d[1537];
    end else if (sel_d0_192[2:0] == 2) begin
        next_mux_d0_192 = input_word_d[1538];
    end else if (sel_d0_192[2:0] == 3) begin
        next_mux_d0_192 = input_word_d[1539];
    end else if (sel_d0_192[2:0] == 4) begin
        next_mux_d0_192 = input_word_d[1540];
    end else if (sel_d0_192[2:0] == 5) begin
        next_mux_d0_192 = input_word_d[1541];
    end else if (sel_d0_192[2:0] == 6) begin
        next_mux_d0_192 = input_word_d[1542];
    end else begin
        next_mux_d0_192 = input_word_d[1543];
    end

    if (sel_d0_193[2:0] == 0) begin
        next_mux_d0_193 = input_word_d[1544];
    end else if (sel_d0_193[2:0] == 1) begin
        next_mux_d0_193 = input_word_d[1545];
    end else if (sel_d0_193[2:0] == 2) begin
        next_mux_d0_193 = input_word_d[1546];
    end else if (sel_d0_193[2:0] == 3) begin
        next_mux_d0_193 = input_word_d[1547];
    end else if (sel_d0_193[2:0] == 4) begin
        next_mux_d0_193 = input_word_d[1548];
    end else if (sel_d0_193[2:0] == 5) begin
        next_mux_d0_193 = input_word_d[1549];
    end else if (sel_d0_193[2:0] == 6) begin
        next_mux_d0_193 = input_word_d[1550];
    end else begin
        next_mux_d0_193 = input_word_d[1551];
    end

    if (sel_d0_194[2:0] == 0) begin
        next_mux_d0_194 = input_word_d[1552];
    end else if (sel_d0_194[2:0] == 1) begin
        next_mux_d0_194 = input_word_d[1553];
    end else if (sel_d0_194[2:0] == 2) begin
        next_mux_d0_194 = input_word_d[1554];
    end else if (sel_d0_194[2:0] == 3) begin
        next_mux_d0_194 = input_word_d[1555];
    end else if (sel_d0_194[2:0] == 4) begin
        next_mux_d0_194 = input_word_d[1556];
    end else if (sel_d0_194[2:0] == 5) begin
        next_mux_d0_194 = input_word_d[1557];
    end else if (sel_d0_194[2:0] == 6) begin
        next_mux_d0_194 = input_word_d[1558];
    end else begin
        next_mux_d0_194 = input_word_d[1559];
    end

    if (sel_d0_195[2:0] == 0) begin
        next_mux_d0_195 = input_word_d[1560];
    end else if (sel_d0_195[2:0] == 1) begin
        next_mux_d0_195 = input_word_d[1561];
    end else if (sel_d0_195[2:0] == 2) begin
        next_mux_d0_195 = input_word_d[1562];
    end else if (sel_d0_195[2:0] == 3) begin
        next_mux_d0_195 = input_word_d[1563];
    end else if (sel_d0_195[2:0] == 4) begin
        next_mux_d0_195 = input_word_d[1564];
    end else if (sel_d0_195[2:0] == 5) begin
        next_mux_d0_195 = input_word_d[1565];
    end else if (sel_d0_195[2:0] == 6) begin
        next_mux_d0_195 = input_word_d[1566];
    end else begin
        next_mux_d0_195 = input_word_d[1567];
    end

    if (sel_d0_196[2:0] == 0) begin
        next_mux_d0_196 = input_word_d[1568];
    end else if (sel_d0_196[2:0] == 1) begin
        next_mux_d0_196 = input_word_d[1569];
    end else if (sel_d0_196[2:0] == 2) begin
        next_mux_d0_196 = input_word_d[1570];
    end else if (sel_d0_196[2:0] == 3) begin
        next_mux_d0_196 = input_word_d[1571];
    end else if (sel_d0_196[2:0] == 4) begin
        next_mux_d0_196 = input_word_d[1572];
    end else if (sel_d0_196[2:0] == 5) begin
        next_mux_d0_196 = input_word_d[1573];
    end else if (sel_d0_196[2:0] == 6) begin
        next_mux_d0_196 = input_word_d[1574];
    end else begin
        next_mux_d0_196 = input_word_d[1575];
    end

    if (sel_d0_197[2:0] == 0) begin
        next_mux_d0_197 = input_word_d[1576];
    end else if (sel_d0_197[2:0] == 1) begin
        next_mux_d0_197 = input_word_d[1577];
    end else if (sel_d0_197[2:0] == 2) begin
        next_mux_d0_197 = input_word_d[1578];
    end else if (sel_d0_197[2:0] == 3) begin
        next_mux_d0_197 = input_word_d[1579];
    end else if (sel_d0_197[2:0] == 4) begin
        next_mux_d0_197 = input_word_d[1580];
    end else if (sel_d0_197[2:0] == 5) begin
        next_mux_d0_197 = input_word_d[1581];
    end else if (sel_d0_197[2:0] == 6) begin
        next_mux_d0_197 = input_word_d[1582];
    end else begin
        next_mux_d0_197 = input_word_d[1583];
    end

    if (sel_d0_198[2:0] == 0) begin
        next_mux_d0_198 = input_word_d[1584];
    end else if (sel_d0_198[2:0] == 1) begin
        next_mux_d0_198 = input_word_d[1585];
    end else if (sel_d0_198[2:0] == 2) begin
        next_mux_d0_198 = input_word_d[1586];
    end else if (sel_d0_198[2:0] == 3) begin
        next_mux_d0_198 = input_word_d[1587];
    end else if (sel_d0_198[2:0] == 4) begin
        next_mux_d0_198 = input_word_d[1588];
    end else if (sel_d0_198[2:0] == 5) begin
        next_mux_d0_198 = input_word_d[1589];
    end else if (sel_d0_198[2:0] == 6) begin
        next_mux_d0_198 = input_word_d[1590];
    end else begin
        next_mux_d0_198 = input_word_d[1591];
    end

    if (sel_d0_199[2:0] == 0) begin
        next_mux_d0_199 = input_word_d[1592];
    end else if (sel_d0_199[2:0] == 1) begin
        next_mux_d0_199 = input_word_d[1593];
    end else if (sel_d0_199[2:0] == 2) begin
        next_mux_d0_199 = input_word_d[1594];
    end else if (sel_d0_199[2:0] == 3) begin
        next_mux_d0_199 = input_word_d[1595];
    end else if (sel_d0_199[2:0] == 4) begin
        next_mux_d0_199 = input_word_d[1596];
    end else if (sel_d0_199[2:0] == 5) begin
        next_mux_d0_199 = input_word_d[1597];
    end else if (sel_d0_199[2:0] == 6) begin
        next_mux_d0_199 = input_word_d[1598];
    end else begin
        next_mux_d0_199 = input_word_d[1599];
    end

    if (sel_d0_200[2:0] == 0) begin
        next_mux_d0_200 = input_word_d[1600];
    end else if (sel_d0_200[2:0] == 1) begin
        next_mux_d0_200 = input_word_d[1601];
    end else if (sel_d0_200[2:0] == 2) begin
        next_mux_d0_200 = input_word_d[1602];
    end else if (sel_d0_200[2:0] == 3) begin
        next_mux_d0_200 = input_word_d[1603];
    end else if (sel_d0_200[2:0] == 4) begin
        next_mux_d0_200 = input_word_d[1604];
    end else if (sel_d0_200[2:0] == 5) begin
        next_mux_d0_200 = input_word_d[1605];
    end else if (sel_d0_200[2:0] == 6) begin
        next_mux_d0_200 = input_word_d[1606];
    end else begin
        next_mux_d0_200 = input_word_d[1607];
    end

    if (sel_d0_201[2:0] == 0) begin
        next_mux_d0_201 = input_word_d[1608];
    end else if (sel_d0_201[2:0] == 1) begin
        next_mux_d0_201 = input_word_d[1609];
    end else if (sel_d0_201[2:0] == 2) begin
        next_mux_d0_201 = input_word_d[1610];
    end else if (sel_d0_201[2:0] == 3) begin
        next_mux_d0_201 = input_word_d[1611];
    end else if (sel_d0_201[2:0] == 4) begin
        next_mux_d0_201 = input_word_d[1612];
    end else if (sel_d0_201[2:0] == 5) begin
        next_mux_d0_201 = input_word_d[1613];
    end else if (sel_d0_201[2:0] == 6) begin
        next_mux_d0_201 = input_word_d[1614];
    end else begin
        next_mux_d0_201 = input_word_d[1615];
    end

    if (sel_d0_202[2:0] == 0) begin
        next_mux_d0_202 = input_word_d[1616];
    end else if (sel_d0_202[2:0] == 1) begin
        next_mux_d0_202 = input_word_d[1617];
    end else if (sel_d0_202[2:0] == 2) begin
        next_mux_d0_202 = input_word_d[1618];
    end else if (sel_d0_202[2:0] == 3) begin
        next_mux_d0_202 = input_word_d[1619];
    end else if (sel_d0_202[2:0] == 4) begin
        next_mux_d0_202 = input_word_d[1620];
    end else if (sel_d0_202[2:0] == 5) begin
        next_mux_d0_202 = input_word_d[1621];
    end else if (sel_d0_202[2:0] == 6) begin
        next_mux_d0_202 = input_word_d[1622];
    end else begin
        next_mux_d0_202 = input_word_d[1623];
    end

    if (sel_d0_203[2:0] == 0) begin
        next_mux_d0_203 = input_word_d[1624];
    end else if (sel_d0_203[2:0] == 1) begin
        next_mux_d0_203 = input_word_d[1625];
    end else if (sel_d0_203[2:0] == 2) begin
        next_mux_d0_203 = input_word_d[1626];
    end else if (sel_d0_203[2:0] == 3) begin
        next_mux_d0_203 = input_word_d[1627];
    end else if (sel_d0_203[2:0] == 4) begin
        next_mux_d0_203 = input_word_d[1628];
    end else if (sel_d0_203[2:0] == 5) begin
        next_mux_d0_203 = input_word_d[1629];
    end else if (sel_d0_203[2:0] == 6) begin
        next_mux_d0_203 = input_word_d[1630];
    end else begin
        next_mux_d0_203 = input_word_d[1631];
    end

    if (sel_d0_204[2:0] == 0) begin
        next_mux_d0_204 = input_word_d[1632];
    end else if (sel_d0_204[2:0] == 1) begin
        next_mux_d0_204 = input_word_d[1633];
    end else if (sel_d0_204[2:0] == 2) begin
        next_mux_d0_204 = input_word_d[1634];
    end else if (sel_d0_204[2:0] == 3) begin
        next_mux_d0_204 = input_word_d[1635];
    end else if (sel_d0_204[2:0] == 4) begin
        next_mux_d0_204 = input_word_d[1636];
    end else if (sel_d0_204[2:0] == 5) begin
        next_mux_d0_204 = input_word_d[1637];
    end else if (sel_d0_204[2:0] == 6) begin
        next_mux_d0_204 = input_word_d[1638];
    end else begin
        next_mux_d0_204 = input_word_d[1639];
    end

    if (sel_d0_205[2:0] == 0) begin
        next_mux_d0_205 = input_word_d[1640];
    end else if (sel_d0_205[2:0] == 1) begin
        next_mux_d0_205 = input_word_d[1641];
    end else if (sel_d0_205[2:0] == 2) begin
        next_mux_d0_205 = input_word_d[1642];
    end else if (sel_d0_205[2:0] == 3) begin
        next_mux_d0_205 = input_word_d[1643];
    end else if (sel_d0_205[2:0] == 4) begin
        next_mux_d0_205 = input_word_d[1644];
    end else if (sel_d0_205[2:0] == 5) begin
        next_mux_d0_205 = input_word_d[1645];
    end else if (sel_d0_205[2:0] == 6) begin
        next_mux_d0_205 = input_word_d[1646];
    end else begin
        next_mux_d0_205 = input_word_d[1647];
    end

    if (sel_d0_206[2:0] == 0) begin
        next_mux_d0_206 = input_word_d[1648];
    end else if (sel_d0_206[2:0] == 1) begin
        next_mux_d0_206 = input_word_d[1649];
    end else if (sel_d0_206[2:0] == 2) begin
        next_mux_d0_206 = input_word_d[1650];
    end else if (sel_d0_206[2:0] == 3) begin
        next_mux_d0_206 = input_word_d[1651];
    end else if (sel_d0_206[2:0] == 4) begin
        next_mux_d0_206 = input_word_d[1652];
    end else if (sel_d0_206[2:0] == 5) begin
        next_mux_d0_206 = input_word_d[1653];
    end else if (sel_d0_206[2:0] == 6) begin
        next_mux_d0_206 = input_word_d[1654];
    end else begin
        next_mux_d0_206 = input_word_d[1655];
    end

    if (sel_d0_207[2:0] == 0) begin
        next_mux_d0_207 = input_word_d[1656];
    end else if (sel_d0_207[2:0] == 1) begin
        next_mux_d0_207 = input_word_d[1657];
    end else if (sel_d0_207[2:0] == 2) begin
        next_mux_d0_207 = input_word_d[1658];
    end else if (sel_d0_207[2:0] == 3) begin
        next_mux_d0_207 = input_word_d[1659];
    end else if (sel_d0_207[2:0] == 4) begin
        next_mux_d0_207 = input_word_d[1660];
    end else if (sel_d0_207[2:0] == 5) begin
        next_mux_d0_207 = input_word_d[1661];
    end else if (sel_d0_207[2:0] == 6) begin
        next_mux_d0_207 = input_word_d[1662];
    end else begin
        next_mux_d0_207 = input_word_d[1663];
    end

    if (sel_d0_208[2:0] == 0) begin
        next_mux_d0_208 = input_word_d[1664];
    end else if (sel_d0_208[2:0] == 1) begin
        next_mux_d0_208 = input_word_d[1665];
    end else if (sel_d0_208[2:0] == 2) begin
        next_mux_d0_208 = input_word_d[1666];
    end else if (sel_d0_208[2:0] == 3) begin
        next_mux_d0_208 = input_word_d[1667];
    end else if (sel_d0_208[2:0] == 4) begin
        next_mux_d0_208 = input_word_d[1668];
    end else if (sel_d0_208[2:0] == 5) begin
        next_mux_d0_208 = input_word_d[1669];
    end else if (sel_d0_208[2:0] == 6) begin
        next_mux_d0_208 = input_word_d[1670];
    end else begin
        next_mux_d0_208 = input_word_d[1671];
    end

    if (sel_d0_209[2:0] == 0) begin
        next_mux_d0_209 = input_word_d[1672];
    end else if (sel_d0_209[2:0] == 1) begin
        next_mux_d0_209 = input_word_d[1673];
    end else if (sel_d0_209[2:0] == 2) begin
        next_mux_d0_209 = input_word_d[1674];
    end else if (sel_d0_209[2:0] == 3) begin
        next_mux_d0_209 = input_word_d[1675];
    end else if (sel_d0_209[2:0] == 4) begin
        next_mux_d0_209 = input_word_d[1676];
    end else if (sel_d0_209[2:0] == 5) begin
        next_mux_d0_209 = input_word_d[1677];
    end else if (sel_d0_209[2:0] == 6) begin
        next_mux_d0_209 = input_word_d[1678];
    end else begin
        next_mux_d0_209 = input_word_d[1679];
    end

    if (sel_d0_210[2:0] == 0) begin
        next_mux_d0_210 = input_word_d[1680];
    end else if (sel_d0_210[2:0] == 1) begin
        next_mux_d0_210 = input_word_d[1681];
    end else if (sel_d0_210[2:0] == 2) begin
        next_mux_d0_210 = input_word_d[1682];
    end else if (sel_d0_210[2:0] == 3) begin
        next_mux_d0_210 = input_word_d[1683];
    end else if (sel_d0_210[2:0] == 4) begin
        next_mux_d0_210 = input_word_d[1684];
    end else if (sel_d0_210[2:0] == 5) begin
        next_mux_d0_210 = input_word_d[1685];
    end else if (sel_d0_210[2:0] == 6) begin
        next_mux_d0_210 = input_word_d[1686];
    end else begin
        next_mux_d0_210 = input_word_d[1687];
    end

    if (sel_d0_211[2:0] == 0) begin
        next_mux_d0_211 = input_word_d[1688];
    end else if (sel_d0_211[2:0] == 1) begin
        next_mux_d0_211 = input_word_d[1689];
    end else if (sel_d0_211[2:0] == 2) begin
        next_mux_d0_211 = input_word_d[1690];
    end else if (sel_d0_211[2:0] == 3) begin
        next_mux_d0_211 = input_word_d[1691];
    end else if (sel_d0_211[2:0] == 4) begin
        next_mux_d0_211 = input_word_d[1692];
    end else if (sel_d0_211[2:0] == 5) begin
        next_mux_d0_211 = input_word_d[1693];
    end else if (sel_d0_211[2:0] == 6) begin
        next_mux_d0_211 = input_word_d[1694];
    end else begin
        next_mux_d0_211 = input_word_d[1695];
    end

    if (sel_d0_212[2:0] == 0) begin
        next_mux_d0_212 = input_word_d[1696];
    end else if (sel_d0_212[2:0] == 1) begin
        next_mux_d0_212 = input_word_d[1697];
    end else if (sel_d0_212[2:0] == 2) begin
        next_mux_d0_212 = input_word_d[1698];
    end else if (sel_d0_212[2:0] == 3) begin
        next_mux_d0_212 = input_word_d[1699];
    end else if (sel_d0_212[2:0] == 4) begin
        next_mux_d0_212 = input_word_d[1700];
    end else if (sel_d0_212[2:0] == 5) begin
        next_mux_d0_212 = input_word_d[1701];
    end else if (sel_d0_212[2:0] == 6) begin
        next_mux_d0_212 = input_word_d[1702];
    end else begin
        next_mux_d0_212 = input_word_d[1703];
    end

    if (sel_d0_213[2:0] == 0) begin
        next_mux_d0_213 = input_word_d[1704];
    end else if (sel_d0_213[2:0] == 1) begin
        next_mux_d0_213 = input_word_d[1705];
    end else if (sel_d0_213[2:0] == 2) begin
        next_mux_d0_213 = input_word_d[1706];
    end else if (sel_d0_213[2:0] == 3) begin
        next_mux_d0_213 = input_word_d[1707];
    end else if (sel_d0_213[2:0] == 4) begin
        next_mux_d0_213 = input_word_d[1708];
    end else if (sel_d0_213[2:0] == 5) begin
        next_mux_d0_213 = input_word_d[1709];
    end else if (sel_d0_213[2:0] == 6) begin
        next_mux_d0_213 = input_word_d[1710];
    end else begin
        next_mux_d0_213 = input_word_d[1711];
    end

    if (sel_d0_214[2:0] == 0) begin
        next_mux_d0_214 = input_word_d[1712];
    end else if (sel_d0_214[2:0] == 1) begin
        next_mux_d0_214 = input_word_d[1713];
    end else if (sel_d0_214[2:0] == 2) begin
        next_mux_d0_214 = input_word_d[1714];
    end else if (sel_d0_214[2:0] == 3) begin
        next_mux_d0_214 = input_word_d[1715];
    end else if (sel_d0_214[2:0] == 4) begin
        next_mux_d0_214 = input_word_d[1716];
    end else if (sel_d0_214[2:0] == 5) begin
        next_mux_d0_214 = input_word_d[1717];
    end else if (sel_d0_214[2:0] == 6) begin
        next_mux_d0_214 = input_word_d[1718];
    end else begin
        next_mux_d0_214 = input_word_d[1719];
    end

    if (sel_d0_215[2:0] == 0) begin
        next_mux_d0_215 = input_word_d[1720];
    end else if (sel_d0_215[2:0] == 1) begin
        next_mux_d0_215 = input_word_d[1721];
    end else if (sel_d0_215[2:0] == 2) begin
        next_mux_d0_215 = input_word_d[1722];
    end else if (sel_d0_215[2:0] == 3) begin
        next_mux_d0_215 = input_word_d[1723];
    end else if (sel_d0_215[2:0] == 4) begin
        next_mux_d0_215 = input_word_d[1724];
    end else if (sel_d0_215[2:0] == 5) begin
        next_mux_d0_215 = input_word_d[1725];
    end else if (sel_d0_215[2:0] == 6) begin
        next_mux_d0_215 = input_word_d[1726];
    end else begin
        next_mux_d0_215 = input_word_d[1727];
    end

    if (sel_d0_216[2:0] == 0) begin
        next_mux_d0_216 = input_word_d[1728];
    end else if (sel_d0_216[2:0] == 1) begin
        next_mux_d0_216 = input_word_d[1729];
    end else if (sel_d0_216[2:0] == 2) begin
        next_mux_d0_216 = input_word_d[1730];
    end else if (sel_d0_216[2:0] == 3) begin
        next_mux_d0_216 = input_word_d[1731];
    end else if (sel_d0_216[2:0] == 4) begin
        next_mux_d0_216 = input_word_d[1732];
    end else if (sel_d0_216[2:0] == 5) begin
        next_mux_d0_216 = input_word_d[1733];
    end else if (sel_d0_216[2:0] == 6) begin
        next_mux_d0_216 = input_word_d[1734];
    end else begin
        next_mux_d0_216 = input_word_d[1735];
    end

    if (sel_d0_217[2:0] == 0) begin
        next_mux_d0_217 = input_word_d[1736];
    end else if (sel_d0_217[2:0] == 1) begin
        next_mux_d0_217 = input_word_d[1737];
    end else if (sel_d0_217[2:0] == 2) begin
        next_mux_d0_217 = input_word_d[1738];
    end else if (sel_d0_217[2:0] == 3) begin
        next_mux_d0_217 = input_word_d[1739];
    end else if (sel_d0_217[2:0] == 4) begin
        next_mux_d0_217 = input_word_d[1740];
    end else if (sel_d0_217[2:0] == 5) begin
        next_mux_d0_217 = input_word_d[1741];
    end else if (sel_d0_217[2:0] == 6) begin
        next_mux_d0_217 = input_word_d[1742];
    end else begin
        next_mux_d0_217 = input_word_d[1743];
    end

    if (sel_d0_218[2:0] == 0) begin
        next_mux_d0_218 = input_word_d[1744];
    end else if (sel_d0_218[2:0] == 1) begin
        next_mux_d0_218 = input_word_d[1745];
    end else if (sel_d0_218[2:0] == 2) begin
        next_mux_d0_218 = input_word_d[1746];
    end else if (sel_d0_218[2:0] == 3) begin
        next_mux_d0_218 = input_word_d[1747];
    end else if (sel_d0_218[2:0] == 4) begin
        next_mux_d0_218 = input_word_d[1748];
    end else if (sel_d0_218[2:0] == 5) begin
        next_mux_d0_218 = input_word_d[1749];
    end else if (sel_d0_218[2:0] == 6) begin
        next_mux_d0_218 = input_word_d[1750];
    end else begin
        next_mux_d0_218 = input_word_d[1751];
    end

    if (sel_d0_219[2:0] == 0) begin
        next_mux_d0_219 = input_word_d[1752];
    end else if (sel_d0_219[2:0] == 1) begin
        next_mux_d0_219 = input_word_d[1753];
    end else if (sel_d0_219[2:0] == 2) begin
        next_mux_d0_219 = input_word_d[1754];
    end else if (sel_d0_219[2:0] == 3) begin
        next_mux_d0_219 = input_word_d[1755];
    end else if (sel_d0_219[2:0] == 4) begin
        next_mux_d0_219 = input_word_d[1756];
    end else if (sel_d0_219[2:0] == 5) begin
        next_mux_d0_219 = input_word_d[1757];
    end else if (sel_d0_219[2:0] == 6) begin
        next_mux_d0_219 = input_word_d[1758];
    end else begin
        next_mux_d0_219 = input_word_d[1759];
    end

    if (sel_d0_220[2:0] == 0) begin
        next_mux_d0_220 = input_word_d[1760];
    end else if (sel_d0_220[2:0] == 1) begin
        next_mux_d0_220 = input_word_d[1761];
    end else if (sel_d0_220[2:0] == 2) begin
        next_mux_d0_220 = input_word_d[1762];
    end else if (sel_d0_220[2:0] == 3) begin
        next_mux_d0_220 = input_word_d[1763];
    end else if (sel_d0_220[2:0] == 4) begin
        next_mux_d0_220 = input_word_d[1764];
    end else if (sel_d0_220[2:0] == 5) begin
        next_mux_d0_220 = input_word_d[1765];
    end else if (sel_d0_220[2:0] == 6) begin
        next_mux_d0_220 = input_word_d[1766];
    end else begin
        next_mux_d0_220 = input_word_d[1767];
    end

    if (sel_d0_221[2:0] == 0) begin
        next_mux_d0_221 = input_word_d[1768];
    end else if (sel_d0_221[2:0] == 1) begin
        next_mux_d0_221 = input_word_d[1769];
    end else if (sel_d0_221[2:0] == 2) begin
        next_mux_d0_221 = input_word_d[1770];
    end else if (sel_d0_221[2:0] == 3) begin
        next_mux_d0_221 = input_word_d[1771];
    end else if (sel_d0_221[2:0] == 4) begin
        next_mux_d0_221 = input_word_d[1772];
    end else if (sel_d0_221[2:0] == 5) begin
        next_mux_d0_221 = input_word_d[1773];
    end else if (sel_d0_221[2:0] == 6) begin
        next_mux_d0_221 = input_word_d[1774];
    end else begin
        next_mux_d0_221 = input_word_d[1775];
    end

    if (sel_d0_222[2:0] == 0) begin
        next_mux_d0_222 = input_word_d[1776];
    end else if (sel_d0_222[2:0] == 1) begin
        next_mux_d0_222 = input_word_d[1777];
    end else if (sel_d0_222[2:0] == 2) begin
        next_mux_d0_222 = input_word_d[1778];
    end else if (sel_d0_222[2:0] == 3) begin
        next_mux_d0_222 = input_word_d[1779];
    end else if (sel_d0_222[2:0] == 4) begin
        next_mux_d0_222 = input_word_d[1780];
    end else if (sel_d0_222[2:0] == 5) begin
        next_mux_d0_222 = input_word_d[1781];
    end else if (sel_d0_222[2:0] == 6) begin
        next_mux_d0_222 = input_word_d[1782];
    end else begin
        next_mux_d0_222 = input_word_d[1783];
    end

    if (sel_d0_223[2:0] == 0) begin
        next_mux_d0_223 = input_word_d[1784];
    end else if (sel_d0_223[2:0] == 1) begin
        next_mux_d0_223 = input_word_d[1785];
    end else if (sel_d0_223[2:0] == 2) begin
        next_mux_d0_223 = input_word_d[1786];
    end else if (sel_d0_223[2:0] == 3) begin
        next_mux_d0_223 = input_word_d[1787];
    end else if (sel_d0_223[2:0] == 4) begin
        next_mux_d0_223 = input_word_d[1788];
    end else if (sel_d0_223[2:0] == 5) begin
        next_mux_d0_223 = input_word_d[1789];
    end else if (sel_d0_223[2:0] == 6) begin
        next_mux_d0_223 = input_word_d[1790];
    end else begin
        next_mux_d0_223 = input_word_d[1791];
    end

    if (sel_d0_224[2:0] == 0) begin
        next_mux_d0_224 = input_word_d[1792];
    end else if (sel_d0_224[2:0] == 1) begin
        next_mux_d0_224 = input_word_d[1793];
    end else if (sel_d0_224[2:0] == 2) begin
        next_mux_d0_224 = input_word_d[1794];
    end else if (sel_d0_224[2:0] == 3) begin
        next_mux_d0_224 = input_word_d[1795];
    end else if (sel_d0_224[2:0] == 4) begin
        next_mux_d0_224 = input_word_d[1796];
    end else if (sel_d0_224[2:0] == 5) begin
        next_mux_d0_224 = input_word_d[1797];
    end else if (sel_d0_224[2:0] == 6) begin
        next_mux_d0_224 = input_word_d[1798];
    end else begin
        next_mux_d0_224 = input_word_d[1799];
    end

    if (sel_d0_225[2:0] == 0) begin
        next_mux_d0_225 = input_word_d[1800];
    end else if (sel_d0_225[2:0] == 1) begin
        next_mux_d0_225 = input_word_d[1801];
    end else if (sel_d0_225[2:0] == 2) begin
        next_mux_d0_225 = input_word_d[1802];
    end else if (sel_d0_225[2:0] == 3) begin
        next_mux_d0_225 = input_word_d[1803];
    end else if (sel_d0_225[2:0] == 4) begin
        next_mux_d0_225 = input_word_d[1804];
    end else if (sel_d0_225[2:0] == 5) begin
        next_mux_d0_225 = input_word_d[1805];
    end else if (sel_d0_225[2:0] == 6) begin
        next_mux_d0_225 = input_word_d[1806];
    end else begin
        next_mux_d0_225 = input_word_d[1807];
    end

    if (sel_d0_226[2:0] == 0) begin
        next_mux_d0_226 = input_word_d[1808];
    end else if (sel_d0_226[2:0] == 1) begin
        next_mux_d0_226 = input_word_d[1809];
    end else if (sel_d0_226[2:0] == 2) begin
        next_mux_d0_226 = input_word_d[1810];
    end else if (sel_d0_226[2:0] == 3) begin
        next_mux_d0_226 = input_word_d[1811];
    end else if (sel_d0_226[2:0] == 4) begin
        next_mux_d0_226 = input_word_d[1812];
    end else if (sel_d0_226[2:0] == 5) begin
        next_mux_d0_226 = input_word_d[1813];
    end else if (sel_d0_226[2:0] == 6) begin
        next_mux_d0_226 = input_word_d[1814];
    end else begin
        next_mux_d0_226 = input_word_d[1815];
    end

    if (sel_d0_227[2:0] == 0) begin
        next_mux_d0_227 = input_word_d[1816];
    end else if (sel_d0_227[2:0] == 1) begin
        next_mux_d0_227 = input_word_d[1817];
    end else if (sel_d0_227[2:0] == 2) begin
        next_mux_d0_227 = input_word_d[1818];
    end else if (sel_d0_227[2:0] == 3) begin
        next_mux_d0_227 = input_word_d[1819];
    end else if (sel_d0_227[2:0] == 4) begin
        next_mux_d0_227 = input_word_d[1820];
    end else if (sel_d0_227[2:0] == 5) begin
        next_mux_d0_227 = input_word_d[1821];
    end else if (sel_d0_227[2:0] == 6) begin
        next_mux_d0_227 = input_word_d[1822];
    end else begin
        next_mux_d0_227 = input_word_d[1823];
    end

    if (sel_d0_228[2:0] == 0) begin
        next_mux_d0_228 = input_word_d[1824];
    end else if (sel_d0_228[2:0] == 1) begin
        next_mux_d0_228 = input_word_d[1825];
    end else if (sel_d0_228[2:0] == 2) begin
        next_mux_d0_228 = input_word_d[1826];
    end else if (sel_d0_228[2:0] == 3) begin
        next_mux_d0_228 = input_word_d[1827];
    end else if (sel_d0_228[2:0] == 4) begin
        next_mux_d0_228 = input_word_d[1828];
    end else if (sel_d0_228[2:0] == 5) begin
        next_mux_d0_228 = input_word_d[1829];
    end else if (sel_d0_228[2:0] == 6) begin
        next_mux_d0_228 = input_word_d[1830];
    end else begin
        next_mux_d0_228 = input_word_d[1831];
    end

    if (sel_d0_229[2:0] == 0) begin
        next_mux_d0_229 = input_word_d[1832];
    end else if (sel_d0_229[2:0] == 1) begin
        next_mux_d0_229 = input_word_d[1833];
    end else if (sel_d0_229[2:0] == 2) begin
        next_mux_d0_229 = input_word_d[1834];
    end else if (sel_d0_229[2:0] == 3) begin
        next_mux_d0_229 = input_word_d[1835];
    end else if (sel_d0_229[2:0] == 4) begin
        next_mux_d0_229 = input_word_d[1836];
    end else if (sel_d0_229[2:0] == 5) begin
        next_mux_d0_229 = input_word_d[1837];
    end else if (sel_d0_229[2:0] == 6) begin
        next_mux_d0_229 = input_word_d[1838];
    end else begin
        next_mux_d0_229 = input_word_d[1839];
    end

    if (sel_d0_230[2:0] == 0) begin
        next_mux_d0_230 = input_word_d[1840];
    end else if (sel_d0_230[2:0] == 1) begin
        next_mux_d0_230 = input_word_d[1841];
    end else if (sel_d0_230[2:0] == 2) begin
        next_mux_d0_230 = input_word_d[1842];
    end else if (sel_d0_230[2:0] == 3) begin
        next_mux_d0_230 = input_word_d[1843];
    end else if (sel_d0_230[2:0] == 4) begin
        next_mux_d0_230 = input_word_d[1844];
    end else if (sel_d0_230[2:0] == 5) begin
        next_mux_d0_230 = input_word_d[1845];
    end else if (sel_d0_230[2:0] == 6) begin
        next_mux_d0_230 = input_word_d[1846];
    end else begin
        next_mux_d0_230 = input_word_d[1847];
    end

    if (sel_d0_231[2:0] == 0) begin
        next_mux_d0_231 = input_word_d[1848];
    end else if (sel_d0_231[2:0] == 1) begin
        next_mux_d0_231 = input_word_d[1849];
    end else if (sel_d0_231[2:0] == 2) begin
        next_mux_d0_231 = input_word_d[1850];
    end else if (sel_d0_231[2:0] == 3) begin
        next_mux_d0_231 = input_word_d[1851];
    end else if (sel_d0_231[2:0] == 4) begin
        next_mux_d0_231 = input_word_d[1852];
    end else if (sel_d0_231[2:0] == 5) begin
        next_mux_d0_231 = input_word_d[1853];
    end else if (sel_d0_231[2:0] == 6) begin
        next_mux_d0_231 = input_word_d[1854];
    end else begin
        next_mux_d0_231 = input_word_d[1855];
    end

    if (sel_d0_232[2:0] == 0) begin
        next_mux_d0_232 = input_word_d[1856];
    end else if (sel_d0_232[2:0] == 1) begin
        next_mux_d0_232 = input_word_d[1857];
    end else if (sel_d0_232[2:0] == 2) begin
        next_mux_d0_232 = input_word_d[1858];
    end else if (sel_d0_232[2:0] == 3) begin
        next_mux_d0_232 = input_word_d[1859];
    end else if (sel_d0_232[2:0] == 4) begin
        next_mux_d0_232 = input_word_d[1860];
    end else if (sel_d0_232[2:0] == 5) begin
        next_mux_d0_232 = input_word_d[1861];
    end else if (sel_d0_232[2:0] == 6) begin
        next_mux_d0_232 = input_word_d[1862];
    end else begin
        next_mux_d0_232 = input_word_d[1863];
    end

    if (sel_d0_233[2:0] == 0) begin
        next_mux_d0_233 = input_word_d[1864];
    end else if (sel_d0_233[2:0] == 1) begin
        next_mux_d0_233 = input_word_d[1865];
    end else if (sel_d0_233[2:0] == 2) begin
        next_mux_d0_233 = input_word_d[1866];
    end else if (sel_d0_233[2:0] == 3) begin
        next_mux_d0_233 = input_word_d[1867];
    end else if (sel_d0_233[2:0] == 4) begin
        next_mux_d0_233 = input_word_d[1868];
    end else if (sel_d0_233[2:0] == 5) begin
        next_mux_d0_233 = input_word_d[1869];
    end else if (sel_d0_233[2:0] == 6) begin
        next_mux_d0_233 = input_word_d[1870];
    end else begin
        next_mux_d0_233 = input_word_d[1871];
    end

    if (sel_d0_234[2:0] == 0) begin
        next_mux_d0_234 = input_word_d[1872];
    end else if (sel_d0_234[2:0] == 1) begin
        next_mux_d0_234 = input_word_d[1873];
    end else if (sel_d0_234[2:0] == 2) begin
        next_mux_d0_234 = input_word_d[1874];
    end else if (sel_d0_234[2:0] == 3) begin
        next_mux_d0_234 = input_word_d[1875];
    end else if (sel_d0_234[2:0] == 4) begin
        next_mux_d0_234 = input_word_d[1876];
    end else if (sel_d0_234[2:0] == 5) begin
        next_mux_d0_234 = input_word_d[1877];
    end else if (sel_d0_234[2:0] == 6) begin
        next_mux_d0_234 = input_word_d[1878];
    end else begin
        next_mux_d0_234 = input_word_d[1879];
    end

    if (sel_d0_235[2:0] == 0) begin
        next_mux_d0_235 = input_word_d[1880];
    end else if (sel_d0_235[2:0] == 1) begin
        next_mux_d0_235 = input_word_d[1881];
    end else if (sel_d0_235[2:0] == 2) begin
        next_mux_d0_235 = input_word_d[1882];
    end else if (sel_d0_235[2:0] == 3) begin
        next_mux_d0_235 = input_word_d[1883];
    end else if (sel_d0_235[2:0] == 4) begin
        next_mux_d0_235 = input_word_d[1884];
    end else if (sel_d0_235[2:0] == 5) begin
        next_mux_d0_235 = input_word_d[1885];
    end else if (sel_d0_235[2:0] == 6) begin
        next_mux_d0_235 = input_word_d[1886];
    end else begin
        next_mux_d0_235 = input_word_d[1887];
    end

    if (sel_d0_236[2:0] == 0) begin
        next_mux_d0_236 = input_word_d[1888];
    end else if (sel_d0_236[2:0] == 1) begin
        next_mux_d0_236 = input_word_d[1889];
    end else if (sel_d0_236[2:0] == 2) begin
        next_mux_d0_236 = input_word_d[1890];
    end else if (sel_d0_236[2:0] == 3) begin
        next_mux_d0_236 = input_word_d[1891];
    end else if (sel_d0_236[2:0] == 4) begin
        next_mux_d0_236 = input_word_d[1892];
    end else if (sel_d0_236[2:0] == 5) begin
        next_mux_d0_236 = input_word_d[1893];
    end else if (sel_d0_236[2:0] == 6) begin
        next_mux_d0_236 = input_word_d[1894];
    end else begin
        next_mux_d0_236 = input_word_d[1895];
    end

    if (sel_d0_237[2:0] == 0) begin
        next_mux_d0_237 = input_word_d[1896];
    end else if (sel_d0_237[2:0] == 1) begin
        next_mux_d0_237 = input_word_d[1897];
    end else if (sel_d0_237[2:0] == 2) begin
        next_mux_d0_237 = input_word_d[1898];
    end else if (sel_d0_237[2:0] == 3) begin
        next_mux_d0_237 = input_word_d[1899];
    end else if (sel_d0_237[2:0] == 4) begin
        next_mux_d0_237 = input_word_d[1900];
    end else if (sel_d0_237[2:0] == 5) begin
        next_mux_d0_237 = input_word_d[1901];
    end else if (sel_d0_237[2:0] == 6) begin
        next_mux_d0_237 = input_word_d[1902];
    end else begin
        next_mux_d0_237 = input_word_d[1903];
    end

    if (sel_d0_238[2:0] == 0) begin
        next_mux_d0_238 = input_word_d[1904];
    end else if (sel_d0_238[2:0] == 1) begin
        next_mux_d0_238 = input_word_d[1905];
    end else if (sel_d0_238[2:0] == 2) begin
        next_mux_d0_238 = input_word_d[1906];
    end else if (sel_d0_238[2:0] == 3) begin
        next_mux_d0_238 = input_word_d[1907];
    end else if (sel_d0_238[2:0] == 4) begin
        next_mux_d0_238 = input_word_d[1908];
    end else if (sel_d0_238[2:0] == 5) begin
        next_mux_d0_238 = input_word_d[1909];
    end else if (sel_d0_238[2:0] == 6) begin
        next_mux_d0_238 = input_word_d[1910];
    end else begin
        next_mux_d0_238 = input_word_d[1911];
    end

    if (sel_d0_239[2:0] == 0) begin
        next_mux_d0_239 = input_word_d[1912];
    end else if (sel_d0_239[2:0] == 1) begin
        next_mux_d0_239 = input_word_d[1913];
    end else if (sel_d0_239[2:0] == 2) begin
        next_mux_d0_239 = input_word_d[1914];
    end else if (sel_d0_239[2:0] == 3) begin
        next_mux_d0_239 = input_word_d[1915];
    end else if (sel_d0_239[2:0] == 4) begin
        next_mux_d0_239 = input_word_d[1916];
    end else if (sel_d0_239[2:0] == 5) begin
        next_mux_d0_239 = input_word_d[1917];
    end else if (sel_d0_239[2:0] == 6) begin
        next_mux_d0_239 = input_word_d[1918];
    end else begin
        next_mux_d0_239 = input_word_d[1919];
    end

    if (sel_d0_240[2:0] == 0) begin
        next_mux_d0_240 = input_word_d[1920];
    end else if (sel_d0_240[2:0] == 1) begin
        next_mux_d0_240 = input_word_d[1921];
    end else if (sel_d0_240[2:0] == 2) begin
        next_mux_d0_240 = input_word_d[1922];
    end else if (sel_d0_240[2:0] == 3) begin
        next_mux_d0_240 = input_word_d[1923];
    end else if (sel_d0_240[2:0] == 4) begin
        next_mux_d0_240 = input_word_d[1924];
    end else if (sel_d0_240[2:0] == 5) begin
        next_mux_d0_240 = input_word_d[1925];
    end else if (sel_d0_240[2:0] == 6) begin
        next_mux_d0_240 = input_word_d[1926];
    end else begin
        next_mux_d0_240 = input_word_d[1927];
    end

    if (sel_d0_241[2:0] == 0) begin
        next_mux_d0_241 = input_word_d[1928];
    end else if (sel_d0_241[2:0] == 1) begin
        next_mux_d0_241 = input_word_d[1929];
    end else if (sel_d0_241[2:0] == 2) begin
        next_mux_d0_241 = input_word_d[1930];
    end else if (sel_d0_241[2:0] == 3) begin
        next_mux_d0_241 = input_word_d[1931];
    end else if (sel_d0_241[2:0] == 4) begin
        next_mux_d0_241 = input_word_d[1932];
    end else if (sel_d0_241[2:0] == 5) begin
        next_mux_d0_241 = input_word_d[1933];
    end else if (sel_d0_241[2:0] == 6) begin
        next_mux_d0_241 = input_word_d[1934];
    end else begin
        next_mux_d0_241 = input_word_d[1935];
    end

    if (sel_d0_242[2:0] == 0) begin
        next_mux_d0_242 = input_word_d[1936];
    end else if (sel_d0_242[2:0] == 1) begin
        next_mux_d0_242 = input_word_d[1937];
    end else if (sel_d0_242[2:0] == 2) begin
        next_mux_d0_242 = input_word_d[1938];
    end else if (sel_d0_242[2:0] == 3) begin
        next_mux_d0_242 = input_word_d[1939];
    end else if (sel_d0_242[2:0] == 4) begin
        next_mux_d0_242 = input_word_d[1940];
    end else if (sel_d0_242[2:0] == 5) begin
        next_mux_d0_242 = input_word_d[1941];
    end else if (sel_d0_242[2:0] == 6) begin
        next_mux_d0_242 = input_word_d[1942];
    end else begin
        next_mux_d0_242 = input_word_d[1943];
    end

    if (sel_d0_243[2:0] == 0) begin
        next_mux_d0_243 = input_word_d[1944];
    end else if (sel_d0_243[2:0] == 1) begin
        next_mux_d0_243 = input_word_d[1945];
    end else if (sel_d0_243[2:0] == 2) begin
        next_mux_d0_243 = input_word_d[1946];
    end else if (sel_d0_243[2:0] == 3) begin
        next_mux_d0_243 = input_word_d[1947];
    end else if (sel_d0_243[2:0] == 4) begin
        next_mux_d0_243 = input_word_d[1948];
    end else if (sel_d0_243[2:0] == 5) begin
        next_mux_d0_243 = input_word_d[1949];
    end else if (sel_d0_243[2:0] == 6) begin
        next_mux_d0_243 = input_word_d[1950];
    end else begin
        next_mux_d0_243 = input_word_d[1951];
    end

    if (sel_d0_244[2:0] == 0) begin
        next_mux_d0_244 = input_word_d[1952];
    end else if (sel_d0_244[2:0] == 1) begin
        next_mux_d0_244 = input_word_d[1953];
    end else if (sel_d0_244[2:0] == 2) begin
        next_mux_d0_244 = input_word_d[1954];
    end else if (sel_d0_244[2:0] == 3) begin
        next_mux_d0_244 = input_word_d[1955];
    end else if (sel_d0_244[2:0] == 4) begin
        next_mux_d0_244 = input_word_d[1956];
    end else if (sel_d0_244[2:0] == 5) begin
        next_mux_d0_244 = input_word_d[1957];
    end else if (sel_d0_244[2:0] == 6) begin
        next_mux_d0_244 = input_word_d[1958];
    end else begin
        next_mux_d0_244 = input_word_d[1959];
    end

    if (sel_d0_245[2:0] == 0) begin
        next_mux_d0_245 = input_word_d[1960];
    end else if (sel_d0_245[2:0] == 1) begin
        next_mux_d0_245 = input_word_d[1961];
    end else if (sel_d0_245[2:0] == 2) begin
        next_mux_d0_245 = input_word_d[1962];
    end else if (sel_d0_245[2:0] == 3) begin
        next_mux_d0_245 = input_word_d[1963];
    end else if (sel_d0_245[2:0] == 4) begin
        next_mux_d0_245 = input_word_d[1964];
    end else if (sel_d0_245[2:0] == 5) begin
        next_mux_d0_245 = input_word_d[1965];
    end else if (sel_d0_245[2:0] == 6) begin
        next_mux_d0_245 = input_word_d[1966];
    end else begin
        next_mux_d0_245 = input_word_d[1967];
    end

    if (sel_d0_246[2:0] == 0) begin
        next_mux_d0_246 = input_word_d[1968];
    end else if (sel_d0_246[2:0] == 1) begin
        next_mux_d0_246 = input_word_d[1969];
    end else if (sel_d0_246[2:0] == 2) begin
        next_mux_d0_246 = input_word_d[1970];
    end else if (sel_d0_246[2:0] == 3) begin
        next_mux_d0_246 = input_word_d[1971];
    end else if (sel_d0_246[2:0] == 4) begin
        next_mux_d0_246 = input_word_d[1972];
    end else if (sel_d0_246[2:0] == 5) begin
        next_mux_d0_246 = input_word_d[1973];
    end else if (sel_d0_246[2:0] == 6) begin
        next_mux_d0_246 = input_word_d[1974];
    end else begin
        next_mux_d0_246 = input_word_d[1975];
    end

    if (sel_d0_247[2:0] == 0) begin
        next_mux_d0_247 = input_word_d[1976];
    end else if (sel_d0_247[2:0] == 1) begin
        next_mux_d0_247 = input_word_d[1977];
    end else if (sel_d0_247[2:0] == 2) begin
        next_mux_d0_247 = input_word_d[1978];
    end else if (sel_d0_247[2:0] == 3) begin
        next_mux_d0_247 = input_word_d[1979];
    end else if (sel_d0_247[2:0] == 4) begin
        next_mux_d0_247 = input_word_d[1980];
    end else if (sel_d0_247[2:0] == 5) begin
        next_mux_d0_247 = input_word_d[1981];
    end else if (sel_d0_247[2:0] == 6) begin
        next_mux_d0_247 = input_word_d[1982];
    end else begin
        next_mux_d0_247 = input_word_d[1983];
    end

    if (sel_d0_248[2:0] == 0) begin
        next_mux_d0_248 = input_word_d[1984];
    end else if (sel_d0_248[2:0] == 1) begin
        next_mux_d0_248 = input_word_d[1985];
    end else if (sel_d0_248[2:0] == 2) begin
        next_mux_d0_248 = input_word_d[1986];
    end else if (sel_d0_248[2:0] == 3) begin
        next_mux_d0_248 = input_word_d[1987];
    end else if (sel_d0_248[2:0] == 4) begin
        next_mux_d0_248 = input_word_d[1988];
    end else if (sel_d0_248[2:0] == 5) begin
        next_mux_d0_248 = input_word_d[1989];
    end else if (sel_d0_248[2:0] == 6) begin
        next_mux_d0_248 = input_word_d[1990];
    end else begin
        next_mux_d0_248 = input_word_d[1991];
    end

    if (sel_d0_249[2:0] == 0) begin
        next_mux_d0_249 = input_word_d[1992];
    end else if (sel_d0_249[2:0] == 1) begin
        next_mux_d0_249 = input_word_d[1993];
    end else if (sel_d0_249[2:0] == 2) begin
        next_mux_d0_249 = input_word_d[1994];
    end else if (sel_d0_249[2:0] == 3) begin
        next_mux_d0_249 = input_word_d[1995];
    end else if (sel_d0_249[2:0] == 4) begin
        next_mux_d0_249 = input_word_d[1996];
    end else if (sel_d0_249[2:0] == 5) begin
        next_mux_d0_249 = input_word_d[1997];
    end else if (sel_d0_249[2:0] == 6) begin
        next_mux_d0_249 = input_word_d[1998];
    end else begin
        next_mux_d0_249 = input_word_d[1999];
    end

    if (sel_d0_250[2:0] == 0) begin
        next_mux_d0_250 = input_word_d[2000];
    end else if (sel_d0_250[2:0] == 1) begin
        next_mux_d0_250 = input_word_d[2001];
    end else if (sel_d0_250[2:0] == 2) begin
        next_mux_d0_250 = input_word_d[2002];
    end else if (sel_d0_250[2:0] == 3) begin
        next_mux_d0_250 = input_word_d[2003];
    end else if (sel_d0_250[2:0] == 4) begin
        next_mux_d0_250 = input_word_d[2004];
    end else if (sel_d0_250[2:0] == 5) begin
        next_mux_d0_250 = input_word_d[2005];
    end else if (sel_d0_250[2:0] == 6) begin
        next_mux_d0_250 = input_word_d[2006];
    end else begin
        next_mux_d0_250 = input_word_d[2007];
    end

    if (sel_d0_251[2:0] == 0) begin
        next_mux_d0_251 = input_word_d[2008];
    end else if (sel_d0_251[2:0] == 1) begin
        next_mux_d0_251 = input_word_d[2009];
    end else if (sel_d0_251[2:0] == 2) begin
        next_mux_d0_251 = input_word_d[2010];
    end else if (sel_d0_251[2:0] == 3) begin
        next_mux_d0_251 = input_word_d[2011];
    end else if (sel_d0_251[2:0] == 4) begin
        next_mux_d0_251 = input_word_d[2012];
    end else if (sel_d0_251[2:0] == 5) begin
        next_mux_d0_251 = input_word_d[2013];
    end else if (sel_d0_251[2:0] == 6) begin
        next_mux_d0_251 = input_word_d[2014];
    end else begin
        next_mux_d0_251 = input_word_d[2015];
    end

    if (sel_d0_252[2:0] == 0) begin
        next_mux_d0_252 = input_word_d[2016];
    end else if (sel_d0_252[2:0] == 1) begin
        next_mux_d0_252 = input_word_d[2017];
    end else if (sel_d0_252[2:0] == 2) begin
        next_mux_d0_252 = input_word_d[2018];
    end else if (sel_d0_252[2:0] == 3) begin
        next_mux_d0_252 = input_word_d[2019];
    end else if (sel_d0_252[2:0] == 4) begin
        next_mux_d0_252 = input_word_d[2020];
    end else if (sel_d0_252[2:0] == 5) begin
        next_mux_d0_252 = input_word_d[2021];
    end else if (sel_d0_252[2:0] == 6) begin
        next_mux_d0_252 = input_word_d[2022];
    end else begin
        next_mux_d0_252 = input_word_d[2023];
    end

    if (sel_d0_253[2:0] == 0) begin
        next_mux_d0_253 = input_word_d[2024];
    end else if (sel_d0_253[2:0] == 1) begin
        next_mux_d0_253 = input_word_d[2025];
    end else if (sel_d0_253[2:0] == 2) begin
        next_mux_d0_253 = input_word_d[2026];
    end else if (sel_d0_253[2:0] == 3) begin
        next_mux_d0_253 = input_word_d[2027];
    end else if (sel_d0_253[2:0] == 4) begin
        next_mux_d0_253 = input_word_d[2028];
    end else if (sel_d0_253[2:0] == 5) begin
        next_mux_d0_253 = input_word_d[2029];
    end else if (sel_d0_253[2:0] == 6) begin
        next_mux_d0_253 = input_word_d[2030];
    end else begin
        next_mux_d0_253 = input_word_d[2031];
    end

    if (sel_d0_254[2:0] == 0) begin
        next_mux_d0_254 = input_word_d[2032];
    end else if (sel_d0_254[2:0] == 1) begin
        next_mux_d0_254 = input_word_d[2033];
    end else if (sel_d0_254[2:0] == 2) begin
        next_mux_d0_254 = input_word_d[2034];
    end else if (sel_d0_254[2:0] == 3) begin
        next_mux_d0_254 = input_word_d[2035];
    end else if (sel_d0_254[2:0] == 4) begin
        next_mux_d0_254 = input_word_d[2036];
    end else if (sel_d0_254[2:0] == 5) begin
        next_mux_d0_254 = input_word_d[2037];
    end else if (sel_d0_254[2:0] == 6) begin
        next_mux_d0_254 = input_word_d[2038];
    end else begin
        next_mux_d0_254 = input_word_d[2039];
    end

    if (sel_d0_255[2:0] == 0) begin
        next_mux_d0_255 = input_word_d[2040];
    end else if (sel_d0_255[2:0] == 1) begin
        next_mux_d0_255 = input_word_d[2041];
    end else if (sel_d0_255[2:0] == 2) begin
        next_mux_d0_255 = input_word_d[2042];
    end else if (sel_d0_255[2:0] == 3) begin
        next_mux_d0_255 = input_word_d[2043];
    end else if (sel_d0_255[2:0] == 4) begin
        next_mux_d0_255 = input_word_d[2044];
    end else if (sel_d0_255[2:0] == 5) begin
        next_mux_d0_255 = input_word_d[2045];
    end else if (sel_d0_255[2:0] == 6) begin
        next_mux_d0_255 = input_word_d[2046];
    end else begin
        next_mux_d0_255 = input_word_d[2047];
    end

    if (sel_d1_0[5:3] == 0) begin
        next_mux_d1_0 = mux_d0_0;
    end else if (sel_d1_0[5:3] == 1) begin
        next_mux_d1_0 = mux_d0_1;
    end else if (sel_d1_0[5:3] == 2) begin
        next_mux_d1_0 = mux_d0_2;
    end else if (sel_d1_0[5:3] == 3) begin
        next_mux_d1_0 = mux_d0_3;
    end else if (sel_d1_0[5:3] == 4) begin
        next_mux_d1_0 = mux_d0_4;
    end else if (sel_d1_0[5:3] == 5) begin
        next_mux_d1_0 = mux_d0_5;
    end else if (sel_d1_0[5:3] == 6) begin
        next_mux_d1_0 = mux_d0_6;
    end else begin
        next_mux_d1_0 = mux_d0_7;
    end

    if (sel_d1_1[5:3] == 0) begin
        next_mux_d1_1 = mux_d0_0;
    end else if (sel_d1_1[5:3] == 1) begin
        next_mux_d1_1 = mux_d0_1;
    end else if (sel_d1_1[5:3] == 2) begin
        next_mux_d1_1 = mux_d0_2;
    end else if (sel_d1_1[5:3] == 3) begin
        next_mux_d1_1 = mux_d0_3;
    end else if (sel_d1_1[5:3] == 4) begin
        next_mux_d1_1 = mux_d0_4;
    end else if (sel_d1_1[5:3] == 5) begin
        next_mux_d1_1 = mux_d0_5;
    end else if (sel_d1_1[5:3] == 6) begin
        next_mux_d1_1 = mux_d0_6;
    end else begin
        next_mux_d1_1 = mux_d0_7;
    end

    if (sel_d1_2[5:3] == 0) begin
        next_mux_d1_2 = mux_d0_0;
    end else if (sel_d1_2[5:3] == 1) begin
        next_mux_d1_2 = mux_d0_1;
    end else if (sel_d1_2[5:3] == 2) begin
        next_mux_d1_2 = mux_d0_2;
    end else if (sel_d1_2[5:3] == 3) begin
        next_mux_d1_2 = mux_d0_3;
    end else if (sel_d1_2[5:3] == 4) begin
        next_mux_d1_2 = mux_d0_4;
    end else if (sel_d1_2[5:3] == 5) begin
        next_mux_d1_2 = mux_d0_5;
    end else if (sel_d1_2[5:3] == 6) begin
        next_mux_d1_2 = mux_d0_6;
    end else begin
        next_mux_d1_2 = mux_d0_7;
    end

    if (sel_d1_3[5:3] == 0) begin
        next_mux_d1_3 = mux_d0_0;
    end else if (sel_d1_3[5:3] == 1) begin
        next_mux_d1_3 = mux_d0_1;
    end else if (sel_d1_3[5:3] == 2) begin
        next_mux_d1_3 = mux_d0_2;
    end else if (sel_d1_3[5:3] == 3) begin
        next_mux_d1_3 = mux_d0_3;
    end else if (sel_d1_3[5:3] == 4) begin
        next_mux_d1_3 = mux_d0_4;
    end else if (sel_d1_3[5:3] == 5) begin
        next_mux_d1_3 = mux_d0_5;
    end else if (sel_d1_3[5:3] == 6) begin
        next_mux_d1_3 = mux_d0_6;
    end else begin
        next_mux_d1_3 = mux_d0_7;
    end

    if (sel_d1_4[5:3] == 0) begin
        next_mux_d1_4 = mux_d0_0;
    end else if (sel_d1_4[5:3] == 1) begin
        next_mux_d1_4 = mux_d0_1;
    end else if (sel_d1_4[5:3] == 2) begin
        next_mux_d1_4 = mux_d0_2;
    end else if (sel_d1_4[5:3] == 3) begin
        next_mux_d1_4 = mux_d0_3;
    end else if (sel_d1_4[5:3] == 4) begin
        next_mux_d1_4 = mux_d0_4;
    end else if (sel_d1_4[5:3] == 5) begin
        next_mux_d1_4 = mux_d0_5;
    end else if (sel_d1_4[5:3] == 6) begin
        next_mux_d1_4 = mux_d0_6;
    end else begin
        next_mux_d1_4 = mux_d0_7;
    end

    if (sel_d1_5[5:3] == 0) begin
        next_mux_d1_5 = mux_d0_0;
    end else if (sel_d1_5[5:3] == 1) begin
        next_mux_d1_5 = mux_d0_1;
    end else if (sel_d1_5[5:3] == 2) begin
        next_mux_d1_5 = mux_d0_2;
    end else if (sel_d1_5[5:3] == 3) begin
        next_mux_d1_5 = mux_d0_3;
    end else if (sel_d1_5[5:3] == 4) begin
        next_mux_d1_5 = mux_d0_4;
    end else if (sel_d1_5[5:3] == 5) begin
        next_mux_d1_5 = mux_d0_5;
    end else if (sel_d1_5[5:3] == 6) begin
        next_mux_d1_5 = mux_d0_6;
    end else begin
        next_mux_d1_5 = mux_d0_7;
    end

    if (sel_d1_6[5:3] == 0) begin
        next_mux_d1_6 = mux_d0_0;
    end else if (sel_d1_6[5:3] == 1) begin
        next_mux_d1_6 = mux_d0_1;
    end else if (sel_d1_6[5:3] == 2) begin
        next_mux_d1_6 = mux_d0_2;
    end else if (sel_d1_6[5:3] == 3) begin
        next_mux_d1_6 = mux_d0_3;
    end else if (sel_d1_6[5:3] == 4) begin
        next_mux_d1_6 = mux_d0_4;
    end else if (sel_d1_6[5:3] == 5) begin
        next_mux_d1_6 = mux_d0_5;
    end else if (sel_d1_6[5:3] == 6) begin
        next_mux_d1_6 = mux_d0_6;
    end else begin
        next_mux_d1_6 = mux_d0_7;
    end

    if (sel_d1_7[5:3] == 0) begin
        next_mux_d1_7 = mux_d0_0;
    end else if (sel_d1_7[5:3] == 1) begin
        next_mux_d1_7 = mux_d0_1;
    end else if (sel_d1_7[5:3] == 2) begin
        next_mux_d1_7 = mux_d0_2;
    end else if (sel_d1_7[5:3] == 3) begin
        next_mux_d1_7 = mux_d0_3;
    end else if (sel_d1_7[5:3] == 4) begin
        next_mux_d1_7 = mux_d0_4;
    end else if (sel_d1_7[5:3] == 5) begin
        next_mux_d1_7 = mux_d0_5;
    end else if (sel_d1_7[5:3] == 6) begin
        next_mux_d1_7 = mux_d0_6;
    end else begin
        next_mux_d1_7 = mux_d0_7;
    end

    if (sel_d1_8[5:3] == 0) begin
        next_mux_d1_8 = mux_d0_0;
    end else if (sel_d1_8[5:3] == 1) begin
        next_mux_d1_8 = mux_d0_1;
    end else if (sel_d1_8[5:3] == 2) begin
        next_mux_d1_8 = mux_d0_2;
    end else if (sel_d1_8[5:3] == 3) begin
        next_mux_d1_8 = mux_d0_3;
    end else if (sel_d1_8[5:3] == 4) begin
        next_mux_d1_8 = mux_d0_4;
    end else if (sel_d1_8[5:3] == 5) begin
        next_mux_d1_8 = mux_d0_5;
    end else if (sel_d1_8[5:3] == 6) begin
        next_mux_d1_8 = mux_d0_6;
    end else begin
        next_mux_d1_8 = mux_d0_7;
    end

    if (sel_d1_9[5:3] == 0) begin
        next_mux_d1_9 = mux_d0_0;
    end else if (sel_d1_9[5:3] == 1) begin
        next_mux_d1_9 = mux_d0_1;
    end else if (sel_d1_9[5:3] == 2) begin
        next_mux_d1_9 = mux_d0_2;
    end else if (sel_d1_9[5:3] == 3) begin
        next_mux_d1_9 = mux_d0_3;
    end else if (sel_d1_9[5:3] == 4) begin
        next_mux_d1_9 = mux_d0_4;
    end else if (sel_d1_9[5:3] == 5) begin
        next_mux_d1_9 = mux_d0_5;
    end else if (sel_d1_9[5:3] == 6) begin
        next_mux_d1_9 = mux_d0_6;
    end else begin
        next_mux_d1_9 = mux_d0_7;
    end

    if (sel_d1_10[5:3] == 0) begin
        next_mux_d1_10 = mux_d0_0;
    end else if (sel_d1_10[5:3] == 1) begin
        next_mux_d1_10 = mux_d0_1;
    end else if (sel_d1_10[5:3] == 2) begin
        next_mux_d1_10 = mux_d0_2;
    end else if (sel_d1_10[5:3] == 3) begin
        next_mux_d1_10 = mux_d0_3;
    end else if (sel_d1_10[5:3] == 4) begin
        next_mux_d1_10 = mux_d0_4;
    end else if (sel_d1_10[5:3] == 5) begin
        next_mux_d1_10 = mux_d0_5;
    end else if (sel_d1_10[5:3] == 6) begin
        next_mux_d1_10 = mux_d0_6;
    end else begin
        next_mux_d1_10 = mux_d0_7;
    end

    if (sel_d1_11[5:3] == 0) begin
        next_mux_d1_11 = mux_d0_0;
    end else if (sel_d1_11[5:3] == 1) begin
        next_mux_d1_11 = mux_d0_1;
    end else if (sel_d1_11[5:3] == 2) begin
        next_mux_d1_11 = mux_d0_2;
    end else if (sel_d1_11[5:3] == 3) begin
        next_mux_d1_11 = mux_d0_3;
    end else if (sel_d1_11[5:3] == 4) begin
        next_mux_d1_11 = mux_d0_4;
    end else if (sel_d1_11[5:3] == 5) begin
        next_mux_d1_11 = mux_d0_5;
    end else if (sel_d1_11[5:3] == 6) begin
        next_mux_d1_11 = mux_d0_6;
    end else begin
        next_mux_d1_11 = mux_d0_7;
    end

    if (sel_d1_12[5:3] == 0) begin
        next_mux_d1_12 = mux_d0_0;
    end else if (sel_d1_12[5:3] == 1) begin
        next_mux_d1_12 = mux_d0_1;
    end else if (sel_d1_12[5:3] == 2) begin
        next_mux_d1_12 = mux_d0_2;
    end else if (sel_d1_12[5:3] == 3) begin
        next_mux_d1_12 = mux_d0_3;
    end else if (sel_d1_12[5:3] == 4) begin
        next_mux_d1_12 = mux_d0_4;
    end else if (sel_d1_12[5:3] == 5) begin
        next_mux_d1_12 = mux_d0_5;
    end else if (sel_d1_12[5:3] == 6) begin
        next_mux_d1_12 = mux_d0_6;
    end else begin
        next_mux_d1_12 = mux_d0_7;
    end

    if (sel_d1_13[5:3] == 0) begin
        next_mux_d1_13 = mux_d0_0;
    end else if (sel_d1_13[5:3] == 1) begin
        next_mux_d1_13 = mux_d0_1;
    end else if (sel_d1_13[5:3] == 2) begin
        next_mux_d1_13 = mux_d0_2;
    end else if (sel_d1_13[5:3] == 3) begin
        next_mux_d1_13 = mux_d0_3;
    end else if (sel_d1_13[5:3] == 4) begin
        next_mux_d1_13 = mux_d0_4;
    end else if (sel_d1_13[5:3] == 5) begin
        next_mux_d1_13 = mux_d0_5;
    end else if (sel_d1_13[5:3] == 6) begin
        next_mux_d1_13 = mux_d0_6;
    end else begin
        next_mux_d1_13 = mux_d0_7;
    end

    if (sel_d1_14[5:3] == 0) begin
        next_mux_d1_14 = mux_d0_0;
    end else if (sel_d1_14[5:3] == 1) begin
        next_mux_d1_14 = mux_d0_1;
    end else if (sel_d1_14[5:3] == 2) begin
        next_mux_d1_14 = mux_d0_2;
    end else if (sel_d1_14[5:3] == 3) begin
        next_mux_d1_14 = mux_d0_3;
    end else if (sel_d1_14[5:3] == 4) begin
        next_mux_d1_14 = mux_d0_4;
    end else if (sel_d1_14[5:3] == 5) begin
        next_mux_d1_14 = mux_d0_5;
    end else if (sel_d1_14[5:3] == 6) begin
        next_mux_d1_14 = mux_d0_6;
    end else begin
        next_mux_d1_14 = mux_d0_7;
    end

    if (sel_d1_15[5:3] == 0) begin
        next_mux_d1_15 = mux_d0_0;
    end else if (sel_d1_15[5:3] == 1) begin
        next_mux_d1_15 = mux_d0_1;
    end else if (sel_d1_15[5:3] == 2) begin
        next_mux_d1_15 = mux_d0_2;
    end else if (sel_d1_15[5:3] == 3) begin
        next_mux_d1_15 = mux_d0_3;
    end else if (sel_d1_15[5:3] == 4) begin
        next_mux_d1_15 = mux_d0_4;
    end else if (sel_d1_15[5:3] == 5) begin
        next_mux_d1_15 = mux_d0_5;
    end else if (sel_d1_15[5:3] == 6) begin
        next_mux_d1_15 = mux_d0_6;
    end else begin
        next_mux_d1_15 = mux_d0_7;
    end

    if (sel_d1_16[5:3] == 0) begin
        next_mux_d1_16 = mux_d0_0;
    end else if (sel_d1_16[5:3] == 1) begin
        next_mux_d1_16 = mux_d0_1;
    end else if (sel_d1_16[5:3] == 2) begin
        next_mux_d1_16 = mux_d0_2;
    end else if (sel_d1_16[5:3] == 3) begin
        next_mux_d1_16 = mux_d0_3;
    end else if (sel_d1_16[5:3] == 4) begin
        next_mux_d1_16 = mux_d0_4;
    end else if (sel_d1_16[5:3] == 5) begin
        next_mux_d1_16 = mux_d0_5;
    end else if (sel_d1_16[5:3] == 6) begin
        next_mux_d1_16 = mux_d0_6;
    end else begin
        next_mux_d1_16 = mux_d0_7;
    end

    if (sel_d1_17[5:3] == 0) begin
        next_mux_d1_17 = mux_d0_0;
    end else if (sel_d1_17[5:3] == 1) begin
        next_mux_d1_17 = mux_d0_1;
    end else if (sel_d1_17[5:3] == 2) begin
        next_mux_d1_17 = mux_d0_2;
    end else if (sel_d1_17[5:3] == 3) begin
        next_mux_d1_17 = mux_d0_3;
    end else if (sel_d1_17[5:3] == 4) begin
        next_mux_d1_17 = mux_d0_4;
    end else if (sel_d1_17[5:3] == 5) begin
        next_mux_d1_17 = mux_d0_5;
    end else if (sel_d1_17[5:3] == 6) begin
        next_mux_d1_17 = mux_d0_6;
    end else begin
        next_mux_d1_17 = mux_d0_7;
    end

    if (sel_d1_18[5:3] == 0) begin
        next_mux_d1_18 = mux_d0_0;
    end else if (sel_d1_18[5:3] == 1) begin
        next_mux_d1_18 = mux_d0_1;
    end else if (sel_d1_18[5:3] == 2) begin
        next_mux_d1_18 = mux_d0_2;
    end else if (sel_d1_18[5:3] == 3) begin
        next_mux_d1_18 = mux_d0_3;
    end else if (sel_d1_18[5:3] == 4) begin
        next_mux_d1_18 = mux_d0_4;
    end else if (sel_d1_18[5:3] == 5) begin
        next_mux_d1_18 = mux_d0_5;
    end else if (sel_d1_18[5:3] == 6) begin
        next_mux_d1_18 = mux_d0_6;
    end else begin
        next_mux_d1_18 = mux_d0_7;
    end

    if (sel_d1_19[5:3] == 0) begin
        next_mux_d1_19 = mux_d0_0;
    end else if (sel_d1_19[5:3] == 1) begin
        next_mux_d1_19 = mux_d0_1;
    end else if (sel_d1_19[5:3] == 2) begin
        next_mux_d1_19 = mux_d0_2;
    end else if (sel_d1_19[5:3] == 3) begin
        next_mux_d1_19 = mux_d0_3;
    end else if (sel_d1_19[5:3] == 4) begin
        next_mux_d1_19 = mux_d0_4;
    end else if (sel_d1_19[5:3] == 5) begin
        next_mux_d1_19 = mux_d0_5;
    end else if (sel_d1_19[5:3] == 6) begin
        next_mux_d1_19 = mux_d0_6;
    end else begin
        next_mux_d1_19 = mux_d0_7;
    end

    if (sel_d1_20[5:3] == 0) begin
        next_mux_d1_20 = mux_d0_0;
    end else if (sel_d1_20[5:3] == 1) begin
        next_mux_d1_20 = mux_d0_1;
    end else if (sel_d1_20[5:3] == 2) begin
        next_mux_d1_20 = mux_d0_2;
    end else if (sel_d1_20[5:3] == 3) begin
        next_mux_d1_20 = mux_d0_3;
    end else if (sel_d1_20[5:3] == 4) begin
        next_mux_d1_20 = mux_d0_4;
    end else if (sel_d1_20[5:3] == 5) begin
        next_mux_d1_20 = mux_d0_5;
    end else if (sel_d1_20[5:3] == 6) begin
        next_mux_d1_20 = mux_d0_6;
    end else begin
        next_mux_d1_20 = mux_d0_7;
    end

    if (sel_d1_21[5:3] == 0) begin
        next_mux_d1_21 = mux_d0_0;
    end else if (sel_d1_21[5:3] == 1) begin
        next_mux_d1_21 = mux_d0_1;
    end else if (sel_d1_21[5:3] == 2) begin
        next_mux_d1_21 = mux_d0_2;
    end else if (sel_d1_21[5:3] == 3) begin
        next_mux_d1_21 = mux_d0_3;
    end else if (sel_d1_21[5:3] == 4) begin
        next_mux_d1_21 = mux_d0_4;
    end else if (sel_d1_21[5:3] == 5) begin
        next_mux_d1_21 = mux_d0_5;
    end else if (sel_d1_21[5:3] == 6) begin
        next_mux_d1_21 = mux_d0_6;
    end else begin
        next_mux_d1_21 = mux_d0_7;
    end

    if (sel_d1_22[5:3] == 0) begin
        next_mux_d1_22 = mux_d0_0;
    end else if (sel_d1_22[5:3] == 1) begin
        next_mux_d1_22 = mux_d0_1;
    end else if (sel_d1_22[5:3] == 2) begin
        next_mux_d1_22 = mux_d0_2;
    end else if (sel_d1_22[5:3] == 3) begin
        next_mux_d1_22 = mux_d0_3;
    end else if (sel_d1_22[5:3] == 4) begin
        next_mux_d1_22 = mux_d0_4;
    end else if (sel_d1_22[5:3] == 5) begin
        next_mux_d1_22 = mux_d0_5;
    end else if (sel_d1_22[5:3] == 6) begin
        next_mux_d1_22 = mux_d0_6;
    end else begin
        next_mux_d1_22 = mux_d0_7;
    end

    if (sel_d1_23[5:3] == 0) begin
        next_mux_d1_23 = mux_d0_0;
    end else if (sel_d1_23[5:3] == 1) begin
        next_mux_d1_23 = mux_d0_1;
    end else if (sel_d1_23[5:3] == 2) begin
        next_mux_d1_23 = mux_d0_2;
    end else if (sel_d1_23[5:3] == 3) begin
        next_mux_d1_23 = mux_d0_3;
    end else if (sel_d1_23[5:3] == 4) begin
        next_mux_d1_23 = mux_d0_4;
    end else if (sel_d1_23[5:3] == 5) begin
        next_mux_d1_23 = mux_d0_5;
    end else if (sel_d1_23[5:3] == 6) begin
        next_mux_d1_23 = mux_d0_6;
    end else begin
        next_mux_d1_23 = mux_d0_7;
    end

    if (sel_d1_24[5:3] == 0) begin
        next_mux_d1_24 = mux_d0_0;
    end else if (sel_d1_24[5:3] == 1) begin
        next_mux_d1_24 = mux_d0_1;
    end else if (sel_d1_24[5:3] == 2) begin
        next_mux_d1_24 = mux_d0_2;
    end else if (sel_d1_24[5:3] == 3) begin
        next_mux_d1_24 = mux_d0_3;
    end else if (sel_d1_24[5:3] == 4) begin
        next_mux_d1_24 = mux_d0_4;
    end else if (sel_d1_24[5:3] == 5) begin
        next_mux_d1_24 = mux_d0_5;
    end else if (sel_d1_24[5:3] == 6) begin
        next_mux_d1_24 = mux_d0_6;
    end else begin
        next_mux_d1_24 = mux_d0_7;
    end

    if (sel_d1_25[5:3] == 0) begin
        next_mux_d1_25 = mux_d0_0;
    end else if (sel_d1_25[5:3] == 1) begin
        next_mux_d1_25 = mux_d0_1;
    end else if (sel_d1_25[5:3] == 2) begin
        next_mux_d1_25 = mux_d0_2;
    end else if (sel_d1_25[5:3] == 3) begin
        next_mux_d1_25 = mux_d0_3;
    end else if (sel_d1_25[5:3] == 4) begin
        next_mux_d1_25 = mux_d0_4;
    end else if (sel_d1_25[5:3] == 5) begin
        next_mux_d1_25 = mux_d0_5;
    end else if (sel_d1_25[5:3] == 6) begin
        next_mux_d1_25 = mux_d0_6;
    end else begin
        next_mux_d1_25 = mux_d0_7;
    end

    if (sel_d1_26[5:3] == 0) begin
        next_mux_d1_26 = mux_d0_0;
    end else if (sel_d1_26[5:3] == 1) begin
        next_mux_d1_26 = mux_d0_1;
    end else if (sel_d1_26[5:3] == 2) begin
        next_mux_d1_26 = mux_d0_2;
    end else if (sel_d1_26[5:3] == 3) begin
        next_mux_d1_26 = mux_d0_3;
    end else if (sel_d1_26[5:3] == 4) begin
        next_mux_d1_26 = mux_d0_4;
    end else if (sel_d1_26[5:3] == 5) begin
        next_mux_d1_26 = mux_d0_5;
    end else if (sel_d1_26[5:3] == 6) begin
        next_mux_d1_26 = mux_d0_6;
    end else begin
        next_mux_d1_26 = mux_d0_7;
    end

    if (sel_d1_27[5:3] == 0) begin
        next_mux_d1_27 = mux_d0_0;
    end else if (sel_d1_27[5:3] == 1) begin
        next_mux_d1_27 = mux_d0_1;
    end else if (sel_d1_27[5:3] == 2) begin
        next_mux_d1_27 = mux_d0_2;
    end else if (sel_d1_27[5:3] == 3) begin
        next_mux_d1_27 = mux_d0_3;
    end else if (sel_d1_27[5:3] == 4) begin
        next_mux_d1_27 = mux_d0_4;
    end else if (sel_d1_27[5:3] == 5) begin
        next_mux_d1_27 = mux_d0_5;
    end else if (sel_d1_27[5:3] == 6) begin
        next_mux_d1_27 = mux_d0_6;
    end else begin
        next_mux_d1_27 = mux_d0_7;
    end

    if (sel_d1_28[5:3] == 0) begin
        next_mux_d1_28 = mux_d0_0;
    end else if (sel_d1_28[5:3] == 1) begin
        next_mux_d1_28 = mux_d0_1;
    end else if (sel_d1_28[5:3] == 2) begin
        next_mux_d1_28 = mux_d0_2;
    end else if (sel_d1_28[5:3] == 3) begin
        next_mux_d1_28 = mux_d0_3;
    end else if (sel_d1_28[5:3] == 4) begin
        next_mux_d1_28 = mux_d0_4;
    end else if (sel_d1_28[5:3] == 5) begin
        next_mux_d1_28 = mux_d0_5;
    end else if (sel_d1_28[5:3] == 6) begin
        next_mux_d1_28 = mux_d0_6;
    end else begin
        next_mux_d1_28 = mux_d0_7;
    end

    if (sel_d1_29[5:3] == 0) begin
        next_mux_d1_29 = mux_d0_0;
    end else if (sel_d1_29[5:3] == 1) begin
        next_mux_d1_29 = mux_d0_1;
    end else if (sel_d1_29[5:3] == 2) begin
        next_mux_d1_29 = mux_d0_2;
    end else if (sel_d1_29[5:3] == 3) begin
        next_mux_d1_29 = mux_d0_3;
    end else if (sel_d1_29[5:3] == 4) begin
        next_mux_d1_29 = mux_d0_4;
    end else if (sel_d1_29[5:3] == 5) begin
        next_mux_d1_29 = mux_d0_5;
    end else if (sel_d1_29[5:3] == 6) begin
        next_mux_d1_29 = mux_d0_6;
    end else begin
        next_mux_d1_29 = mux_d0_7;
    end

    if (sel_d1_30[5:3] == 0) begin
        next_mux_d1_30 = mux_d0_0;
    end else if (sel_d1_30[5:3] == 1) begin
        next_mux_d1_30 = mux_d0_1;
    end else if (sel_d1_30[5:3] == 2) begin
        next_mux_d1_30 = mux_d0_2;
    end else if (sel_d1_30[5:3] == 3) begin
        next_mux_d1_30 = mux_d0_3;
    end else if (sel_d1_30[5:3] == 4) begin
        next_mux_d1_30 = mux_d0_4;
    end else if (sel_d1_30[5:3] == 5) begin
        next_mux_d1_30 = mux_d0_5;
    end else if (sel_d1_30[5:3] == 6) begin
        next_mux_d1_30 = mux_d0_6;
    end else begin
        next_mux_d1_30 = mux_d0_7;
    end

    if (sel_d1_31[5:3] == 0) begin
        next_mux_d1_31 = mux_d0_0;
    end else if (sel_d1_31[5:3] == 1) begin
        next_mux_d1_31 = mux_d0_1;
    end else if (sel_d1_31[5:3] == 2) begin
        next_mux_d1_31 = mux_d0_2;
    end else if (sel_d1_31[5:3] == 3) begin
        next_mux_d1_31 = mux_d0_3;
    end else if (sel_d1_31[5:3] == 4) begin
        next_mux_d1_31 = mux_d0_4;
    end else if (sel_d1_31[5:3] == 5) begin
        next_mux_d1_31 = mux_d0_5;
    end else if (sel_d1_31[5:3] == 6) begin
        next_mux_d1_31 = mux_d0_6;
    end else begin
        next_mux_d1_31 = mux_d0_7;
    end

    if (sel_d2_0[8:6] == 0) begin
        next_mux_d2_0 = mux_d1_0;
    end else if (sel_d2_0[8:6] == 1) begin
        next_mux_d2_0 = mux_d1_1;
    end else if (sel_d2_0[8:6] == 2) begin
        next_mux_d2_0 = mux_d1_2;
    end else if (sel_d2_0[8:6] == 3) begin
        next_mux_d2_0 = mux_d1_3;
    end else if (sel_d2_0[8:6] == 4) begin
        next_mux_d2_0 = mux_d1_4;
    end else if (sel_d2_0[8:6] == 5) begin
        next_mux_d2_0 = mux_d1_5;
    end else if (sel_d2_0[8:6] == 6) begin
        next_mux_d2_0 = mux_d1_6;
    end else begin
        next_mux_d2_0 = mux_d1_7;
    end

    if (sel_d2_1[8:6] == 0) begin
        next_mux_d2_1 = mux_d1_0;
    end else if (sel_d2_1[8:6] == 1) begin
        next_mux_d2_1 = mux_d1_1;
    end else if (sel_d2_1[8:6] == 2) begin
        next_mux_d2_1 = mux_d1_2;
    end else if (sel_d2_1[8:6] == 3) begin
        next_mux_d2_1 = mux_d1_3;
    end else if (sel_d2_1[8:6] == 4) begin
        next_mux_d2_1 = mux_d1_4;
    end else if (sel_d2_1[8:6] == 5) begin
        next_mux_d2_1 = mux_d1_5;
    end else if (sel_d2_1[8:6] == 6) begin
        next_mux_d2_1 = mux_d1_6;
    end else begin
        next_mux_d2_1 = mux_d1_7;
    end

    if (sel_d2_2[8:6] == 0) begin
        next_mux_d2_2 = mux_d1_0;
    end else if (sel_d2_2[8:6] == 1) begin
        next_mux_d2_2 = mux_d1_1;
    end else if (sel_d2_2[8:6] == 2) begin
        next_mux_d2_2 = mux_d1_2;
    end else if (sel_d2_2[8:6] == 3) begin
        next_mux_d2_2 = mux_d1_3;
    end else if (sel_d2_2[8:6] == 4) begin
        next_mux_d2_2 = mux_d1_4;
    end else if (sel_d2_2[8:6] == 5) begin
        next_mux_d2_2 = mux_d1_5;
    end else if (sel_d2_2[8:6] == 6) begin
        next_mux_d2_2 = mux_d1_6;
    end else begin
        next_mux_d2_2 = mux_d1_7;
    end

    if (sel_d2_3[8:6] == 0) begin
        next_mux_d2_3 = mux_d1_0;
    end else if (sel_d2_3[8:6] == 1) begin
        next_mux_d2_3 = mux_d1_1;
    end else if (sel_d2_3[8:6] == 2) begin
        next_mux_d2_3 = mux_d1_2;
    end else if (sel_d2_3[8:6] == 3) begin
        next_mux_d2_3 = mux_d1_3;
    end else if (sel_d2_3[8:6] == 4) begin
        next_mux_d2_3 = mux_d1_4;
    end else if (sel_d2_3[8:6] == 5) begin
        next_mux_d2_3 = mux_d1_5;
    end else if (sel_d2_3[8:6] == 6) begin
        next_mux_d2_3 = mux_d1_6;
    end else begin
        next_mux_d2_3 = mux_d1_7;
    end

    if (sel_d3_0[10:9] == 0) begin
        next_mux_d3_0 = mux_d2_0;
    end else if (sel_d3_0[10:9] == 1) begin
        next_mux_d3_0 = mux_d2_1;
    end else if (sel_d3_0[10:9] == 2) begin
        next_mux_d3_0 = mux_d2_2;
    end else begin
        next_mux_d3_0 = mux_d2_3;
    end

end

endmodule
