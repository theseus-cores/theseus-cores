
/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : pfb_512Mmax_16iw_16ow_32tps_dp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data                                                     
//
//
/*****************************************************************************/


module pfb_512Mmax_16iw_16ow_32tps_dp_rom
(
  input clk, 
  input wea,
  input [13:0] addra,
  input [13:0] addrb,
  input [24:0] dia,
  output [24:0] dob
);

(* rom_style = "block" *) reg [24:0] rom [16383:0];
reg [13:0] addra_d;
reg [13:0] addrb_d;
reg [24:0] dob_d;
reg [24:0] rom_pipea;
reg [24:0] dia_d;
reg wea_d;

assign dob = dob_d;

initial
begin
    rom[0] = 25'b1111111111111111111111111;
    rom[1] = 25'b1111111111111111111111111;
    rom[2] = 25'b1111111111111111111111111;
    rom[3] = 25'b1111111111111111111111111;
    rom[4] = 25'b1111111111111111111111111;
    rom[5] = 25'b1111111111111111111111111;
    rom[6] = 25'b1111111111111111111111111;
    rom[7] = 25'b1111111111111111111111111;
    rom[8] = 25'b1111111111111111111111111;
    rom[9] = 25'b1111111111111111111111111;
    rom[10] = 25'b1111111111111111111111111;
    rom[11] = 25'b1111111111111111111111111;
    rom[12] = 25'b1111111111111111111111111;
    rom[13] = 25'b1111111111111111111111111;
    rom[14] = 25'b1111111111111111111111111;
    rom[15] = 25'b1111111111111111111111111;
    rom[16] = 25'b1111111111111111111111111;
    rom[17] = 25'b1111111111111111111111111;
    rom[18] = 25'b1111111111111111111111111;
    rom[19] = 25'b1111111111111111111111111;
    rom[20] = 25'b1111111111111111111111111;
    rom[21] = 25'b1111111111111111111111111;
    rom[22] = 25'b1111111111111111111111111;
    rom[23] = 25'b1111111111111111111111111;
    rom[24] = 25'b1111111111111111111111111;
    rom[25] = 25'b1111111111111111111111111;
    rom[26] = 25'b1111111111111111111111111;
    rom[27] = 25'b1111111111111111111111111;
    rom[28] = 25'b1111111111111111111111111;
    rom[29] = 25'b1111111111111111111111111;
    rom[30] = 25'b1111111111111111111111111;
    rom[31] = 25'b1111111111111111111111111;
    rom[32] = 25'b1111111111111111111111111;
    rom[33] = 25'b1111111111111111111111111;
    rom[34] = 25'b1111111111111111111111111;
    rom[35] = 25'b1111111111111111111111111;
    rom[36] = 25'b1111111111111111111111111;
    rom[37] = 25'b1111111111111111111111111;
    rom[38] = 25'b1111111111111111111111111;
    rom[39] = 25'b1111111111111111111111111;
    rom[40] = 25'b1111111111111111111111111;
    rom[41] = 25'b1111111111111111111111111;
    rom[42] = 25'b1111111111111111111111111;
    rom[43] = 25'b1111111111111111111111111;
    rom[44] = 25'b1111111111111111111111111;
    rom[45] = 25'b1111111111111111111111111;
    rom[46] = 25'b1111111111111111111111111;
    rom[47] = 25'b1111111111111111111111111;
    rom[48] = 25'b1111111111111111111111111;
    rom[49] = 25'b1111111111111111111111111;
    rom[50] = 25'b1111111111111111111111111;
    rom[51] = 25'b1111111111111111111111111;
    rom[52] = 25'b1111111111111111111111111;
    rom[53] = 25'b1111111111111111111111111;
    rom[54] = 25'b1111111111111111111111111;
    rom[55] = 25'b1111111111111111111111111;
    rom[56] = 25'b1111111111111111111111111;
    rom[57] = 25'b1111111111111111111111111;
    rom[58] = 25'b1111111111111111111111111;
    rom[59] = 25'b1111111111111111111111111;
    rom[60] = 25'b1111111111111111111111111;
    rom[61] = 25'b1111111111111111111111111;
    rom[62] = 25'b1111111111111111111111111;
    rom[63] = 25'b1111111111111111111111111;
    rom[64] = 25'b1111111111111111111111111;
    rom[65] = 25'b1111111111111111111111111;
    rom[66] = 25'b1111111111111111111111111;
    rom[67] = 25'b1111111111111111111111111;
    rom[68] = 25'b1111111111111111111111111;
    rom[69] = 25'b1111111111111111111111111;
    rom[70] = 25'b1111111111111111111111111;
    rom[71] = 25'b1111111111111111111111111;
    rom[72] = 25'b1111111111111111111111111;
    rom[73] = 25'b1111111111111111111111111;
    rom[74] = 25'b1111111111111111111111111;
    rom[75] = 25'b1111111111111111111111111;
    rom[76] = 25'b1111111111111111111111111;
    rom[77] = 25'b1111111111111111111111111;
    rom[78] = 25'b1111111111111111111111111;
    rom[79] = 25'b1111111111111111111111111;
    rom[80] = 25'b1111111111111111111111111;
    rom[81] = 25'b1111111111111111111111111;
    rom[82] = 25'b1111111111111111111111111;
    rom[83] = 25'b1111111111111111111111111;
    rom[84] = 25'b1111111111111111111111111;
    rom[85] = 25'b1111111111111111111111111;
    rom[86] = 25'b1111111111111111111111111;
    rom[87] = 25'b1111111111111111111111111;
    rom[88] = 25'b1111111111111111111111111;
    rom[89] = 25'b1111111111111111111111111;
    rom[90] = 25'b1111111111111111111111111;
    rom[91] = 25'b1111111111111111111111111;
    rom[92] = 25'b1111111111111111111111111;
    rom[93] = 25'b1111111111111111111111111;
    rom[94] = 25'b1111111111111111111111111;
    rom[95] = 25'b1111111111111111111111111;
    rom[96] = 25'b1111111111111111111111111;
    rom[97] = 25'b1111111111111111111111111;
    rom[98] = 25'b1111111111111111111111111;
    rom[99] = 25'b1111111111111111111111111;
    rom[100] = 25'b1111111111111111111111111;
    rom[101] = 25'b1111111111111111111111111;
    rom[102] = 25'b1111111111111111111111111;
    rom[103] = 25'b1111111111111111111111111;
    rom[104] = 25'b1111111111111111111111111;
    rom[105] = 25'b1111111111111111111111111;
    rom[106] = 25'b1111111111111111111111111;
    rom[107] = 25'b1111111111111111111111111;
    rom[108] = 25'b1111111111111111111111111;
    rom[109] = 25'b1111111111111111111111111;
    rom[110] = 25'b1111111111111111111111111;
    rom[111] = 25'b1111111111111111111111111;
    rom[112] = 25'b1111111111111111111111111;
    rom[113] = 25'b1111111111111111111111111;
    rom[114] = 25'b1111111111111111111111111;
    rom[115] = 25'b1111111111111111111111111;
    rom[116] = 25'b1111111111111111111111111;
    rom[117] = 25'b1111111111111111111111111;
    rom[118] = 25'b1111111111111111111111111;
    rom[119] = 25'b1111111111111111111111111;
    rom[120] = 25'b1111111111111111111111111;
    rom[121] = 25'b1111111111111111111111111;
    rom[122] = 25'b1111111111111111111111111;
    rom[123] = 25'b1111111111111111111111111;
    rom[124] = 25'b1111111111111111111111111;
    rom[125] = 25'b1111111111111111111111111;
    rom[126] = 25'b1111111111111111111111111;
    rom[127] = 25'b1111111111111111111111111;
    rom[128] = 25'b1111111111111111111111111;
    rom[129] = 25'b1111111111111111111111111;
    rom[130] = 25'b1111111111111111111111111;
    rom[131] = 25'b1111111111111111111111111;
    rom[132] = 25'b1111111111111111111111111;
    rom[133] = 25'b1111111111111111111111111;
    rom[134] = 25'b1111111111111111111111111;
    rom[135] = 25'b1111111111111111111111111;
    rom[136] = 25'b1111111111111111111111111;
    rom[137] = 25'b1111111111111111111111111;
    rom[138] = 25'b1111111111111111111111111;
    rom[139] = 25'b1111111111111111111111111;
    rom[140] = 25'b1111111111111111111111111;
    rom[141] = 25'b1111111111111111111111111;
    rom[142] = 25'b1111111111111111111111111;
    rom[143] = 25'b1111111111111111111111111;
    rom[144] = 25'b1111111111111111111111111;
    rom[145] = 25'b1111111111111111111111111;
    rom[146] = 25'b1111111111111111111111111;
    rom[147] = 25'b1111111111111111111111111;
    rom[148] = 25'b1111111111111111111111111;
    rom[149] = 25'b1111111111111111111111111;
    rom[150] = 25'b1111111111111111111111111;
    rom[151] = 25'b1111111111111111111111111;
    rom[152] = 25'b1111111111111111111111111;
    rom[153] = 25'b1111111111111111111111111;
    rom[154] = 25'b1111111111111111111111111;
    rom[155] = 25'b1111111111111111111111111;
    rom[156] = 25'b1111111111111111111111111;
    rom[157] = 25'b1111111111111111111111111;
    rom[158] = 25'b1111111111111111111111111;
    rom[159] = 25'b1111111111111111111111111;
    rom[160] = 25'b1111111111111111111111111;
    rom[161] = 25'b1111111111111111111111111;
    rom[162] = 25'b1111111111111111111111111;
    rom[163] = 25'b1111111111111111111111111;
    rom[164] = 25'b1111111111111111111111111;
    rom[165] = 25'b1111111111111111111111111;
    rom[166] = 25'b1111111111111111111111111;
    rom[167] = 25'b1111111111111111111111111;
    rom[168] = 25'b1111111111111111111111111;
    rom[169] = 25'b1111111111111111111111111;
    rom[170] = 25'b1111111111111111111111111;
    rom[171] = 25'b1111111111111111111111111;
    rom[172] = 25'b1111111111111111111111111;
    rom[173] = 25'b1111111111111111111111111;
    rom[174] = 25'b1111111111111111111111111;
    rom[175] = 25'b1111111111111111111111111;
    rom[176] = 25'b1111111111111111111111111;
    rom[177] = 25'b1111111111111111111111111;
    rom[178] = 25'b1111111111111111111111111;
    rom[179] = 25'b1111111111111111111111111;
    rom[180] = 25'b1111111111111111111111111;
    rom[181] = 25'b1111111111111111111111111;
    rom[182] = 25'b1111111111111111111111111;
    rom[183] = 25'b1111111111111111111111111;
    rom[184] = 25'b1111111111111111111111111;
    rom[185] = 25'b1111111111111111111111111;
    rom[186] = 25'b1111111111111111111111111;
    rom[187] = 25'b1111111111111111111111111;
    rom[188] = 25'b1111111111111111111111111;
    rom[189] = 25'b1111111111111111111111111;
    rom[190] = 25'b1111111111111111111111111;
    rom[191] = 25'b1111111111111111111111111;
    rom[192] = 25'b1111111111111111111111111;
    rom[193] = 25'b1111111111111111111111111;
    rom[194] = 25'b1111111111111111111111111;
    rom[195] = 25'b1111111111111111111111111;
    rom[196] = 25'b1111111111111111111111111;
    rom[197] = 25'b1111111111111111111111111;
    rom[198] = 25'b1111111111111111111111111;
    rom[199] = 25'b1111111111111111111111111;
    rom[200] = 25'b1111111111111111111111111;
    rom[201] = 25'b1111111111111111111111111;
    rom[202] = 25'b1111111111111111111111111;
    rom[203] = 25'b1111111111111111111111111;
    rom[204] = 25'b1111111111111111111111111;
    rom[205] = 25'b1111111111111111111111111;
    rom[206] = 25'b1111111111111111111111111;
    rom[207] = 25'b1111111111111111111111111;
    rom[208] = 25'b1111111111111111111111111;
    rom[209] = 25'b1111111111111111111111111;
    rom[210] = 25'b1111111111111111111111111;
    rom[211] = 25'b1111111111111111111111111;
    rom[212] = 25'b1111111111111111111111111;
    rom[213] = 25'b1111111111111111111111111;
    rom[214] = 25'b1111111111111111111111111;
    rom[215] = 25'b1111111111111111111111111;
    rom[216] = 25'b1111111111111111111111111;
    rom[217] = 25'b1111111111111111111111111;
    rom[218] = 25'b1111111111111111111111111;
    rom[219] = 25'b1111111111111111111111111;
    rom[220] = 25'b1111111111111111111111111;
    rom[221] = 25'b1111111111111111111111111;
    rom[222] = 25'b1111111111111111111111111;
    rom[223] = 25'b1111111111111111111111111;
    rom[224] = 25'b1111111111111111111111111;
    rom[225] = 25'b1111111111111111111111111;
    rom[226] = 25'b1111111111111111111111111;
    rom[227] = 25'b1111111111111111111111111;
    rom[228] = 25'b1111111111111111111111111;
    rom[229] = 25'b1111111111111111111111111;
    rom[230] = 25'b1111111111111111111111111;
    rom[231] = 25'b1111111111111111111111111;
    rom[232] = 25'b1111111111111111111111111;
    rom[233] = 25'b1111111111111111111111111;
    rom[234] = 25'b1111111111111111111111111;
    rom[235] = 25'b1111111111111111111111111;
    rom[236] = 25'b1111111111111111111111111;
    rom[237] = 25'b1111111111111111111111111;
    rom[238] = 25'b1111111111111111111111111;
    rom[239] = 25'b1111111111111111111111111;
    rom[240] = 25'b1111111111111111111111111;
    rom[241] = 25'b1111111111111111111111111;
    rom[242] = 25'b1111111111111111111111111;
    rom[243] = 25'b1111111111111111111111111;
    rom[244] = 25'b1111111111111111111111111;
    rom[245] = 25'b1111111111111111111111111;
    rom[246] = 25'b1111111111111111111111111;
    rom[247] = 25'b1111111111111111111111111;
    rom[248] = 25'b1111111111111111111111111;
    rom[249] = 25'b1111111111111111111111111;
    rom[250] = 25'b1111111111111111111111111;
    rom[251] = 25'b1111111111111111111111111;
    rom[252] = 25'b1111111111111111111111111;
    rom[253] = 25'b1111111111111111111111111;
    rom[254] = 25'b1111111111111111111111111;
    rom[255] = 25'b1111111111111111111111111;
    rom[256] = 25'b1111111111111111111111111;
    rom[257] = 25'b1111111111111111111111111;
    rom[258] = 25'b1111111111111111111111111;
    rom[259] = 25'b1111111111111111111111111;
    rom[260] = 25'b1111111111111111111111111;
    rom[261] = 25'b1111111111111111111111111;
    rom[262] = 25'b1111111111111111111111111;
    rom[263] = 25'b1111111111111111111111111;
    rom[264] = 25'b1111111111111111111111111;
    rom[265] = 25'b1111111111111111111111111;
    rom[266] = 25'b1111111111111111111111111;
    rom[267] = 25'b1111111111111111111111111;
    rom[268] = 25'b1111111111111111111111111;
    rom[269] = 25'b1111111111111111111111111;
    rom[270] = 25'b1111111111111111111111111;
    rom[271] = 25'b1111111111111111111111111;
    rom[272] = 25'b1111111111111111111111111;
    rom[273] = 25'b1111111111111111111111111;
    rom[274] = 25'b1111111111111111111111111;
    rom[275] = 25'b1111111111111111111111111;
    rom[276] = 25'b1111111111111111111111111;
    rom[277] = 25'b1111111111111111111111111;
    rom[278] = 25'b1111111111111111111111111;
    rom[279] = 25'b1111111111111111111111111;
    rom[280] = 25'b1111111111111111111111111;
    rom[281] = 25'b1111111111111111111111111;
    rom[282] = 25'b1111111111111111111111111;
    rom[283] = 25'b1111111111111111111111111;
    rom[284] = 25'b1111111111111111111111111;
    rom[285] = 25'b1111111111111111111111111;
    rom[286] = 25'b1111111111111111111111111;
    rom[287] = 25'b1111111111111111111111111;
    rom[288] = 25'b1111111111111111111111111;
    rom[289] = 25'b1111111111111111111111111;
    rom[290] = 25'b0000000000000000000000000;
    rom[291] = 25'b0000000000000000000000000;
    rom[292] = 25'b0000000000000000000000000;
    rom[293] = 25'b0000000000000000000000000;
    rom[294] = 25'b0000000000000000000000000;
    rom[295] = 25'b0000000000000000000000000;
    rom[296] = 25'b0000000000000000000000000;
    rom[297] = 25'b0000000000000000000000000;
    rom[298] = 25'b0000000000000000000000000;
    rom[299] = 25'b0000000000000000000000000;
    rom[300] = 25'b0000000000000000000000000;
    rom[301] = 25'b0000000000000000000000000;
    rom[302] = 25'b0000000000000000000000000;
    rom[303] = 25'b0000000000000000000000000;
    rom[304] = 25'b0000000000000000000000000;
    rom[305] = 25'b0000000000000000000000000;
    rom[306] = 25'b0000000000000000000000000;
    rom[307] = 25'b0000000000000000000000000;
    rom[308] = 25'b0000000000000000000000000;
    rom[309] = 25'b0000000000000000000000000;
    rom[310] = 25'b0000000000000000000000000;
    rom[311] = 25'b0000000000000000000000000;
    rom[312] = 25'b0000000000000000000000000;
    rom[313] = 25'b0000000000000000000000000;
    rom[314] = 25'b0000000000000000000000000;
    rom[315] = 25'b0000000000000000000000000;
    rom[316] = 25'b0000000000000000000000000;
    rom[317] = 25'b0000000000000000000000000;
    rom[318] = 25'b0000000000000000000000000;
    rom[319] = 25'b0000000000000000000000000;
    rom[320] = 25'b0000000000000000000000000;
    rom[321] = 25'b0000000000000000000000000;
    rom[322] = 25'b0000000000000000000000000;
    rom[323] = 25'b0000000000000000000000000;
    rom[324] = 25'b0000000000000000000000000;
    rom[325] = 25'b0000000000000000000000000;
    rom[326] = 25'b0000000000000000000000000;
    rom[327] = 25'b0000000000000000000000000;
    rom[328] = 25'b0000000000000000000000000;
    rom[329] = 25'b0000000000000000000000000;
    rom[330] = 25'b0000000000000000000000000;
    rom[331] = 25'b0000000000000000000000000;
    rom[332] = 25'b0000000000000000000000000;
    rom[333] = 25'b0000000000000000000000000;
    rom[334] = 25'b0000000000000000000000000;
    rom[335] = 25'b0000000000000000000000000;
    rom[336] = 25'b0000000000000000000000000;
    rom[337] = 25'b0000000000000000000000000;
    rom[338] = 25'b0000000000000000000000000;
    rom[339] = 25'b0000000000000000000000000;
    rom[340] = 25'b0000000000000000000000000;
    rom[341] = 25'b0000000000000000000000000;
    rom[342] = 25'b0000000000000000000000000;
    rom[343] = 25'b0000000000000000000000000;
    rom[344] = 25'b0000000000000000000000000;
    rom[345] = 25'b0000000000000000000000000;
    rom[346] = 25'b0000000000000000000000000;
    rom[347] = 25'b0000000000000000000000000;
    rom[348] = 25'b0000000000000000000000000;
    rom[349] = 25'b0000000000000000000000000;
    rom[350] = 25'b0000000000000000000000000;
    rom[351] = 25'b0000000000000000000000000;
    rom[352] = 25'b0000000000000000000000000;
    rom[353] = 25'b0000000000000000000000000;
    rom[354] = 25'b0000000000000000000000000;
    rom[355] = 25'b0000000000000000000000000;
    rom[356] = 25'b0000000000000000000000000;
    rom[357] = 25'b0000000000000000000000000;
    rom[358] = 25'b0000000000000000000000000;
    rom[359] = 25'b0000000000000000000000000;
    rom[360] = 25'b0000000000000000000000000;
    rom[361] = 25'b0000000000000000000000000;
    rom[362] = 25'b0000000000000000000000000;
    rom[363] = 25'b0000000000000000000000000;
    rom[364] = 25'b0000000000000000000000000;
    rom[365] = 25'b0000000000000000000000000;
    rom[366] = 25'b0000000000000000000000000;
    rom[367] = 25'b0000000000000000000000000;
    rom[368] = 25'b0000000000000000000000000;
    rom[369] = 25'b0000000000000000000000000;
    rom[370] = 25'b0000000000000000000000000;
    rom[371] = 25'b0000000000000000000000000;
    rom[372] = 25'b0000000000000000000000000;
    rom[373] = 25'b0000000000000000000000000;
    rom[374] = 25'b0000000000000000000000000;
    rom[375] = 25'b0000000000000000000000000;
    rom[376] = 25'b0000000000000000000000000;
    rom[377] = 25'b0000000000000000000000000;
    rom[378] = 25'b0000000000000000000000000;
    rom[379] = 25'b0000000000000000000000000;
    rom[380] = 25'b0000000000000000000000000;
    rom[381] = 25'b0000000000000000000000000;
    rom[382] = 25'b0000000000000000000000000;
    rom[383] = 25'b0000000000000000000000000;
    rom[384] = 25'b0000000000000000000000000;
    rom[385] = 25'b0000000000000000000000000;
    rom[386] = 25'b0000000000000000000000000;
    rom[387] = 25'b0000000000000000000000000;
    rom[388] = 25'b0000000000000000000000000;
    rom[389] = 25'b0000000000000000000000000;
    rom[390] = 25'b0000000000000000000000000;
    rom[391] = 25'b0000000000000000000000000;
    rom[392] = 25'b0000000000000000000000000;
    rom[393] = 25'b0000000000000000000000000;
    rom[394] = 25'b0000000000000000000000000;
    rom[395] = 25'b0000000000000000000000000;
    rom[396] = 25'b0000000000000000000000000;
    rom[397] = 25'b0000000000000000000000000;
    rom[398] = 25'b0000000000000000000000000;
    rom[399] = 25'b0000000000000000000000000;
    rom[400] = 25'b0000000000000000000000000;
    rom[401] = 25'b0000000000000000000000000;
    rom[402] = 25'b0000000000000000000000000;
    rom[403] = 25'b0000000000000000000000000;
    rom[404] = 25'b0000000000000000000000000;
    rom[405] = 25'b0000000000000000000000000;
    rom[406] = 25'b0000000000000000000000000;
    rom[407] = 25'b0000000000000000000000000;
    rom[408] = 25'b0000000000000000000000000;
    rom[409] = 25'b0000000000000000000000000;
    rom[410] = 25'b0000000000000000000000000;
    rom[411] = 25'b0000000000000000000000000;
    rom[412] = 25'b0000000000000000000000000;
    rom[413] = 25'b0000000000000000000000000;
    rom[414] = 25'b0000000000000000000000000;
    rom[415] = 25'b0000000000000000000000000;
    rom[416] = 25'b0000000000000000000000000;
    rom[417] = 25'b0000000000000000000000000;
    rom[418] = 25'b0000000000000000000000000;
    rom[419] = 25'b0000000000000000000000000;
    rom[420] = 25'b0000000000000000000000000;
    rom[421] = 25'b0000000000000000000000000;
    rom[422] = 25'b0000000000000000000000000;
    rom[423] = 25'b0000000000000000000000000;
    rom[424] = 25'b0000000000000000000000000;
    rom[425] = 25'b0000000000000000000000000;
    rom[426] = 25'b0000000000000000000000000;
    rom[427] = 25'b0000000000000000000000000;
    rom[428] = 25'b0000000000000000000000000;
    rom[429] = 25'b0000000000000000000000000;
    rom[430] = 25'b0000000000000000000000000;
    rom[431] = 25'b0000000000000000000000000;
    rom[432] = 25'b0000000000000000000000000;
    rom[433] = 25'b0000000000000000000000000;
    rom[434] = 25'b0000000000000000000000000;
    rom[435] = 25'b0000000000000000000000000;
    rom[436] = 25'b0000000000000000000000000;
    rom[437] = 25'b0000000000000000000000000;
    rom[438] = 25'b0000000000000000000000000;
    rom[439] = 25'b0000000000000000000000000;
    rom[440] = 25'b0000000000000000000000000;
    rom[441] = 25'b0000000000000000000000000;
    rom[442] = 25'b0000000000000000000000000;
    rom[443] = 25'b0000000000000000000000000;
    rom[444] = 25'b0000000000000000000000000;
    rom[445] = 25'b0000000000000000000000000;
    rom[446] = 25'b0000000000000000000000000;
    rom[447] = 25'b0000000000000000000000000;
    rom[448] = 25'b0000000000000000000000000;
    rom[449] = 25'b0000000000000000000000000;
    rom[450] = 25'b0000000000000000000000000;
    rom[451] = 25'b0000000000000000000000001;
    rom[452] = 25'b0000000000000000000000001;
    rom[453] = 25'b0000000000000000000000001;
    rom[454] = 25'b0000000000000000000000001;
    rom[455] = 25'b0000000000000000000000001;
    rom[456] = 25'b0000000000000000000000001;
    rom[457] = 25'b0000000000000000000000001;
    rom[458] = 25'b0000000000000000000000001;
    rom[459] = 25'b0000000000000000000000001;
    rom[460] = 25'b0000000000000000000000001;
    rom[461] = 25'b0000000000000000000000001;
    rom[462] = 25'b0000000000000000000000001;
    rom[463] = 25'b0000000000000000000000001;
    rom[464] = 25'b0000000000000000000000001;
    rom[465] = 25'b0000000000000000000000001;
    rom[466] = 25'b0000000000000000000000001;
    rom[467] = 25'b0000000000000000000000001;
    rom[468] = 25'b0000000000000000000000001;
    rom[469] = 25'b0000000000000000000000001;
    rom[470] = 25'b0000000000000000000000001;
    rom[471] = 25'b0000000000000000000000001;
    rom[472] = 25'b0000000000000000000000001;
    rom[473] = 25'b0000000000000000000000001;
    rom[474] = 25'b0000000000000000000000001;
    rom[475] = 25'b0000000000000000000000001;
    rom[476] = 25'b0000000000000000000000001;
    rom[477] = 25'b0000000000000000000000001;
    rom[478] = 25'b0000000000000000000000001;
    rom[479] = 25'b0000000000000000000000001;
    rom[480] = 25'b0000000000000000000000001;
    rom[481] = 25'b0000000000000000000000001;
    rom[482] = 25'b0000000000000000000000001;
    rom[483] = 25'b0000000000000000000000001;
    rom[484] = 25'b0000000000000000000000001;
    rom[485] = 25'b0000000000000000000000010;
    rom[486] = 25'b0000000000000000000000010;
    rom[487] = 25'b0000000000000000000000010;
    rom[488] = 25'b0000000000000000000000010;
    rom[489] = 25'b0000000000000000000000010;
    rom[490] = 25'b0000000000000000000000010;
    rom[491] = 25'b0000000000000000000000010;
    rom[492] = 25'b0000000000000000000000010;
    rom[493] = 25'b0000000000000000000000010;
    rom[494] = 25'b0000000000000000000000010;
    rom[495] = 25'b0000000000000000000000010;
    rom[496] = 25'b0000000000000000000000010;
    rom[497] = 25'b0000000000000000000000010;
    rom[498] = 25'b0000000000000000000000010;
    rom[499] = 25'b0000000000000000000000010;
    rom[500] = 25'b0000000000000000000000010;
    rom[501] = 25'b0000000000000000000000010;
    rom[502] = 25'b0000000000000000000000010;
    rom[503] = 25'b0000000000000000000000010;
    rom[504] = 25'b0000000000000000000000010;
    rom[505] = 25'b0000000000000000000000010;
    rom[506] = 25'b0000000000000000000000010;
    rom[507] = 25'b0000000000000000000000010;
    rom[508] = 25'b0000000000000000000000010;
    rom[509] = 25'b0000000000000000000000010;
    rom[510] = 25'b0000000000000000000000010;
    rom[511] = 25'b0000000000000000000000010;
    rom[512] = 25'b0000000000000000000000010;
    rom[513] = 25'b0000000000000000000000010;
    rom[514] = 25'b0000000000000000000000010;
    rom[515] = 25'b0000000000000000000000010;
    rom[516] = 25'b0000000000000000000000010;
    rom[517] = 25'b0000000000000000000000011;
    rom[518] = 25'b0000000000000000000000011;
    rom[519] = 25'b0000000000000000000000011;
    rom[520] = 25'b0000000000000000000000011;
    rom[521] = 25'b0000000000000000000000011;
    rom[522] = 25'b0000000000000000000000011;
    rom[523] = 25'b0000000000000000000000011;
    rom[524] = 25'b0000000000000000000000011;
    rom[525] = 25'b0000000000000000000000011;
    rom[526] = 25'b0000000000000000000000011;
    rom[527] = 25'b0000000000000000000000011;
    rom[528] = 25'b0000000000000000000000011;
    rom[529] = 25'b0000000000000000000000011;
    rom[530] = 25'b0000000000000000000000011;
    rom[531] = 25'b0000000000000000000000011;
    rom[532] = 25'b0000000000000000000000011;
    rom[533] = 25'b0000000000000000000000011;
    rom[534] = 25'b0000000000000000000000011;
    rom[535] = 25'b0000000000000000000000011;
    rom[536] = 25'b0000000000000000000000011;
    rom[537] = 25'b0000000000000000000000011;
    rom[538] = 25'b0000000000000000000000011;
    rom[539] = 25'b0000000000000000000000011;
    rom[540] = 25'b0000000000000000000000011;
    rom[541] = 25'b0000000000000000000000011;
    rom[542] = 25'b0000000000000000000000011;
    rom[543] = 25'b0000000000000000000000011;
    rom[544] = 25'b0000000000000000000000011;
    rom[545] = 25'b0000000000000000000000011;
    rom[546] = 25'b0000000000000000000000100;
    rom[547] = 25'b0000000000000000000000100;
    rom[548] = 25'b0000000000000000000000100;
    rom[549] = 25'b0000000000000000000000100;
    rom[550] = 25'b0000000000000000000000100;
    rom[551] = 25'b0000000000000000000000100;
    rom[552] = 25'b0000000000000000000000100;
    rom[553] = 25'b0000000000000000000000100;
    rom[554] = 25'b0000000000000000000000100;
    rom[555] = 25'b0000000000000000000000100;
    rom[556] = 25'b0000000000000000000000100;
    rom[557] = 25'b0000000000000000000000100;
    rom[558] = 25'b0000000000000000000000100;
    rom[559] = 25'b0000000000000000000000100;
    rom[560] = 25'b0000000000000000000000100;
    rom[561] = 25'b0000000000000000000000100;
    rom[562] = 25'b0000000000000000000000100;
    rom[563] = 25'b0000000000000000000000100;
    rom[564] = 25'b0000000000000000000000100;
    rom[565] = 25'b0000000000000000000000100;
    rom[566] = 25'b0000000000000000000000100;
    rom[567] = 25'b0000000000000000000000100;
    rom[568] = 25'b0000000000000000000000100;
    rom[569] = 25'b0000000000000000000000100;
    rom[570] = 25'b0000000000000000000000100;
    rom[571] = 25'b0000000000000000000000100;
    rom[572] = 25'b0000000000000000000000100;
    rom[573] = 25'b0000000000000000000000100;
    rom[574] = 25'b0000000000000000000000100;
    rom[575] = 25'b0000000000000000000000101;
    rom[576] = 25'b0000000000000000000000101;
    rom[577] = 25'b0000000000000000000000101;
    rom[578] = 25'b0000000000000000000000101;
    rom[579] = 25'b0000000000000000000000101;
    rom[580] = 25'b0000000000000000000000101;
    rom[581] = 25'b0000000000000000000000101;
    rom[582] = 25'b0000000000000000000000101;
    rom[583] = 25'b0000000000000000000000101;
    rom[584] = 25'b0000000000000000000000101;
    rom[585] = 25'b0000000000000000000000101;
    rom[586] = 25'b0000000000000000000000101;
    rom[587] = 25'b0000000000000000000000101;
    rom[588] = 25'b0000000000000000000000101;
    rom[589] = 25'b0000000000000000000000101;
    rom[590] = 25'b0000000000000000000000101;
    rom[591] = 25'b0000000000000000000000101;
    rom[592] = 25'b0000000000000000000000101;
    rom[593] = 25'b0000000000000000000000101;
    rom[594] = 25'b0000000000000000000000101;
    rom[595] = 25'b0000000000000000000000101;
    rom[596] = 25'b0000000000000000000000101;
    rom[597] = 25'b0000000000000000000000101;
    rom[598] = 25'b0000000000000000000000101;
    rom[599] = 25'b0000000000000000000000101;
    rom[600] = 25'b0000000000000000000000101;
    rom[601] = 25'b0000000000000000000000101;
    rom[602] = 25'b0000000000000000000000101;
    rom[603] = 25'b0000000000000000000000101;
    rom[604] = 25'b0000000000000000000000101;
    rom[605] = 25'b0000000000000000000000101;
    rom[606] = 25'b0000000000000000000000101;
    rom[607] = 25'b0000000000000000000000101;
    rom[608] = 25'b0000000000000000000000101;
    rom[609] = 25'b0000000000000000000000101;
    rom[610] = 25'b0000000000000000000000101;
    rom[611] = 25'b0000000000000000000000101;
    rom[612] = 25'b0000000000000000000000101;
    rom[613] = 25'b0000000000000000000000101;
    rom[614] = 25'b0000000000000000000000101;
    rom[615] = 25'b0000000000000000000000101;
    rom[616] = 25'b0000000000000000000000101;
    rom[617] = 25'b0000000000000000000000101;
    rom[618] = 25'b0000000000000000000000101;
    rom[619] = 25'b0000000000000000000000101;
    rom[620] = 25'b0000000000000000000000101;
    rom[621] = 25'b0000000000000000000000101;
    rom[622] = 25'b0000000000000000000000101;
    rom[623] = 25'b0000000000000000000000101;
    rom[624] = 25'b0000000000000000000000101;
    rom[625] = 25'b0000000000000000000000101;
    rom[626] = 25'b0000000000000000000000101;
    rom[627] = 25'b0000000000000000000000101;
    rom[628] = 25'b0000000000000000000000101;
    rom[629] = 25'b0000000000000000000000101;
    rom[630] = 25'b0000000000000000000000101;
    rom[631] = 25'b0000000000000000000000101;
    rom[632] = 25'b0000000000000000000000101;
    rom[633] = 25'b0000000000000000000000101;
    rom[634] = 25'b0000000000000000000000110;
    rom[635] = 25'b0000000000000000000000110;
    rom[636] = 25'b0000000000000000000000110;
    rom[637] = 25'b0000000000000000000000110;
    rom[638] = 25'b0000000000000000000000110;
    rom[639] = 25'b0000000000000000000000110;
    rom[640] = 25'b0000000000000000000000110;
    rom[641] = 25'b0000000000000000000000110;
    rom[642] = 25'b0000000000000000000000110;
    rom[643] = 25'b0000000000000000000000110;
    rom[644] = 25'b0000000000000000000000110;
    rom[645] = 25'b0000000000000000000000110;
    rom[646] = 25'b0000000000000000000000110;
    rom[647] = 25'b0000000000000000000000110;
    rom[648] = 25'b0000000000000000000000110;
    rom[649] = 25'b0000000000000000000000110;
    rom[650] = 25'b0000000000000000000000110;
    rom[651] = 25'b0000000000000000000000110;
    rom[652] = 25'b0000000000000000000000110;
    rom[653] = 25'b0000000000000000000000110;
    rom[654] = 25'b0000000000000000000000110;
    rom[655] = 25'b0000000000000000000000110;
    rom[656] = 25'b0000000000000000000000110;
    rom[657] = 25'b0000000000000000000000110;
    rom[658] = 25'b0000000000000000000000110;
    rom[659] = 25'b0000000000000000000000110;
    rom[660] = 25'b0000000000000000000000110;
    rom[661] = 25'b0000000000000000000000110;
    rom[662] = 25'b0000000000000000000000110;
    rom[663] = 25'b0000000000000000000000110;
    rom[664] = 25'b0000000000000000000000110;
    rom[665] = 25'b0000000000000000000000110;
    rom[666] = 25'b0000000000000000000000110;
    rom[667] = 25'b0000000000000000000000110;
    rom[668] = 25'b0000000000000000000000111;
    rom[669] = 25'b0000000000000000000000111;
    rom[670] = 25'b0000000000000000000000111;
    rom[671] = 25'b0000000000000000000000111;
    rom[672] = 25'b0000000000000000000000111;
    rom[673] = 25'b0000000000000000000000111;
    rom[674] = 25'b0000000000000000000000111;
    rom[675] = 25'b0000000000000000000000111;
    rom[676] = 25'b0000000000000000000000111;
    rom[677] = 25'b0000000000000000000000111;
    rom[678] = 25'b0000000000000000000000111;
    rom[679] = 25'b0000000000000000000000111;
    rom[680] = 25'b0000000000000000000000111;
    rom[681] = 25'b0000000000000000000000111;
    rom[682] = 25'b0000000000000000000000111;
    rom[683] = 25'b0000000000000000000000111;
    rom[684] = 25'b0000000000000000000000111;
    rom[685] = 25'b0000000000000000000000111;
    rom[686] = 25'b0000000000000000000000111;
    rom[687] = 25'b0000000000000000000000111;
    rom[688] = 25'b0000000000000000000000111;
    rom[689] = 25'b0000000000000000000000111;
    rom[690] = 25'b0000000000000000000000111;
    rom[691] = 25'b0000000000000000000000111;
    rom[692] = 25'b0000000000000000000000111;
    rom[693] = 25'b0000000000000000000000111;
    rom[694] = 25'b0000000000000000000000111;
    rom[695] = 25'b0000000000000000000000111;
    rom[696] = 25'b0000000000000000000000111;
    rom[697] = 25'b0000000000000000000000111;
    rom[698] = 25'b0000000000000000000000111;
    rom[699] = 25'b0000000000000000000000111;
    rom[700] = 25'b0000000000000000000000111;
    rom[701] = 25'b0000000000000000000000111;
    rom[702] = 25'b0000000000000000000000111;
    rom[703] = 25'b0000000000000000000000111;
    rom[704] = 25'b0000000000000000000000111;
    rom[705] = 25'b0000000000000000000000111;
    rom[706] = 25'b0000000000000000000000111;
    rom[707] = 25'b0000000000000000000000111;
    rom[708] = 25'b0000000000000000000000111;
    rom[709] = 25'b0000000000000000000000111;
    rom[710] = 25'b0000000000000000000001000;
    rom[711] = 25'b0000000000000000000001000;
    rom[712] = 25'b0000000000000000000001000;
    rom[713] = 25'b0000000000000000000001000;
    rom[714] = 25'b0000000000000000000001000;
    rom[715] = 25'b0000000000000000000001000;
    rom[716] = 25'b0000000000000000000001000;
    rom[717] = 25'b0000000000000000000001000;
    rom[718] = 25'b0000000000000000000001000;
    rom[719] = 25'b0000000000000000000001000;
    rom[720] = 25'b0000000000000000000001000;
    rom[721] = 25'b0000000000000000000001000;
    rom[722] = 25'b0000000000000000000001000;
    rom[723] = 25'b0000000000000000000001000;
    rom[724] = 25'b0000000000000000000001000;
    rom[725] = 25'b0000000000000000000001000;
    rom[726] = 25'b0000000000000000000001000;
    rom[727] = 25'b0000000000000000000001000;
    rom[728] = 25'b0000000000000000000001000;
    rom[729] = 25'b0000000000000000000001000;
    rom[730] = 25'b0000000000000000000001000;
    rom[731] = 25'b0000000000000000000001000;
    rom[732] = 25'b0000000000000000000001000;
    rom[733] = 25'b0000000000000000000001000;
    rom[734] = 25'b0000000000000000000001000;
    rom[735] = 25'b0000000000000000000001000;
    rom[736] = 25'b0000000000000000000001000;
    rom[737] = 25'b0000000000000000000001000;
    rom[738] = 25'b0000000000000000000001000;
    rom[739] = 25'b0000000000000000000001000;
    rom[740] = 25'b0000000000000000000001000;
    rom[741] = 25'b0000000000000000000001000;
    rom[742] = 25'b0000000000000000000001000;
    rom[743] = 25'b0000000000000000000001000;
    rom[744] = 25'b0000000000000000000001000;
    rom[745] = 25'b0000000000000000000001000;
    rom[746] = 25'b0000000000000000000001000;
    rom[747] = 25'b0000000000000000000001000;
    rom[748] = 25'b0000000000000000000001000;
    rom[749] = 25'b0000000000000000000001000;
    rom[750] = 25'b0000000000000000000001000;
    rom[751] = 25'b0000000000000000000001000;
    rom[752] = 25'b0000000000000000000001000;
    rom[753] = 25'b0000000000000000000001000;
    rom[754] = 25'b0000000000000000000001000;
    rom[755] = 25'b0000000000000000000001000;
    rom[756] = 25'b0000000000000000000001000;
    rom[757] = 25'b0000000000000000000001000;
    rom[758] = 25'b0000000000000000000001000;
    rom[759] = 25'b0000000000000000000001000;
    rom[760] = 25'b0000000000000000000001000;
    rom[761] = 25'b0000000000000000000001000;
    rom[762] = 25'b0000000000000000000001000;
    rom[763] = 25'b0000000000000000000001000;
    rom[764] = 25'b0000000000000000000001000;
    rom[765] = 25'b0000000000000000000001000;
    rom[766] = 25'b0000000000000000000001000;
    rom[767] = 25'b0000000000000000000001000;
    rom[768] = 25'b0000000000000000000001000;
    rom[769] = 25'b0000000000000000000001000;
    rom[770] = 25'b0000000000000000000001000;
    rom[771] = 25'b0000000000000000000001000;
    rom[772] = 25'b0000000000000000000001000;
    rom[773] = 25'b0000000000000000000001000;
    rom[774] = 25'b0000000000000000000001000;
    rom[775] = 25'b0000000000000000000001000;
    rom[776] = 25'b0000000000000000000001000;
    rom[777] = 25'b0000000000000000000001000;
    rom[778] = 25'b0000000000000000000001000;
    rom[779] = 25'b0000000000000000000001000;
    rom[780] = 25'b0000000000000000000001000;
    rom[781] = 25'b0000000000000000000001000;
    rom[782] = 25'b0000000000000000000001000;
    rom[783] = 25'b0000000000000000000001000;
    rom[784] = 25'b0000000000000000000001000;
    rom[785] = 25'b0000000000000000000001000;
    rom[786] = 25'b0000000000000000000001000;
    rom[787] = 25'b0000000000000000000001000;
    rom[788] = 25'b0000000000000000000001000;
    rom[789] = 25'b0000000000000000000001000;
    rom[790] = 25'b0000000000000000000001000;
    rom[791] = 25'b0000000000000000000001000;
    rom[792] = 25'b0000000000000000000001000;
    rom[793] = 25'b0000000000000000000001000;
    rom[794] = 25'b0000000000000000000001000;
    rom[795] = 25'b0000000000000000000001000;
    rom[796] = 25'b0000000000000000000001000;
    rom[797] = 25'b0000000000000000000001000;
    rom[798] = 25'b0000000000000000000001000;
    rom[799] = 25'b0000000000000000000001000;
    rom[800] = 25'b0000000000000000000001000;
    rom[801] = 25'b0000000000000000000001000;
    rom[802] = 25'b0000000000000000000001000;
    rom[803] = 25'b0000000000000000000001000;
    rom[804] = 25'b0000000000000000000001000;
    rom[805] = 25'b0000000000000000000001000;
    rom[806] = 25'b0000000000000000000001000;
    rom[807] = 25'b0000000000000000000001000;
    rom[808] = 25'b0000000000000000000001000;
    rom[809] = 25'b0000000000000000000001000;
    rom[810] = 25'b0000000000000000000001000;
    rom[811] = 25'b0000000000000000000001000;
    rom[812] = 25'b0000000000000000000001000;
    rom[813] = 25'b0000000000000000000001000;
    rom[814] = 25'b0000000000000000000001000;
    rom[815] = 25'b0000000000000000000001000;
    rom[816] = 25'b0000000000000000000001000;
    rom[817] = 25'b0000000000000000000001000;
    rom[818] = 25'b0000000000000000000001000;
    rom[819] = 25'b0000000000000000000001000;
    rom[820] = 25'b0000000000000000000001000;
    rom[821] = 25'b0000000000000000000000111;
    rom[822] = 25'b0000000000000000000000111;
    rom[823] = 25'b0000000000000000000000111;
    rom[824] = 25'b0000000000000000000000111;
    rom[825] = 25'b0000000000000000000000111;
    rom[826] = 25'b0000000000000000000000111;
    rom[827] = 25'b0000000000000000000000111;
    rom[828] = 25'b0000000000000000000000111;
    rom[829] = 25'b0000000000000000000000111;
    rom[830] = 25'b0000000000000000000000111;
    rom[831] = 25'b0000000000000000000000111;
    rom[832] = 25'b0000000000000000000000111;
    rom[833] = 25'b0000000000000000000000111;
    rom[834] = 25'b0000000000000000000000111;
    rom[835] = 25'b0000000000000000000000111;
    rom[836] = 25'b0000000000000000000000111;
    rom[837] = 25'b0000000000000000000000111;
    rom[838] = 25'b0000000000000000000000111;
    rom[839] = 25'b0000000000000000000000111;
    rom[840] = 25'b0000000000000000000000111;
    rom[841] = 25'b0000000000000000000000111;
    rom[842] = 25'b0000000000000000000000111;
    rom[843] = 25'b0000000000000000000000111;
    rom[844] = 25'b0000000000000000000000111;
    rom[845] = 25'b0000000000000000000000111;
    rom[846] = 25'b0000000000000000000000111;
    rom[847] = 25'b0000000000000000000000111;
    rom[848] = 25'b0000000000000000000000111;
    rom[849] = 25'b0000000000000000000000111;
    rom[850] = 25'b0000000000000000000000111;
    rom[851] = 25'b0000000000000000000000111;
    rom[852] = 25'b0000000000000000000000111;
    rom[853] = 25'b0000000000000000000000110;
    rom[854] = 25'b0000000000000000000000110;
    rom[855] = 25'b0000000000000000000000110;
    rom[856] = 25'b0000000000000000000000110;
    rom[857] = 25'b0000000000000000000000110;
    rom[858] = 25'b0000000000000000000000110;
    rom[859] = 25'b0000000000000000000000110;
    rom[860] = 25'b0000000000000000000000110;
    rom[861] = 25'b0000000000000000000000110;
    rom[862] = 25'b0000000000000000000000110;
    rom[863] = 25'b0000000000000000000000110;
    rom[864] = 25'b0000000000000000000000110;
    rom[865] = 25'b0000000000000000000000110;
    rom[866] = 25'b0000000000000000000000110;
    rom[867] = 25'b0000000000000000000000110;
    rom[868] = 25'b0000000000000000000000110;
    rom[869] = 25'b0000000000000000000000110;
    rom[870] = 25'b0000000000000000000000110;
    rom[871] = 25'b0000000000000000000000110;
    rom[872] = 25'b0000000000000000000000110;
    rom[873] = 25'b0000000000000000000000110;
    rom[874] = 25'b0000000000000000000000101;
    rom[875] = 25'b0000000000000000000000101;
    rom[876] = 25'b0000000000000000000000101;
    rom[877] = 25'b0000000000000000000000101;
    rom[878] = 25'b0000000000000000000000101;
    rom[879] = 25'b0000000000000000000000101;
    rom[880] = 25'b0000000000000000000000101;
    rom[881] = 25'b0000000000000000000000101;
    rom[882] = 25'b0000000000000000000000101;
    rom[883] = 25'b0000000000000000000000101;
    rom[884] = 25'b0000000000000000000000101;
    rom[885] = 25'b0000000000000000000000101;
    rom[886] = 25'b0000000000000000000000101;
    rom[887] = 25'b0000000000000000000000101;
    rom[888] = 25'b0000000000000000000000101;
    rom[889] = 25'b0000000000000000000000101;
    rom[890] = 25'b0000000000000000000000101;
    rom[891] = 25'b0000000000000000000000101;
    rom[892] = 25'b0000000000000000000000101;
    rom[893] = 25'b0000000000000000000000101;
    rom[894] = 25'b0000000000000000000000101;
    rom[895] = 25'b0000000000000000000000101;
    rom[896] = 25'b0000000000000000000000101;
    rom[897] = 25'b0000000000000000000000101;
    rom[898] = 25'b0000000000000000000000101;
    rom[899] = 25'b0000000000000000000000101;
    rom[900] = 25'b0000000000000000000000101;
    rom[901] = 25'b0000000000000000000000101;
    rom[902] = 25'b0000000000000000000000101;
    rom[903] = 25'b0000000000000000000000101;
    rom[904] = 25'b0000000000000000000000101;
    rom[905] = 25'b0000000000000000000000101;
    rom[906] = 25'b0000000000000000000000100;
    rom[907] = 25'b0000000000000000000000100;
    rom[908] = 25'b0000000000000000000000100;
    rom[909] = 25'b0000000000000000000000100;
    rom[910] = 25'b0000000000000000000000100;
    rom[911] = 25'b0000000000000000000000100;
    rom[912] = 25'b0000000000000000000000100;
    rom[913] = 25'b0000000000000000000000100;
    rom[914] = 25'b0000000000000000000000100;
    rom[915] = 25'b0000000000000000000000100;
    rom[916] = 25'b0000000000000000000000100;
    rom[917] = 25'b0000000000000000000000100;
    rom[918] = 25'b0000000000000000000000100;
    rom[919] = 25'b0000000000000000000000011;
    rom[920] = 25'b0000000000000000000000011;
    rom[921] = 25'b0000000000000000000000011;
    rom[922] = 25'b0000000000000000000000011;
    rom[923] = 25'b0000000000000000000000011;
    rom[924] = 25'b0000000000000000000000011;
    rom[925] = 25'b0000000000000000000000011;
    rom[926] = 25'b0000000000000000000000011;
    rom[927] = 25'b0000000000000000000000011;
    rom[928] = 25'b0000000000000000000000011;
    rom[929] = 25'b0000000000000000000000011;
    rom[930] = 25'b0000000000000000000000010;
    rom[931] = 25'b0000000000000000000000010;
    rom[932] = 25'b0000000000000000000000010;
    rom[933] = 25'b0000000000000000000000010;
    rom[934] = 25'b0000000000000000000000010;
    rom[935] = 25'b0000000000000000000000010;
    rom[936] = 25'b0000000000000000000000010;
    rom[937] = 25'b0000000000000000000000010;
    rom[938] = 25'b0000000000000000000000010;
    rom[939] = 25'b0000000000000000000000010;
    rom[940] = 25'b0000000000000000000000010;
    rom[941] = 25'b0000000000000000000000001;
    rom[942] = 25'b0000000000000000000000001;
    rom[943] = 25'b0000000000000000000000001;
    rom[944] = 25'b0000000000000000000000001;
    rom[945] = 25'b0000000000000000000000001;
    rom[946] = 25'b0000000000000000000000001;
    rom[947] = 25'b0000000000000000000000001;
    rom[948] = 25'b0000000000000000000000001;
    rom[949] = 25'b0000000000000000000000001;
    rom[950] = 25'b0000000000000000000000001;
    rom[951] = 25'b0000000000000000000000000;
    rom[952] = 25'b0000000000000000000000000;
    rom[953] = 25'b0000000000000000000000000;
    rom[954] = 25'b0000000000000000000000000;
    rom[955] = 25'b0000000000000000000000000;
    rom[956] = 25'b0000000000000000000000000;
    rom[957] = 25'b0000000000000000000000000;
    rom[958] = 25'b0000000000000000000000000;
    rom[959] = 25'b0000000000000000000000000;
    rom[960] = 25'b0000000000000000000000000;
    rom[961] = 25'b0000000000000000000000000;
    rom[962] = 25'b0000000000000000000000000;
    rom[963] = 25'b0000000000000000000000000;
    rom[964] = 25'b0000000000000000000000000;
    rom[965] = 25'b0000000000000000000000000;
    rom[966] = 25'b0000000000000000000000000;
    rom[967] = 25'b0000000000000000000000000;
    rom[968] = 25'b0000000000000000000000000;
    rom[969] = 25'b0000000000000000000000000;
    rom[970] = 25'b0000000000000000000000000;
    rom[971] = 25'b0000000000000000000000000;
    rom[972] = 25'b0000000000000000000000000;
    rom[973] = 25'b0000000000000000000000000;
    rom[974] = 25'b0000000000000000000000000;
    rom[975] = 25'b0000000000000000000000000;
    rom[976] = 25'b0000000000000000000000000;
    rom[977] = 25'b0000000000000000000000000;
    rom[978] = 25'b1111111111111111111111111;
    rom[979] = 25'b1111111111111111111111111;
    rom[980] = 25'b1111111111111111111111111;
    rom[981] = 25'b1111111111111111111111111;
    rom[982] = 25'b1111111111111111111111111;
    rom[983] = 25'b1111111111111111111111111;
    rom[984] = 25'b1111111111111111111111111;
    rom[985] = 25'b1111111111111111111111111;
    rom[986] = 25'b1111111111111111111111110;
    rom[987] = 25'b1111111111111111111111110;
    rom[988] = 25'b1111111111111111111111110;
    rom[989] = 25'b1111111111111111111111110;
    rom[990] = 25'b1111111111111111111111110;
    rom[991] = 25'b1111111111111111111111110;
    rom[992] = 25'b1111111111111111111111110;
    rom[993] = 25'b1111111111111111111111110;
    rom[994] = 25'b1111111111111111111111101;
    rom[995] = 25'b1111111111111111111111101;
    rom[996] = 25'b1111111111111111111111101;
    rom[997] = 25'b1111111111111111111111101;
    rom[998] = 25'b1111111111111111111111101;
    rom[999] = 25'b1111111111111111111111101;
    rom[1000] = 25'b1111111111111111111111101;
    rom[1001] = 25'b1111111111111111111111100;
    rom[1002] = 25'b1111111111111111111111100;
    rom[1003] = 25'b1111111111111111111111100;
    rom[1004] = 25'b1111111111111111111111100;
    rom[1005] = 25'b1111111111111111111111100;
    rom[1006] = 25'b1111111111111111111111100;
    rom[1007] = 25'b1111111111111111111111100;
    rom[1008] = 25'b1111111111111111111111011;
    rom[1009] = 25'b1111111111111111111111011;
    rom[1010] = 25'b1111111111111111111111011;
    rom[1011] = 25'b1111111111111111111111011;
    rom[1012] = 25'b1111111111111111111111011;
    rom[1013] = 25'b1111111111111111111111011;
    rom[1014] = 25'b1111111111111111111111011;
    rom[1015] = 25'b1111111111111111111111010;
    rom[1016] = 25'b1111111111111111111111010;
    rom[1017] = 25'b1111111111111111111111010;
    rom[1018] = 25'b1111111111111111111111010;
    rom[1019] = 25'b1111111111111111111111010;
    rom[1020] = 25'b1111111111111111111111010;
    rom[1021] = 25'b1111111111111111111111010;
    rom[1022] = 25'b1111111111111111111111010;
    rom[1023] = 25'b1111111111111111111111010;
    rom[1024] = 25'b1111111111111111111111010;
    rom[1025] = 25'b1111111111111111111111010;
    rom[1026] = 25'b1111111111111111111111010;
    rom[1027] = 25'b1111111111111111111111010;
    rom[1028] = 25'b1111111111111111111111010;
    rom[1029] = 25'b1111111111111111111111001;
    rom[1030] = 25'b1111111111111111111111001;
    rom[1031] = 25'b1111111111111111111111001;
    rom[1032] = 25'b1111111111111111111111001;
    rom[1033] = 25'b1111111111111111111111001;
    rom[1034] = 25'b1111111111111111111111001;
    rom[1035] = 25'b1111111111111111111111000;
    rom[1036] = 25'b1111111111111111111111000;
    rom[1037] = 25'b1111111111111111111111000;
    rom[1038] = 25'b1111111111111111111111000;
    rom[1039] = 25'b1111111111111111111111000;
    rom[1040] = 25'b1111111111111111111111000;
    rom[1041] = 25'b1111111111111111111110111;
    rom[1042] = 25'b1111111111111111111110111;
    rom[1043] = 25'b1111111111111111111110111;
    rom[1044] = 25'b1111111111111111111110111;
    rom[1045] = 25'b1111111111111111111110111;
    rom[1046] = 25'b1111111111111111111110111;
    rom[1047] = 25'b1111111111111111111110111;
    rom[1048] = 25'b1111111111111111111110110;
    rom[1049] = 25'b1111111111111111111110110;
    rom[1050] = 25'b1111111111111111111110110;
    rom[1051] = 25'b1111111111111111111110110;
    rom[1052] = 25'b1111111111111111111110110;
    rom[1053] = 25'b1111111111111111111110110;
    rom[1054] = 25'b1111111111111111111110101;
    rom[1055] = 25'b1111111111111111111110101;
    rom[1056] = 25'b1111111111111111111110101;
    rom[1057] = 25'b1111111111111111111110101;
    rom[1058] = 25'b1111111111111111111110101;
    rom[1059] = 25'b1111111111111111111110100;
    rom[1060] = 25'b1111111111111111111110100;
    rom[1061] = 25'b1111111111111111111110100;
    rom[1062] = 25'b1111111111111111111110100;
    rom[1063] = 25'b1111111111111111111110100;
    rom[1064] = 25'b1111111111111111111110100;
    rom[1065] = 25'b1111111111111111111110100;
    rom[1066] = 25'b1111111111111111111110100;
    rom[1067] = 25'b1111111111111111111110100;
    rom[1068] = 25'b1111111111111111111110100;
    rom[1069] = 25'b1111111111111111111110100;
    rom[1070] = 25'b1111111111111111111110100;
    rom[1071] = 25'b1111111111111111111110011;
    rom[1072] = 25'b1111111111111111111110011;
    rom[1073] = 25'b1111111111111111111110011;
    rom[1074] = 25'b1111111111111111111110011;
    rom[1075] = 25'b1111111111111111111110011;
    rom[1076] = 25'b1111111111111111111110011;
    rom[1077] = 25'b1111111111111111111110010;
    rom[1078] = 25'b1111111111111111111110010;
    rom[1079] = 25'b1111111111111111111110010;
    rom[1080] = 25'b1111111111111111111110010;
    rom[1081] = 25'b1111111111111111111110010;
    rom[1082] = 25'b1111111111111111111110001;
    rom[1083] = 25'b1111111111111111111110001;
    rom[1084] = 25'b1111111111111111111110001;
    rom[1085] = 25'b1111111111111111111110001;
    rom[1086] = 25'b1111111111111111111110001;
    rom[1087] = 25'b1111111111111111111110001;
    rom[1088] = 25'b1111111111111111111110000;
    rom[1089] = 25'b1111111111111111111110000;
    rom[1090] = 25'b1111111111111111111110000;
    rom[1091] = 25'b1111111111111111111110000;
    rom[1092] = 25'b1111111111111111111110000;
    rom[1093] = 25'b1111111111111111111101111;
    rom[1094] = 25'b1111111111111111111101111;
    rom[1095] = 25'b1111111111111111111101111;
    rom[1096] = 25'b1111111111111111111101111;
    rom[1097] = 25'b1111111111111111111101111;
    rom[1098] = 25'b1111111111111111111101110;
    rom[1099] = 25'b1111111111111111111101110;
    rom[1100] = 25'b1111111111111111111101110;
    rom[1101] = 25'b1111111111111111111101110;
    rom[1102] = 25'b1111111111111111111101110;
    rom[1103] = 25'b1111111111111111111101110;
    rom[1104] = 25'b1111111111111111111101110;
    rom[1105] = 25'b1111111111111111111101110;
    rom[1106] = 25'b1111111111111111111101110;
    rom[1107] = 25'b1111111111111111111101110;
    rom[1108] = 25'b1111111111111111111101110;
    rom[1109] = 25'b1111111111111111111101101;
    rom[1110] = 25'b1111111111111111111101101;
    rom[1111] = 25'b1111111111111111111101101;
    rom[1112] = 25'b1111111111111111111101101;
    rom[1113] = 25'b1111111111111111111101101;
    rom[1114] = 25'b1111111111111111111101100;
    rom[1115] = 25'b1111111111111111111101100;
    rom[1116] = 25'b1111111111111111111101100;
    rom[1117] = 25'b1111111111111111111101100;
    rom[1118] = 25'b1111111111111111111101100;
    rom[1119] = 25'b1111111111111111111101011;
    rom[1120] = 25'b1111111111111111111101011;
    rom[1121] = 25'b1111111111111111111101011;
    rom[1122] = 25'b1111111111111111111101011;
    rom[1123] = 25'b1111111111111111111101011;
    rom[1124] = 25'b1111111111111111111101010;
    rom[1125] = 25'b1111111111111111111101010;
    rom[1126] = 25'b1111111111111111111101010;
    rom[1127] = 25'b1111111111111111111101010;
    rom[1128] = 25'b1111111111111111111101010;
    rom[1129] = 25'b1111111111111111111101010;
    rom[1130] = 25'b1111111111111111111101001;
    rom[1131] = 25'b1111111111111111111101001;
    rom[1132] = 25'b1111111111111111111101001;
    rom[1133] = 25'b1111111111111111111101001;
    rom[1134] = 25'b1111111111111111111101001;
    rom[1135] = 25'b1111111111111111111101001;
    rom[1136] = 25'b1111111111111111111101001;
    rom[1137] = 25'b1111111111111111111101001;
    rom[1138] = 25'b1111111111111111111101001;
    rom[1139] = 25'b1111111111111111111101001;
    rom[1140] = 25'b1111111111111111111101000;
    rom[1141] = 25'b1111111111111111111101000;
    rom[1142] = 25'b1111111111111111111101000;
    rom[1143] = 25'b1111111111111111111101000;
    rom[1144] = 25'b1111111111111111111101000;
    rom[1145] = 25'b1111111111111111111100111;
    rom[1146] = 25'b1111111111111111111100111;
    rom[1147] = 25'b1111111111111111111100111;
    rom[1148] = 25'b1111111111111111111100111;
    rom[1149] = 25'b1111111111111111111100111;
    rom[1150] = 25'b1111111111111111111100110;
    rom[1151] = 25'b1111111111111111111100110;
    rom[1152] = 25'b1111111111111111111100110;
    rom[1153] = 25'b1111111111111111111100110;
    rom[1154] = 25'b1111111111111111111100110;
    rom[1155] = 25'b1111111111111111111100101;
    rom[1156] = 25'b1111111111111111111100101;
    rom[1157] = 25'b1111111111111111111100101;
    rom[1158] = 25'b1111111111111111111100101;
    rom[1159] = 25'b1111111111111111111100101;
    rom[1160] = 25'b1111111111111111111100100;
    rom[1161] = 25'b1111111111111111111100100;
    rom[1162] = 25'b1111111111111111111100100;
    rom[1163] = 25'b1111111111111111111100100;
    rom[1164] = 25'b1111111111111111111100100;
    rom[1165] = 25'b1111111111111111111100011;
    rom[1166] = 25'b1111111111111111111100011;
    rom[1167] = 25'b1111111111111111111100011;
    rom[1168] = 25'b1111111111111111111100011;
    rom[1169] = 25'b1111111111111111111100011;
    rom[1170] = 25'b1111111111111111111100011;
    rom[1171] = 25'b1111111111111111111100011;
    rom[1172] = 25'b1111111111111111111100011;
    rom[1173] = 25'b1111111111111111111100011;
    rom[1174] = 25'b1111111111111111111100011;
    rom[1175] = 25'b1111111111111111111100010;
    rom[1176] = 25'b1111111111111111111100010;
    rom[1177] = 25'b1111111111111111111100010;
    rom[1178] = 25'b1111111111111111111100010;
    rom[1179] = 25'b1111111111111111111100010;
    rom[1180] = 25'b1111111111111111111100001;
    rom[1181] = 25'b1111111111111111111100001;
    rom[1182] = 25'b1111111111111111111100001;
    rom[1183] = 25'b1111111111111111111100001;
    rom[1184] = 25'b1111111111111111111100001;
    rom[1185] = 25'b1111111111111111111100000;
    rom[1186] = 25'b1111111111111111111100000;
    rom[1187] = 25'b1111111111111111111100000;
    rom[1188] = 25'b1111111111111111111100000;
    rom[1189] = 25'b1111111111111111111100000;
    rom[1190] = 25'b1111111111111111111011111;
    rom[1191] = 25'b1111111111111111111011111;
    rom[1192] = 25'b1111111111111111111011111;
    rom[1193] = 25'b1111111111111111111011111;
    rom[1194] = 25'b1111111111111111111011111;
    rom[1195] = 25'b1111111111111111111011110;
    rom[1196] = 25'b1111111111111111111011110;
    rom[1197] = 25'b1111111111111111111011110;
    rom[1198] = 25'b1111111111111111111011110;
    rom[1199] = 25'b1111111111111111111011110;
    rom[1200] = 25'b1111111111111111111011101;
    rom[1201] = 25'b1111111111111111111011101;
    rom[1202] = 25'b1111111111111111111011101;
    rom[1203] = 25'b1111111111111111111011101;
    rom[1204] = 25'b1111111111111111111011101;
    rom[1205] = 25'b1111111111111111111011101;
    rom[1206] = 25'b1111111111111111111011101;
    rom[1207] = 25'b1111111111111111111011101;
    rom[1208] = 25'b1111111111111111111011101;
    rom[1209] = 25'b1111111111111111111011101;
    rom[1210] = 25'b1111111111111111111011101;
    rom[1211] = 25'b1111111111111111111011100;
    rom[1212] = 25'b1111111111111111111011100;
    rom[1213] = 25'b1111111111111111111011100;
    rom[1214] = 25'b1111111111111111111011100;
    rom[1215] = 25'b1111111111111111111011100;
    rom[1216] = 25'b1111111111111111111011011;
    rom[1217] = 25'b1111111111111111111011011;
    rom[1218] = 25'b1111111111111111111011011;
    rom[1219] = 25'b1111111111111111111011011;
    rom[1220] = 25'b1111111111111111111011011;
    rom[1221] = 25'b1111111111111111111011011;
    rom[1222] = 25'b1111111111111111111011010;
    rom[1223] = 25'b1111111111111111111011010;
    rom[1224] = 25'b1111111111111111111011010;
    rom[1225] = 25'b1111111111111111111011010;
    rom[1226] = 25'b1111111111111111111011010;
    rom[1227] = 25'b1111111111111111111011001;
    rom[1228] = 25'b1111111111111111111011001;
    rom[1229] = 25'b1111111111111111111011001;
    rom[1230] = 25'b1111111111111111111011001;
    rom[1231] = 25'b1111111111111111111011001;
    rom[1232] = 25'b1111111111111111111011001;
    rom[1233] = 25'b1111111111111111111011000;
    rom[1234] = 25'b1111111111111111111011000;
    rom[1235] = 25'b1111111111111111111011000;
    rom[1236] = 25'b1111111111111111111011000;
    rom[1237] = 25'b1111111111111111111011000;
    rom[1238] = 25'b1111111111111111111011000;
    rom[1239] = 25'b1111111111111111111011000;
    rom[1240] = 25'b1111111111111111111011000;
    rom[1241] = 25'b1111111111111111111011000;
    rom[1242] = 25'b1111111111111111111011000;
    rom[1243] = 25'b1111111111111111111011000;
    rom[1244] = 25'b1111111111111111111011000;
    rom[1245] = 25'b1111111111111111111010111;
    rom[1246] = 25'b1111111111111111111010111;
    rom[1247] = 25'b1111111111111111111010111;
    rom[1248] = 25'b1111111111111111111010111;
    rom[1249] = 25'b1111111111111111111010111;
    rom[1250] = 25'b1111111111111111111010111;
    rom[1251] = 25'b1111111111111111111010110;
    rom[1252] = 25'b1111111111111111111010110;
    rom[1253] = 25'b1111111111111111111010110;
    rom[1254] = 25'b1111111111111111111010110;
    rom[1255] = 25'b1111111111111111111010110;
    rom[1256] = 25'b1111111111111111111010110;
    rom[1257] = 25'b1111111111111111111010101;
    rom[1258] = 25'b1111111111111111111010101;
    rom[1259] = 25'b1111111111111111111010101;
    rom[1260] = 25'b1111111111111111111010101;
    rom[1261] = 25'b1111111111111111111010101;
    rom[1262] = 25'b1111111111111111111010101;
    rom[1263] = 25'b1111111111111111111010100;
    rom[1264] = 25'b1111111111111111111010100;
    rom[1265] = 25'b1111111111111111111010100;
    rom[1266] = 25'b1111111111111111111010100;
    rom[1267] = 25'b1111111111111111111010100;
    rom[1268] = 25'b1111111111111111111010100;
    rom[1269] = 25'b1111111111111111111010100;
    rom[1270] = 25'b1111111111111111111010011;
    rom[1271] = 25'b1111111111111111111010011;
    rom[1272] = 25'b1111111111111111111010011;
    rom[1273] = 25'b1111111111111111111010011;
    rom[1274] = 25'b1111111111111111111010011;
    rom[1275] = 25'b1111111111111111111010011;
    rom[1276] = 25'b1111111111111111111010011;
    rom[1277] = 25'b1111111111111111111010010;
    rom[1278] = 25'b1111111111111111111010010;
    rom[1279] = 25'b1111111111111111111010010;
    rom[1280] = 25'b1111111111111111111010010;
    rom[1281] = 25'b1111111111111111111010010;
    rom[1282] = 25'b1111111111111111111010010;
    rom[1283] = 25'b1111111111111111111010010;
    rom[1284] = 25'b1111111111111111111010010;
    rom[1285] = 25'b1111111111111111111010010;
    rom[1286] = 25'b1111111111111111111010010;
    rom[1287] = 25'b1111111111111111111010010;
    rom[1288] = 25'b1111111111111111111010010;
    rom[1289] = 25'b1111111111111111111010010;
    rom[1290] = 25'b1111111111111111111010010;
    rom[1291] = 25'b1111111111111111111010010;
    rom[1292] = 25'b1111111111111111111010010;
    rom[1293] = 25'b1111111111111111111010001;
    rom[1294] = 25'b1111111111111111111010001;
    rom[1295] = 25'b1111111111111111111010001;
    rom[1296] = 25'b1111111111111111111010001;
    rom[1297] = 25'b1111111111111111111010001;
    rom[1298] = 25'b1111111111111111111010001;
    rom[1299] = 25'b1111111111111111111010001;
    rom[1300] = 25'b1111111111111111111010001;
    rom[1301] = 25'b1111111111111111111010001;
    rom[1302] = 25'b1111111111111111111010000;
    rom[1303] = 25'b1111111111111111111010000;
    rom[1304] = 25'b1111111111111111111010000;
    rom[1305] = 25'b1111111111111111111010000;
    rom[1306] = 25'b1111111111111111111010000;
    rom[1307] = 25'b1111111111111111111010000;
    rom[1308] = 25'b1111111111111111111010000;
    rom[1309] = 25'b1111111111111111111010000;
    rom[1310] = 25'b1111111111111111111010000;
    rom[1311] = 25'b1111111111111111111010000;
    rom[1312] = 25'b1111111111111111111001111;
    rom[1313] = 25'b1111111111111111111001111;
    rom[1314] = 25'b1111111111111111111001111;
    rom[1315] = 25'b1111111111111111111001111;
    rom[1316] = 25'b1111111111111111111001111;
    rom[1317] = 25'b1111111111111111111001111;
    rom[1318] = 25'b1111111111111111111001111;
    rom[1319] = 25'b1111111111111111111001111;
    rom[1320] = 25'b1111111111111111111001111;
    rom[1321] = 25'b1111111111111111111001111;
    rom[1322] = 25'b1111111111111111111001111;
    rom[1323] = 25'b1111111111111111111001111;
    rom[1324] = 25'b1111111111111111111001110;
    rom[1325] = 25'b1111111111111111111001110;
    rom[1326] = 25'b1111111111111111111001110;
    rom[1327] = 25'b1111111111111111111001110;
    rom[1328] = 25'b1111111111111111111001110;
    rom[1329] = 25'b1111111111111111111001110;
    rom[1330] = 25'b1111111111111111111001110;
    rom[1331] = 25'b1111111111111111111001110;
    rom[1332] = 25'b1111111111111111111001110;
    rom[1333] = 25'b1111111111111111111001110;
    rom[1334] = 25'b1111111111111111111001110;
    rom[1335] = 25'b1111111111111111111001110;
    rom[1336] = 25'b1111111111111111111001110;
    rom[1337] = 25'b1111111111111111111001110;
    rom[1338] = 25'b1111111111111111111001110;
    rom[1339] = 25'b1111111111111111111001110;
    rom[1340] = 25'b1111111111111111111001110;
    rom[1341] = 25'b1111111111111111111001110;
    rom[1342] = 25'b1111111111111111111001101;
    rom[1343] = 25'b1111111111111111111001101;
    rom[1344] = 25'b1111111111111111111001101;
    rom[1345] = 25'b1111111111111111111001101;
    rom[1346] = 25'b1111111111111111111001101;
    rom[1347] = 25'b1111111111111111111001101;
    rom[1348] = 25'b1111111111111111111001101;
    rom[1349] = 25'b1111111111111111111001101;
    rom[1350] = 25'b1111111111111111111001101;
    rom[1351] = 25'b1111111111111111111001101;
    rom[1352] = 25'b1111111111111111111001101;
    rom[1353] = 25'b1111111111111111111001101;
    rom[1354] = 25'b1111111111111111111001101;
    rom[1355] = 25'b1111111111111111111001101;
    rom[1356] = 25'b1111111111111111111001101;
    rom[1357] = 25'b1111111111111111111001101;
    rom[1358] = 25'b1111111111111111111001101;
    rom[1359] = 25'b1111111111111111111001101;
    rom[1360] = 25'b1111111111111111111001101;
    rom[1361] = 25'b1111111111111111111001101;
    rom[1362] = 25'b1111111111111111111001101;
    rom[1363] = 25'b1111111111111111111001101;
    rom[1364] = 25'b1111111111111111111001101;
    rom[1365] = 25'b1111111111111111111001101;
    rom[1366] = 25'b1111111111111111111001101;
    rom[1367] = 25'b1111111111111111111001101;
    rom[1368] = 25'b1111111111111111111001101;
    rom[1369] = 25'b1111111111111111111001101;
    rom[1370] = 25'b1111111111111111111001101;
    rom[1371] = 25'b1111111111111111111001101;
    rom[1372] = 25'b1111111111111111111001101;
    rom[1373] = 25'b1111111111111111111001101;
    rom[1374] = 25'b1111111111111111111001101;
    rom[1375] = 25'b1111111111111111111001101;
    rom[1376] = 25'b1111111111111111111001101;
    rom[1377] = 25'b1111111111111111111001101;
    rom[1378] = 25'b1111111111111111111001101;
    rom[1379] = 25'b1111111111111111111001101;
    rom[1380] = 25'b1111111111111111111001101;
    rom[1381] = 25'b1111111111111111111001101;
    rom[1382] = 25'b1111111111111111111001101;
    rom[1383] = 25'b1111111111111111111001110;
    rom[1384] = 25'b1111111111111111111001110;
    rom[1385] = 25'b1111111111111111111001110;
    rom[1386] = 25'b1111111111111111111001110;
    rom[1387] = 25'b1111111111111111111001110;
    rom[1388] = 25'b1111111111111111111001110;
    rom[1389] = 25'b1111111111111111111001110;
    rom[1390] = 25'b1111111111111111111001110;
    rom[1391] = 25'b1111111111111111111001110;
    rom[1392] = 25'b1111111111111111111001110;
    rom[1393] = 25'b1111111111111111111001110;
    rom[1394] = 25'b1111111111111111111001110;
    rom[1395] = 25'b1111111111111111111001110;
    rom[1396] = 25'b1111111111111111111001110;
    rom[1397] = 25'b1111111111111111111001110;
    rom[1398] = 25'b1111111111111111111001110;
    rom[1399] = 25'b1111111111111111111001111;
    rom[1400] = 25'b1111111111111111111001111;
    rom[1401] = 25'b1111111111111111111001111;
    rom[1402] = 25'b1111111111111111111001111;
    rom[1403] = 25'b1111111111111111111001111;
    rom[1404] = 25'b1111111111111111111001111;
    rom[1405] = 25'b1111111111111111111001111;
    rom[1406] = 25'b1111111111111111111001111;
    rom[1407] = 25'b1111111111111111111001111;
    rom[1408] = 25'b1111111111111111111001111;
    rom[1409] = 25'b1111111111111111111010000;
    rom[1410] = 25'b1111111111111111111010000;
    rom[1411] = 25'b1111111111111111111010000;
    rom[1412] = 25'b1111111111111111111010000;
    rom[1413] = 25'b1111111111111111111010000;
    rom[1414] = 25'b1111111111111111111010000;
    rom[1415] = 25'b1111111111111111111010000;
    rom[1416] = 25'b1111111111111111111010000;
    rom[1417] = 25'b1111111111111111111010001;
    rom[1418] = 25'b1111111111111111111010001;
    rom[1419] = 25'b1111111111111111111010001;
    rom[1420] = 25'b1111111111111111111010001;
    rom[1421] = 25'b1111111111111111111010001;
    rom[1422] = 25'b1111111111111111111010001;
    rom[1423] = 25'b1111111111111111111010001;
    rom[1424] = 25'b1111111111111111111010010;
    rom[1425] = 25'b1111111111111111111010010;
    rom[1426] = 25'b1111111111111111111010010;
    rom[1427] = 25'b1111111111111111111010010;
    rom[1428] = 25'b1111111111111111111010010;
    rom[1429] = 25'b1111111111111111111010010;
    rom[1430] = 25'b1111111111111111111010010;
    rom[1431] = 25'b1111111111111111111010010;
    rom[1432] = 25'b1111111111111111111010010;
    rom[1433] = 25'b1111111111111111111010010;
    rom[1434] = 25'b1111111111111111111010010;
    rom[1435] = 25'b1111111111111111111010010;
    rom[1436] = 25'b1111111111111111111010011;
    rom[1437] = 25'b1111111111111111111010011;
    rom[1438] = 25'b1111111111111111111010011;
    rom[1439] = 25'b1111111111111111111010011;
    rom[1440] = 25'b1111111111111111111010011;
    rom[1441] = 25'b1111111111111111111010011;
    rom[1442] = 25'b1111111111111111111010100;
    rom[1443] = 25'b1111111111111111111010100;
    rom[1444] = 25'b1111111111111111111010100;
    rom[1445] = 25'b1111111111111111111010100;
    rom[1446] = 25'b1111111111111111111010100;
    rom[1447] = 25'b1111111111111111111010101;
    rom[1448] = 25'b1111111111111111111010101;
    rom[1449] = 25'b1111111111111111111010101;
    rom[1450] = 25'b1111111111111111111010101;
    rom[1451] = 25'b1111111111111111111010110;
    rom[1452] = 25'b1111111111111111111010110;
    rom[1453] = 25'b1111111111111111111010110;
    rom[1454] = 25'b1111111111111111111010110;
    rom[1455] = 25'b1111111111111111111010111;
    rom[1456] = 25'b1111111111111111111010111;
    rom[1457] = 25'b1111111111111111111010111;
    rom[1458] = 25'b1111111111111111111010111;
    rom[1459] = 25'b1111111111111111111011000;
    rom[1460] = 25'b1111111111111111111011000;
    rom[1461] = 25'b1111111111111111111011000;
    rom[1462] = 25'b1111111111111111111011000;
    rom[1463] = 25'b1111111111111111111011000;
    rom[1464] = 25'b1111111111111111111011000;
    rom[1465] = 25'b1111111111111111111011000;
    rom[1466] = 25'b1111111111111111111011000;
    rom[1467] = 25'b1111111111111111111011001;
    rom[1468] = 25'b1111111111111111111011001;
    rom[1469] = 25'b1111111111111111111011001;
    rom[1470] = 25'b1111111111111111111011001;
    rom[1471] = 25'b1111111111111111111011010;
    rom[1472] = 25'b1111111111111111111011010;
    rom[1473] = 25'b1111111111111111111011010;
    rom[1474] = 25'b1111111111111111111011011;
    rom[1475] = 25'b1111111111111111111011011;
    rom[1476] = 25'b1111111111111111111011011;
    rom[1477] = 25'b1111111111111111111011100;
    rom[1478] = 25'b1111111111111111111011100;
    rom[1479] = 25'b1111111111111111111011100;
    rom[1480] = 25'b1111111111111111111011100;
    rom[1481] = 25'b1111111111111111111011101;
    rom[1482] = 25'b1111111111111111111011101;
    rom[1483] = 25'b1111111111111111111011101;
    rom[1484] = 25'b1111111111111111111011101;
    rom[1485] = 25'b1111111111111111111011101;
    rom[1486] = 25'b1111111111111111111011101;
    rom[1487] = 25'b1111111111111111111011110;
    rom[1488] = 25'b1111111111111111111011110;
    rom[1489] = 25'b1111111111111111111011110;
    rom[1490] = 25'b1111111111111111111011111;
    rom[1491] = 25'b1111111111111111111011111;
    rom[1492] = 25'b1111111111111111111100000;
    rom[1493] = 25'b1111111111111111111100000;
    rom[1494] = 25'b1111111111111111111100000;
    rom[1495] = 25'b1111111111111111111100001;
    rom[1496] = 25'b1111111111111111111100001;
    rom[1497] = 25'b1111111111111111111100001;
    rom[1498] = 25'b1111111111111111111100010;
    rom[1499] = 25'b1111111111111111111100010;
    rom[1500] = 25'b1111111111111111111100010;
    rom[1501] = 25'b1111111111111111111100011;
    rom[1502] = 25'b1111111111111111111100011;
    rom[1503] = 25'b1111111111111111111100011;
    rom[1504] = 25'b1111111111111111111100011;
    rom[1505] = 25'b1111111111111111111100011;
    rom[1506] = 25'b1111111111111111111100100;
    rom[1507] = 25'b1111111111111111111100100;
    rom[1508] = 25'b1111111111111111111100101;
    rom[1509] = 25'b1111111111111111111100101;
    rom[1510] = 25'b1111111111111111111100101;
    rom[1511] = 25'b1111111111111111111100110;
    rom[1512] = 25'b1111111111111111111100110;
    rom[1513] = 25'b1111111111111111111100111;
    rom[1514] = 25'b1111111111111111111100111;
    rom[1515] = 25'b1111111111111111111101000;
    rom[1516] = 25'b1111111111111111111101000;
    rom[1517] = 25'b1111111111111111111101000;
    rom[1518] = 25'b1111111111111111111101001;
    rom[1519] = 25'b1111111111111111111101001;
    rom[1520] = 25'b1111111111111111111101001;
    rom[1521] = 25'b1111111111111111111101001;
    rom[1522] = 25'b1111111111111111111101010;
    rom[1523] = 25'b1111111111111111111101010;
    rom[1524] = 25'b1111111111111111111101011;
    rom[1525] = 25'b1111111111111111111101011;
    rom[1526] = 25'b1111111111111111111101100;
    rom[1527] = 25'b1111111111111111111101100;
    rom[1528] = 25'b1111111111111111111101100;
    rom[1529] = 25'b1111111111111111111101101;
    rom[1530] = 25'b1111111111111111111101101;
    rom[1531] = 25'b1111111111111111111101110;
    rom[1532] = 25'b1111111111111111111101110;
    rom[1533] = 25'b1111111111111111111101110;
    rom[1534] = 25'b1111111111111111111101110;
    rom[1535] = 25'b1111111111111111111101111;
    rom[1536] = 25'b1111111111111111111101111;
    rom[1537] = 25'b1111111111111111111110000;
    rom[1538] = 25'b1111111111111111111110000;
    rom[1539] = 25'b1111111111111111111110001;
    rom[1540] = 25'b1111111111111111111110001;
    rom[1541] = 25'b1111111111111111111110010;
    rom[1542] = 25'b1111111111111111111110010;
    rom[1543] = 25'b1111111111111111111110011;
    rom[1544] = 25'b1111111111111111111110100;
    rom[1545] = 25'b1111111111111111111110100;
    rom[1546] = 25'b1111111111111111111110100;
    rom[1547] = 25'b1111111111111111111110100;
    rom[1548] = 25'b1111111111111111111110101;
    rom[1549] = 25'b1111111111111111111110101;
    rom[1550] = 25'b1111111111111111111110110;
    rom[1551] = 25'b1111111111111111111110110;
    rom[1552] = 25'b1111111111111111111110111;
    rom[1553] = 25'b1111111111111111111110111;
    rom[1554] = 25'b1111111111111111111111000;
    rom[1555] = 25'b1111111111111111111111001;
    rom[1556] = 25'b1111111111111111111111001;
    rom[1557] = 25'b1111111111111111111111010;
    rom[1558] = 25'b1111111111111111111111010;
    rom[1559] = 25'b1111111111111111111111010;
    rom[1560] = 25'b1111111111111111111111010;
    rom[1561] = 25'b1111111111111111111111011;
    rom[1562] = 25'b1111111111111111111111100;
    rom[1563] = 25'b1111111111111111111111100;
    rom[1564] = 25'b1111111111111111111111101;
    rom[1565] = 25'b1111111111111111111111101;
    rom[1566] = 25'b1111111111111111111111110;
    rom[1567] = 25'b1111111111111111111111111;
    rom[1568] = 25'b1111111111111111111111111;
    rom[1569] = 25'b0000000000000000000000000;
    rom[1570] = 25'b0000000000000000000000000;
    rom[1571] = 25'b0000000000000000000000000;
    rom[1572] = 25'b0000000000000000000000000;
    rom[1573] = 25'b0000000000000000000000000;
    rom[1574] = 25'b0000000000000000000000001;
    rom[1575] = 25'b0000000000000000000000001;
    rom[1576] = 25'b0000000000000000000000010;
    rom[1577] = 25'b0000000000000000000000011;
    rom[1578] = 25'b0000000000000000000000011;
    rom[1579] = 25'b0000000000000000000000100;
    rom[1580] = 25'b0000000000000000000000101;
    rom[1581] = 25'b0000000000000000000000101;
    rom[1582] = 25'b0000000000000000000000101;
    rom[1583] = 25'b0000000000000000000000110;
    rom[1584] = 25'b0000000000000000000000110;
    rom[1585] = 25'b0000000000000000000000111;
    rom[1586] = 25'b0000000000000000000001000;
    rom[1587] = 25'b0000000000000000000001000;
    rom[1588] = 25'b0000000000000000000001001;
    rom[1589] = 25'b0000000000000000000001010;
    rom[1590] = 25'b0000000000000000000001010;
    rom[1591] = 25'b0000000000000000000001011;
    rom[1592] = 25'b0000000000000000000001011;
    rom[1593] = 25'b0000000000000000000001011;
    rom[1594] = 25'b0000000000000000000001100;
    rom[1595] = 25'b0000000000000000000001101;
    rom[1596] = 25'b0000000000000000000001101;
    rom[1597] = 25'b0000000000000000000001110;
    rom[1598] = 25'b0000000000000000000001111;
    rom[1599] = 25'b0000000000000000000010000;
    rom[1600] = 25'b0000000000000000000010000;
    rom[1601] = 25'b0000000000000000000010001;
    rom[1602] = 25'b0000000000000000000010001;
    rom[1603] = 25'b0000000000000000000010001;
    rom[1604] = 25'b0000000000000000000010010;
    rom[1605] = 25'b0000000000000000000010011;
    rom[1606] = 25'b0000000000000000000010100;
    rom[1607] = 25'b0000000000000000000010100;
    rom[1608] = 25'b0000000000000000000010101;
    rom[1609] = 25'b0000000000000000000010110;
    rom[1610] = 25'b0000000000000000000010110;
    rom[1611] = 25'b0000000000000000000010110;
    rom[1612] = 25'b0000000000000000000010111;
    rom[1613] = 25'b0000000000000000000011000;
    rom[1614] = 25'b0000000000000000000011001;
    rom[1615] = 25'b0000000000000000000011001;
    rom[1616] = 25'b0000000000000000000011010;
    rom[1617] = 25'b0000000000000000000011011;
    rom[1618] = 25'b0000000000000000000011100;
    rom[1619] = 25'b0000000000000000000011100;
    rom[1620] = 25'b0000000000000000000011100;
    rom[1621] = 25'b0000000000000000000011101;
    rom[1622] = 25'b0000000000000000000011110;
    rom[1623] = 25'b0000000000000000000011110;
    rom[1624] = 25'b0000000000000000000011111;
    rom[1625] = 25'b0000000000000000000100000;
    rom[1626] = 25'b0000000000000000000100001;
    rom[1627] = 25'b0000000000000000000100010;
    rom[1628] = 25'b0000000000000000000100010;
    rom[1629] = 25'b0000000000000000000100010;
    rom[1630] = 25'b0000000000000000000100011;
    rom[1631] = 25'b0000000000000000000100100;
    rom[1632] = 25'b0000000000000000000100101;
    rom[1633] = 25'b0000000000000000000100101;
    rom[1634] = 25'b0000000000000000000100110;
    rom[1635] = 25'b0000000000000000000100111;
    rom[1636] = 25'b0000000000000000000100111;
    rom[1637] = 25'b0000000000000000000101000;
    rom[1638] = 25'b0000000000000000000101000;
    rom[1639] = 25'b0000000000000000000101001;
    rom[1640] = 25'b0000000000000000000101010;
    rom[1641] = 25'b0000000000000000000101011;
    rom[1642] = 25'b0000000000000000000101100;
    rom[1643] = 25'b0000000000000000000101101;
    rom[1644] = 25'b0000000000000000000101101;
    rom[1645] = 25'b0000000000000000000101101;
    rom[1646] = 25'b0000000000000000000101110;
    rom[1647] = 25'b0000000000000000000101111;
    rom[1648] = 25'b0000000000000000000110000;
    rom[1649] = 25'b0000000000000000000110001;
    rom[1650] = 25'b0000000000000000000110001;
    rom[1651] = 25'b0000000000000000000110010;
    rom[1652] = 25'b0000000000000000000110011;
    rom[1653] = 25'b0000000000000000000110011;
    rom[1654] = 25'b0000000000000000000110100;
    rom[1655] = 25'b0000000000000000000110101;
    rom[1656] = 25'b0000000000000000000110110;
    rom[1657] = 25'b0000000000000000000110111;
    rom[1658] = 25'b0000000000000000000110111;
    rom[1659] = 25'b0000000000000000000111000;
    rom[1660] = 25'b0000000000000000000111000;
    rom[1661] = 25'b0000000000000000000111001;
    rom[1662] = 25'b0000000000000000000111010;
    rom[1663] = 25'b0000000000000000000111011;
    rom[1664] = 25'b0000000000000000000111100;
    rom[1665] = 25'b0000000000000000000111101;
    rom[1666] = 25'b0000000000000000000111101;
    rom[1667] = 25'b0000000000000000000111110;
    rom[1668] = 25'b0000000000000000000111110;
    rom[1669] = 25'b0000000000000000000111111;
    rom[1670] = 25'b0000000000000000001000000;
    rom[1671] = 25'b0000000000000000001000001;
    rom[1672] = 25'b0000000000000000001000010;
    rom[1673] = 25'b0000000000000000001000011;
    rom[1674] = 25'b0000000000000000001000100;
    rom[1675] = 25'b0000000000000000001000100;
    rom[1676] = 25'b0000000000000000001000100;
    rom[1677] = 25'b0000000000000000001000101;
    rom[1678] = 25'b0000000000000000001000110;
    rom[1679] = 25'b0000000000000000001000111;
    rom[1680] = 25'b0000000000000000001001000;
    rom[1681] = 25'b0000000000000000001001001;
    rom[1682] = 25'b0000000000000000001001001;
    rom[1683] = 25'b0000000000000000001001010;
    rom[1684] = 25'b0000000000000000001001011;
    rom[1685] = 25'b0000000000000000001001100;
    rom[1686] = 25'b0000000000000000001001101;
    rom[1687] = 25'b0000000000000000001001110;
    rom[1688] = 25'b0000000000000000001001110;
    rom[1689] = 25'b0000000000000000001001111;
    rom[1690] = 25'b0000000000000000001001111;
    rom[1691] = 25'b0000000000000000001010000;
    rom[1692] = 25'b0000000000000000001010001;
    rom[1693] = 25'b0000000000000000001010010;
    rom[1694] = 25'b0000000000000000001010011;
    rom[1695] = 25'b0000000000000000001010100;
    rom[1696] = 25'b0000000000000000001010101;
    rom[1697] = 25'b0000000000000000001010101;
    rom[1698] = 25'b0000000000000000001010110;
    rom[1699] = 25'b0000000000000000001010111;
    rom[1700] = 25'b0000000000000000001011000;
    rom[1701] = 25'b0000000000000000001011001;
    rom[1702] = 25'b0000000000000000001011010;
    rom[1703] = 25'b0000000000000000001011011;
    rom[1704] = 25'b0000000000000000001011011;
    rom[1705] = 25'b0000000000000000001011011;
    rom[1706] = 25'b0000000000000000001011100;
    rom[1707] = 25'b0000000000000000001011101;
    rom[1708] = 25'b0000000000000000001011110;
    rom[1709] = 25'b0000000000000000001011111;
    rom[1710] = 25'b0000000000000000001100000;
    rom[1711] = 25'b0000000000000000001100000;
    rom[1712] = 25'b0000000000000000001100001;
    rom[1713] = 25'b0000000000000000001100010;
    rom[1714] = 25'b0000000000000000001100011;
    rom[1715] = 25'b0000000000000000001100100;
    rom[1716] = 25'b0000000000000000001100101;
    rom[1717] = 25'b0000000000000000001100110;
    rom[1718] = 25'b0000000000000000001100110;
    rom[1719] = 25'b0000000000000000001100111;
    rom[1720] = 25'b0000000000000000001101000;
    rom[1721] = 25'b0000000000000000001101001;
    rom[1722] = 25'b0000000000000000001101010;
    rom[1723] = 25'b0000000000000000001101011;
    rom[1724] = 25'b0000000000000000001101100;
    rom[1725] = 25'b0000000000000000001101100;
    rom[1726] = 25'b0000000000000000001101101;
    rom[1727] = 25'b0000000000000000001101110;
    rom[1728] = 25'b0000000000000000001101111;
    rom[1729] = 25'b0000000000000000001110000;
    rom[1730] = 25'b0000000000000000001110001;
    rom[1731] = 25'b0000000000000000001110001;
    rom[1732] = 25'b0000000000000000001110010;
    rom[1733] = 25'b0000000000000000001110011;
    rom[1734] = 25'b0000000000000000001110100;
    rom[1735] = 25'b0000000000000000001110101;
    rom[1736] = 25'b0000000000000000001110110;
    rom[1737] = 25'b0000000000000000001110111;
    rom[1738] = 25'b0000000000000000001110111;
    rom[1739] = 25'b0000000000000000001111000;
    rom[1740] = 25'b0000000000000000001111000;
    rom[1741] = 25'b0000000000000000001111001;
    rom[1742] = 25'b0000000000000000001111010;
    rom[1743] = 25'b0000000000000000001111011;
    rom[1744] = 25'b0000000000000000001111100;
    rom[1745] = 25'b0000000000000000001111101;
    rom[1746] = 25'b0000000000000000001111101;
    rom[1747] = 25'b0000000000000000001111110;
    rom[1748] = 25'b0000000000000000001111111;
    rom[1749] = 25'b0000000000000000010000000;
    rom[1750] = 25'b0000000000000000010000001;
    rom[1751] = 25'b0000000000000000010000010;
    rom[1752] = 25'b0000000000000000010000010;
    rom[1753] = 25'b0000000000000000010000011;
    rom[1754] = 25'b0000000000000000010000100;
    rom[1755] = 25'b0000000000000000010000101;
    rom[1756] = 25'b0000000000000000010000110;
    rom[1757] = 25'b0000000000000000010000111;
    rom[1758] = 25'b0000000000000000010001000;
    rom[1759] = 25'b0000000000000000010001000;
    rom[1760] = 25'b0000000000000000010001001;
    rom[1761] = 25'b0000000000000000010001010;
    rom[1762] = 25'b0000000000000000010001011;
    rom[1763] = 25'b0000000000000000010001100;
    rom[1764] = 25'b0000000000000000010001101;
    rom[1765] = 25'b0000000000000000010001110;
    rom[1766] = 25'b0000000000000000010001110;
    rom[1767] = 25'b0000000000000000010001111;
    rom[1768] = 25'b0000000000000000010010000;
    rom[1769] = 25'b0000000000000000010010001;
    rom[1770] = 25'b0000000000000000010010010;
    rom[1771] = 25'b0000000000000000010010011;
    rom[1772] = 25'b0000000000000000010010011;
    rom[1773] = 25'b0000000000000000010010100;
    rom[1774] = 25'b0000000000000000010010101;
    rom[1775] = 25'b0000000000000000010010110;
    rom[1776] = 25'b0000000000000000010010111;
    rom[1777] = 25'b0000000000000000010011000;
    rom[1778] = 25'b0000000000000000010011001;
    rom[1779] = 25'b0000000000000000010011001;
    rom[1780] = 25'b0000000000000000010011010;
    rom[1781] = 25'b0000000000000000010011010;
    rom[1782] = 25'b0000000000000000010011011;
    rom[1783] = 25'b0000000000000000010011100;
    rom[1784] = 25'b0000000000000000010011101;
    rom[1785] = 25'b0000000000000000010011110;
    rom[1786] = 25'b0000000000000000010011111;
    rom[1787] = 25'b0000000000000000010011111;
    rom[1788] = 25'b0000000000000000010100000;
    rom[1789] = 25'b0000000000000000010100001;
    rom[1790] = 25'b0000000000000000010100010;
    rom[1791] = 25'b0000000000000000010100011;
    rom[1792] = 25'b0000000000000000010100100;
    rom[1793] = 25'b0000000000000000010100100;
    rom[1794] = 25'b0000000000000000010100101;
    rom[1795] = 25'b0000000000000000010100110;
    rom[1796] = 25'b0000000000000000010100111;
    rom[1797] = 25'b0000000000000000010101000;
    rom[1798] = 25'b0000000000000000010101001;
    rom[1799] = 25'b0000000000000000010101010;
    rom[1800] = 25'b0000000000000000010101010;
    rom[1801] = 25'b0000000000000000010101010;
    rom[1802] = 25'b0000000000000000010101011;
    rom[1803] = 25'b0000000000000000010101100;
    rom[1804] = 25'b0000000000000000010101101;
    rom[1805] = 25'b0000000000000000010101110;
    rom[1806] = 25'b0000000000000000010101111;
    rom[1807] = 25'b0000000000000000010110000;
    rom[1808] = 25'b0000000000000000010110000;
    rom[1809] = 25'b0000000000000000010110001;
    rom[1810] = 25'b0000000000000000010110010;
    rom[1811] = 25'b0000000000000000010110011;
    rom[1812] = 25'b0000000000000000010110011;
    rom[1813] = 25'b0000000000000000010110100;
    rom[1814] = 25'b0000000000000000010110101;
    rom[1815] = 25'b0000000000000000010110110;
    rom[1816] = 25'b0000000000000000010110110;
    rom[1817] = 25'b0000000000000000010110111;
    rom[1818] = 25'b0000000000000000010111000;
    rom[1819] = 25'b0000000000000000010111001;
    rom[1820] = 25'b0000000000000000010111010;
    rom[1821] = 25'b0000000000000000010111010;
    rom[1822] = 25'b0000000000000000010111011;
    rom[1823] = 25'b0000000000000000010111011;
    rom[1824] = 25'b0000000000000000010111100;
    rom[1825] = 25'b0000000000000000010111101;
    rom[1826] = 25'b0000000000000000010111110;
    rom[1827] = 25'b0000000000000000010111111;
    rom[1828] = 25'b0000000000000000010111111;
    rom[1829] = 25'b0000000000000000011000000;
    rom[1830] = 25'b0000000000000000011000001;
    rom[1831] = 25'b0000000000000000011000001;
    rom[1832] = 25'b0000000000000000011000010;
    rom[1833] = 25'b0000000000000000011000011;
    rom[1834] = 25'b0000000000000000011000011;
    rom[1835] = 25'b0000000000000000011000100;
    rom[1836] = 25'b0000000000000000011000101;
    rom[1837] = 25'b0000000000000000011000110;
    rom[1838] = 25'b0000000000000000011000111;
    rom[1839] = 25'b0000000000000000011000111;
    rom[1840] = 25'b0000000000000000011000111;
    rom[1841] = 25'b0000000000000000011001000;
    rom[1842] = 25'b0000000000000000011001001;
    rom[1843] = 25'b0000000000000000011001010;
    rom[1844] = 25'b0000000000000000011001011;
    rom[1845] = 25'b0000000000000000011001011;
    rom[1846] = 25'b0000000000000000011001100;
    rom[1847] = 25'b0000000000000000011001100;
    rom[1848] = 25'b0000000000000000011001101;
    rom[1849] = 25'b0000000000000000011001101;
    rom[1850] = 25'b0000000000000000011001110;
    rom[1851] = 25'b0000000000000000011001111;
    rom[1852] = 25'b0000000000000000011010000;
    rom[1853] = 25'b0000000000000000011010001;
    rom[1854] = 25'b0000000000000000011010001;
    rom[1855] = 25'b0000000000000000011010010;
    rom[1856] = 25'b0000000000000000011010010;
    rom[1857] = 25'b0000000000000000011010011;
    rom[1858] = 25'b0000000000000000011010011;
    rom[1859] = 25'b0000000000000000011010100;
    rom[1860] = 25'b0000000000000000011010101;
    rom[1861] = 25'b0000000000000000011010101;
    rom[1862] = 25'b0000000000000000011010110;
    rom[1863] = 25'b0000000000000000011010111;
    rom[1864] = 25'b0000000000000000011011000;
    rom[1865] = 25'b0000000000000000011011000;
    rom[1866] = 25'b0000000000000000011011000;
    rom[1867] = 25'b0000000000000000011011001;
    rom[1868] = 25'b0000000000000000011011001;
    rom[1869] = 25'b0000000000000000011011010;
    rom[1870] = 25'b0000000000000000011011011;
    rom[1871] = 25'b0000000000000000011011011;
    rom[1872] = 25'b0000000000000000011011100;
    rom[1873] = 25'b0000000000000000011011101;
    rom[1874] = 25'b0000000000000000011011101;
    rom[1875] = 25'b0000000000000000011011101;
    rom[1876] = 25'b0000000000000000011011110;
    rom[1877] = 25'b0000000000000000011011110;
    rom[1878] = 25'b0000000000000000011011111;
    rom[1879] = 25'b0000000000000000011011111;
    rom[1880] = 25'b0000000000000000011100000;
    rom[1881] = 25'b0000000000000000011100001;
    rom[1882] = 25'b0000000000000000011100001;
    rom[1883] = 25'b0000000000000000011100010;
    rom[1884] = 25'b0000000000000000011100010;
    rom[1885] = 25'b0000000000000000011100011;
    rom[1886] = 25'b0000000000000000011100011;
    rom[1887] = 25'b0000000000000000011100011;
    rom[1888] = 25'b0000000000000000011100100;
    rom[1889] = 25'b0000000000000000011100100;
    rom[1890] = 25'b0000000000000000011100101;
    rom[1891] = 25'b0000000000000000011100101;
    rom[1892] = 25'b0000000000000000011100110;
    rom[1893] = 25'b0000000000000000011100110;
    rom[1894] = 25'b0000000000000000011100111;
    rom[1895] = 25'b0000000000000000011101000;
    rom[1896] = 25'b0000000000000000011101000;
    rom[1897] = 25'b0000000000000000011101001;
    rom[1898] = 25'b0000000000000000011101001;
    rom[1899] = 25'b0000000000000000011101001;
    rom[1900] = 25'b0000000000000000011101001;
    rom[1901] = 25'b0000000000000000011101001;
    rom[1902] = 25'b0000000000000000011101010;
    rom[1903] = 25'b0000000000000000011101010;
    rom[1904] = 25'b0000000000000000011101011;
    rom[1905] = 25'b0000000000000000011101011;
    rom[1906] = 25'b0000000000000000011101100;
    rom[1907] = 25'b0000000000000000011101100;
    rom[1908] = 25'b0000000000000000011101101;
    rom[1909] = 25'b0000000000000000011101101;
    rom[1910] = 25'b0000000000000000011101101;
    rom[1911] = 25'b0000000000000000011101110;
    rom[1912] = 25'b0000000000000000011101110;
    rom[1913] = 25'b0000000000000000011101110;
    rom[1914] = 25'b0000000000000000011101110;
    rom[1915] = 25'b0000000000000000011101110;
    rom[1916] = 25'b0000000000000000011101111;
    rom[1917] = 25'b0000000000000000011101111;
    rom[1918] = 25'b0000000000000000011110000;
    rom[1919] = 25'b0000000000000000011110000;
    rom[1920] = 25'b0000000000000000011110000;
    rom[1921] = 25'b0000000000000000011110001;
    rom[1922] = 25'b0000000000000000011110001;
    rom[1923] = 25'b0000000000000000011110001;
    rom[1924] = 25'b0000000000000000011110001;
    rom[1925] = 25'b0000000000000000011110010;
    rom[1926] = 25'b0000000000000000011110010;
    rom[1927] = 25'b0000000000000000011110010;
    rom[1928] = 25'b0000000000000000011110011;
    rom[1929] = 25'b0000000000000000011110011;
    rom[1930] = 25'b0000000000000000011110011;
    rom[1931] = 25'b0000000000000000011110011;
    rom[1932] = 25'b0000000000000000011110100;
    rom[1933] = 25'b0000000000000000011110100;
    rom[1934] = 25'b0000000000000000011110100;
    rom[1935] = 25'b0000000000000000011110100;
    rom[1936] = 25'b0000000000000000011110100;
    rom[1937] = 25'b0000000000000000011110100;
    rom[1938] = 25'b0000000000000000011110100;
    rom[1939] = 25'b0000000000000000011110100;
    rom[1940] = 25'b0000000000000000011110100;
    rom[1941] = 25'b0000000000000000011110100;
    rom[1942] = 25'b0000000000000000011110101;
    rom[1943] = 25'b0000000000000000011110101;
    rom[1944] = 25'b0000000000000000011110101;
    rom[1945] = 25'b0000000000000000011110101;
    rom[1946] = 25'b0000000000000000011110101;
    rom[1947] = 25'b0000000000000000011110101;
    rom[1948] = 25'b0000000000000000011110101;
    rom[1949] = 25'b0000000000000000011110101;
    rom[1950] = 25'b0000000000000000011110101;
    rom[1951] = 25'b0000000000000000011110101;
    rom[1952] = 25'b0000000000000000011110110;
    rom[1953] = 25'b0000000000000000011110110;
    rom[1954] = 25'b0000000000000000011110110;
    rom[1955] = 25'b0000000000000000011110110;
    rom[1956] = 25'b0000000000000000011110110;
    rom[1957] = 25'b0000000000000000011110110;
    rom[1958] = 25'b0000000000000000011110110;
    rom[1959] = 25'b0000000000000000011110110;
    rom[1960] = 25'b0000000000000000011110110;
    rom[1961] = 25'b0000000000000000011110110;
    rom[1962] = 25'b0000000000000000011110110;
    rom[1963] = 25'b0000000000000000011110110;
    rom[1964] = 25'b0000000000000000011110101;
    rom[1965] = 25'b0000000000000000011110101;
    rom[1966] = 25'b0000000000000000011110101;
    rom[1967] = 25'b0000000000000000011110101;
    rom[1968] = 25'b0000000000000000011110101;
    rom[1969] = 25'b0000000000000000011110101;
    rom[1970] = 25'b0000000000000000011110101;
    rom[1971] = 25'b0000000000000000011110101;
    rom[1972] = 25'b0000000000000000011110101;
    rom[1973] = 25'b0000000000000000011110100;
    rom[1974] = 25'b0000000000000000011110100;
    rom[1975] = 25'b0000000000000000011110100;
    rom[1976] = 25'b0000000000000000011110100;
    rom[1977] = 25'b0000000000000000011110100;
    rom[1978] = 25'b0000000000000000011110100;
    rom[1979] = 25'b0000000000000000011110100;
    rom[1980] = 25'b0000000000000000011110100;
    rom[1981] = 25'b0000000000000000011110100;
    rom[1982] = 25'b0000000000000000011110100;
    rom[1983] = 25'b0000000000000000011110011;
    rom[1984] = 25'b0000000000000000011110011;
    rom[1985] = 25'b0000000000000000011110011;
    rom[1986] = 25'b0000000000000000011110010;
    rom[1987] = 25'b0000000000000000011110010;
    rom[1988] = 25'b0000000000000000011110010;
    rom[1989] = 25'b0000000000000000011110010;
    rom[1990] = 25'b0000000000000000011110001;
    rom[1991] = 25'b0000000000000000011110001;
    rom[1992] = 25'b0000000000000000011110000;
    rom[1993] = 25'b0000000000000000011110000;
    rom[1994] = 25'b0000000000000000011110000;
    rom[1995] = 25'b0000000000000000011101111;
    rom[1996] = 25'b0000000000000000011101111;
    rom[1997] = 25'b0000000000000000011101110;
    rom[1998] = 25'b0000000000000000011101110;
    rom[1999] = 25'b0000000000000000011101110;
    rom[2000] = 25'b0000000000000000011101110;
    rom[2001] = 25'b0000000000000000011101110;
    rom[2002] = 25'b0000000000000000011101101;
    rom[2003] = 25'b0000000000000000011101101;
    rom[2004] = 25'b0000000000000000011101100;
    rom[2005] = 25'b0000000000000000011101100;
    rom[2006] = 25'b0000000000000000011101011;
    rom[2007] = 25'b0000000000000000011101011;
    rom[2008] = 25'b0000000000000000011101010;
    rom[2009] = 25'b0000000000000000011101010;
    rom[2010] = 25'b0000000000000000011101001;
    rom[2011] = 25'b0000000000000000011101001;
    rom[2012] = 25'b0000000000000000011101001;
    rom[2013] = 25'b0000000000000000011101000;
    rom[2014] = 25'b0000000000000000011101000;
    rom[2015] = 25'b0000000000000000011100111;
    rom[2016] = 25'b0000000000000000011100110;
    rom[2017] = 25'b0000000000000000011100110;
    rom[2018] = 25'b0000000000000000011100101;
    rom[2019] = 25'b0000000000000000011100100;
    rom[2020] = 25'b0000000000000000011100011;
    rom[2021] = 25'b0000000000000000011100011;
    rom[2022] = 25'b0000000000000000011100011;
    rom[2023] = 25'b0000000000000000011100010;
    rom[2024] = 25'b0000000000000000011100010;
    rom[2025] = 25'b0000000000000000011100001;
    rom[2026] = 25'b0000000000000000011100000;
    rom[2027] = 25'b0000000000000000011011111;
    rom[2028] = 25'b0000000000000000011011110;
    rom[2029] = 25'b0000000000000000011011110;
    rom[2030] = 25'b0000000000000000011011101;
    rom[2031] = 25'b0000000000000000011011101;
    rom[2032] = 25'b0000000000000000011011100;
    rom[2033] = 25'b0000000000000000011011011;
    rom[2034] = 25'b0000000000000000011011010;
    rom[2035] = 25'b0000000000000000011011001;
    rom[2036] = 25'b0000000000000000011011001;
    rom[2037] = 25'b0000000000000000011011000;
    rom[2038] = 25'b0000000000000000011011000;
    rom[2039] = 25'b0000000000000000011010111;
    rom[2040] = 25'b0000000000000000011010110;
    rom[2041] = 25'b0000000000000000011010101;
    rom[2042] = 25'b0000000000000000011010100;
    rom[2043] = 25'b0000000000000000011010011;
    rom[2044] = 25'b0000000000000000011010010;
    rom[2045] = 25'b0000000000000000011010010;
    rom[2046] = 25'b0000000000000000011010001;
    rom[2047] = 25'b0000000000000000011010000;
    rom[2048] = 25'b0000000000000000011001111;
    rom[2049] = 25'b0000000000000000011001101;
    rom[2050] = 25'b0000000000000000011001100;
    rom[2051] = 25'b0000000000000000011001100;
    rom[2052] = 25'b0000000000000000011001011;
    rom[2053] = 25'b0000000000000000011001010;
    rom[2054] = 25'b0000000000000000011001001;
    rom[2055] = 25'b0000000000000000011001000;
    rom[2056] = 25'b0000000000000000011000111;
    rom[2057] = 25'b0000000000000000011000110;
    rom[2058] = 25'b0000000000000000011000101;
    rom[2059] = 25'b0000000000000000011000100;
    rom[2060] = 25'b0000000000000000011000011;
    rom[2061] = 25'b0000000000000000011000001;
    rom[2062] = 25'b0000000000000000011000001;
    rom[2063] = 25'b0000000000000000011000000;
    rom[2064] = 25'b0000000000000000010111111;
    rom[2065] = 25'b0000000000000000010111101;
    rom[2066] = 25'b0000000000000000010111100;
    rom[2067] = 25'b0000000000000000010111011;
    rom[2068] = 25'b0000000000000000010111010;
    rom[2069] = 25'b0000000000000000010111001;
    rom[2070] = 25'b0000000000000000010111000;
    rom[2071] = 25'b0000000000000000010110110;
    rom[2072] = 25'b0000000000000000010110110;
    rom[2073] = 25'b0000000000000000010110100;
    rom[2074] = 25'b0000000000000000010110011;
    rom[2075] = 25'b0000000000000000010110001;
    rom[2076] = 25'b0000000000000000010110000;
    rom[2077] = 25'b0000000000000000010110000;
    rom[2078] = 25'b0000000000000000010101110;
    rom[2079] = 25'b0000000000000000010101101;
    rom[2080] = 25'b0000000000000000010101011;
    rom[2081] = 25'b0000000000000000010101010;
    rom[2082] = 25'b0000000000000000010101001;
    rom[2083] = 25'b0000000000000000010100111;
    rom[2084] = 25'b0000000000000000010100110;
    rom[2085] = 25'b0000000000000000010100100;
    rom[2086] = 25'b0000000000000000010100100;
    rom[2087] = 25'b0000000000000000010100010;
    rom[2088] = 25'b0000000000000000010100000;
    rom[2089] = 25'b0000000000000000010011111;
    rom[2090] = 25'b0000000000000000010011110;
    rom[2091] = 25'b0000000000000000010011100;
    rom[2092] = 25'b0000000000000000010011011;
    rom[2093] = 25'b0000000000000000010011001;
    rom[2094] = 25'b0000000000000000010011000;
    rom[2095] = 25'b0000000000000000010010111;
    rom[2096] = 25'b0000000000000000010010101;
    rom[2097] = 25'b0000000000000000010010011;
    rom[2098] = 25'b0000000000000000010010010;
    rom[2099] = 25'b0000000000000000010010000;
    rom[2100] = 25'b0000000000000000010001111;
    rom[2101] = 25'b0000000000000000010001110;
    rom[2102] = 25'b0000000000000000010001100;
    rom[2103] = 25'b0000000000000000010001010;
    rom[2104] = 25'b0000000000000000010001000;
    rom[2105] = 25'b0000000000000000010000111;
    rom[2106] = 25'b0000000000000000010000101;
    rom[2107] = 25'b0000000000000000010000100;
    rom[2108] = 25'b0000000000000000010000010;
    rom[2109] = 25'b0000000000000000010000001;
    rom[2110] = 25'b0000000000000000001111111;
    rom[2111] = 25'b0000000000000000001111101;
    rom[2112] = 25'b0000000000000000001111100;
    rom[2113] = 25'b0000000000000000001111010;
    rom[2114] = 25'b0000000000000000001111000;
    rom[2115] = 25'b0000000000000000001110111;
    rom[2116] = 25'b0000000000000000001110101;
    rom[2117] = 25'b0000000000000000001110011;
    rom[2118] = 25'b0000000000000000001110001;
    rom[2119] = 25'b0000000000000000001101111;
    rom[2120] = 25'b0000000000000000001101101;
    rom[2121] = 25'b0000000000000000001101100;
    rom[2122] = 25'b0000000000000000001101010;
    rom[2123] = 25'b0000000000000000001101000;
    rom[2124] = 25'b0000000000000000001100110;
    rom[2125] = 25'b0000000000000000001100101;
    rom[2126] = 25'b0000000000000000001100010;
    rom[2127] = 25'b0000000000000000001100000;
    rom[2128] = 25'b0000000000000000001011111;
    rom[2129] = 25'b0000000000000000001011101;
    rom[2130] = 25'b0000000000000000001011011;
    rom[2131] = 25'b0000000000000000001011001;
    rom[2132] = 25'b0000000000000000001010111;
    rom[2133] = 25'b0000000000000000001010101;
    rom[2134] = 25'b0000000000000000001010011;
    rom[2135] = 25'b0000000000000000001010001;
    rom[2136] = 25'b0000000000000000001001111;
    rom[2137] = 25'b0000000000000000001001101;
    rom[2138] = 25'b0000000000000000001001011;
    rom[2139] = 25'b0000000000000000001001001;
    rom[2140] = 25'b0000000000000000001000111;
    rom[2141] = 25'b0000000000000000001000101;
    rom[2142] = 25'b0000000000000000001000011;
    rom[2143] = 25'b0000000000000000001000001;
    rom[2144] = 25'b0000000000000000000111110;
    rom[2145] = 25'b0000000000000000000111101;
    rom[2146] = 25'b0000000000000000000111010;
    rom[2147] = 25'b0000000000000000000111000;
    rom[2148] = 25'b0000000000000000000110110;
    rom[2149] = 25'b0000000000000000000110100;
    rom[2150] = 25'b0000000000000000000110010;
    rom[2151] = 25'b0000000000000000000110000;
    rom[2152] = 25'b0000000000000000000101101;
    rom[2153] = 25'b0000000000000000000101100;
    rom[2154] = 25'b0000000000000000000101001;
    rom[2155] = 25'b0000000000000000000100111;
    rom[2156] = 25'b0000000000000000000100101;
    rom[2157] = 25'b0000000000000000000100010;
    rom[2158] = 25'b0000000000000000000100000;
    rom[2159] = 25'b0000000000000000000011110;
    rom[2160] = 25'b0000000000000000000011100;
    rom[2161] = 25'b0000000000000000000011001;
    rom[2162] = 25'b0000000000000000000010111;
    rom[2163] = 25'b0000000000000000000010101;
    rom[2164] = 25'b0000000000000000000010010;
    rom[2165] = 25'b0000000000000000000010000;
    rom[2166] = 25'b0000000000000000000001110;
    rom[2167] = 25'b0000000000000000000001011;
    rom[2168] = 25'b0000000000000000000001001;
    rom[2169] = 25'b0000000000000000000000110;
    rom[2170] = 25'b0000000000000000000000100;
    rom[2171] = 25'b0000000000000000000000001;
    rom[2172] = 25'b0000000000000000000000000;
    rom[2173] = 25'b1111111111111111111111110;
    rom[2174] = 25'b1111111111111111111111011;
    rom[2175] = 25'b1111111111111111111111001;
    rom[2176] = 25'b1111111111111111111110110;
    rom[2177] = 25'b1111111111111111111110100;
    rom[2178] = 25'b1111111111111111111110001;
    rom[2179] = 25'b1111111111111111111101110;
    rom[2180] = 25'b1111111111111111111101100;
    rom[2181] = 25'b1111111111111111111101001;
    rom[2182] = 25'b1111111111111111111100111;
    rom[2183] = 25'b1111111111111111111100100;
    rom[2184] = 25'b1111111111111111111100010;
    rom[2185] = 25'b1111111111111111111011111;
    rom[2186] = 25'b1111111111111111111011101;
    rom[2187] = 25'b1111111111111111111011010;
    rom[2188] = 25'b1111111111111111111011000;
    rom[2189] = 25'b1111111111111111111010101;
    rom[2190] = 25'b1111111111111111111010010;
    rom[2191] = 25'b1111111111111111111010000;
    rom[2192] = 25'b1111111111111111111001100;
    rom[2193] = 25'b1111111111111111111001010;
    rom[2194] = 25'b1111111111111111111000111;
    rom[2195] = 25'b1111111111111111111000101;
    rom[2196] = 25'b1111111111111111111000010;
    rom[2197] = 25'b1111111111111111111000000;
    rom[2198] = 25'b1111111111111111110111100;
    rom[2199] = 25'b1111111111111111110111010;
    rom[2200] = 25'b1111111111111111110110111;
    rom[2201] = 25'b1111111111111111110110101;
    rom[2202] = 25'b1111111111111111110110001;
    rom[2203] = 25'b1111111111111111110101111;
    rom[2204] = 25'b1111111111111111110101100;
    rom[2205] = 25'b1111111111111111110101001;
    rom[2206] = 25'b1111111111111111110100110;
    rom[2207] = 25'b1111111111111111110100100;
    rom[2208] = 25'b1111111111111111110100000;
    rom[2209] = 25'b1111111111111111110011110;
    rom[2210] = 25'b1111111111111111110011011;
    rom[2211] = 25'b1111111111111111110011000;
    rom[2212] = 25'b1111111111111111110010101;
    rom[2213] = 25'b1111111111111111110010011;
    rom[2214] = 25'b1111111111111111110001111;
    rom[2215] = 25'b1111111111111111110001101;
    rom[2216] = 25'b1111111111111111110001001;
    rom[2217] = 25'b1111111111111111110000111;
    rom[2218] = 25'b1111111111111111110000011;
    rom[2219] = 25'b1111111111111111110000001;
    rom[2220] = 25'b1111111111111111101111101;
    rom[2221] = 25'b1111111111111111101111011;
    rom[2222] = 25'b1111111111111111101110111;
    rom[2223] = 25'b1111111111111111101110101;
    rom[2224] = 25'b1111111111111111101110001;
    rom[2225] = 25'b1111111111111111101101111;
    rom[2226] = 25'b1111111111111111101101100;
    rom[2227] = 25'b1111111111111111101101001;
    rom[2228] = 25'b1111111111111111101100110;
    rom[2229] = 25'b1111111111111111101100010;
    rom[2230] = 25'b1111111111111111101100000;
    rom[2231] = 25'b1111111111111111101011100;
    rom[2232] = 25'b1111111111111111101011001;
    rom[2233] = 25'b1111111111111111101010110;
    rom[2234] = 25'b1111111111111111101010011;
    rom[2235] = 25'b1111111111111111101010000;
    rom[2236] = 25'b1111111111111111101001101;
    rom[2237] = 25'b1111111111111111101001001;
    rom[2238] = 25'b1111111111111111101000110;
    rom[2239] = 25'b1111111111111111101000100;
    rom[2240] = 25'b1111111111111111101000000;
    rom[2241] = 25'b1111111111111111100111101;
    rom[2242] = 25'b1111111111111111100111010;
    rom[2243] = 25'b1111111111111111100110111;
    rom[2244] = 25'b1111111111111111100110011;
    rom[2245] = 25'b1111111111111111100110000;
    rom[2246] = 25'b1111111111111111100101101;
    rom[2247] = 25'b1111111111111111100101010;
    rom[2248] = 25'b1111111111111111100100111;
    rom[2249] = 25'b1111111111111111100100011;
    rom[2250] = 25'b1111111111111111100100000;
    rom[2251] = 25'b1111111111111111100011100;
    rom[2252] = 25'b1111111111111111100011010;
    rom[2253] = 25'b1111111111111111100010110;
    rom[2254] = 25'b1111111111111111100010011;
    rom[2255] = 25'b1111111111111111100010000;
    rom[2256] = 25'b1111111111111111100001100;
    rom[2257] = 25'b1111111111111111100001001;
    rom[2258] = 25'b1111111111111111100000101;
    rom[2259] = 25'b1111111111111111100000010;
    rom[2260] = 25'b1111111111111111100000000;
    rom[2261] = 25'b1111111111111111011111100;
    rom[2262] = 25'b1111111111111111011111001;
    rom[2263] = 25'b1111111111111111011110101;
    rom[2264] = 25'b1111111111111111011110010;
    rom[2265] = 25'b1111111111111111011101110;
    rom[2266] = 25'b1111111111111111011101011;
    rom[2267] = 25'b1111111111111111011101000;
    rom[2268] = 25'b1111111111111111011100100;
    rom[2269] = 25'b1111111111111111011100001;
    rom[2270] = 25'b1111111111111111011011101;
    rom[2271] = 25'b1111111111111111011011010;
    rom[2272] = 25'b1111111111111111011010111;
    rom[2273] = 25'b1111111111111111011010011;
    rom[2274] = 25'b1111111111111111011010000;
    rom[2275] = 25'b1111111111111111011001100;
    rom[2276] = 25'b1111111111111111011001001;
    rom[2277] = 25'b1111111111111111011000110;
    rom[2278] = 25'b1111111111111111011000010;
    rom[2279] = 25'b1111111111111111010111111;
    rom[2280] = 25'b1111111111111111010111011;
    rom[2281] = 25'b1111111111111111010110111;
    rom[2282] = 25'b1111111111111111010110100;
    rom[2283] = 25'b1111111111111111010110000;
    rom[2284] = 25'b1111111111111111010101101;
    rom[2285] = 25'b1111111111111111010101010;
    rom[2286] = 25'b1111111111111111010100110;
    rom[2287] = 25'b1111111111111111010100011;
    rom[2288] = 25'b1111111111111111010011111;
    rom[2289] = 25'b1111111111111111010011100;
    rom[2290] = 25'b1111111111111111010011000;
    rom[2291] = 25'b1111111111111111010010100;
    rom[2292] = 25'b1111111111111111010010001;
    rom[2293] = 25'b1111111111111111010001110;
    rom[2294] = 25'b1111111111111111010001010;
    rom[2295] = 25'b1111111111111111010000111;
    rom[2296] = 25'b1111111111111111010000010;
    rom[2297] = 25'b1111111111111111001111111;
    rom[2298] = 25'b1111111111111111001111100;
    rom[2299] = 25'b1111111111111111001111000;
    rom[2300] = 25'b1111111111111111001110101;
    rom[2301] = 25'b1111111111111111001110001;
    rom[2302] = 25'b1111111111111111001101101;
    rom[2303] = 25'b1111111111111111001101010;
    rom[2304] = 25'b1111111111111111001100110;
    rom[2305] = 25'b1111111111111111001100011;
    rom[2306] = 25'b1111111111111111001011111;
    rom[2307] = 25'b1111111111111111001011011;
    rom[2308] = 25'b1111111111111111001011000;
    rom[2309] = 25'b1111111111111111001010101;
    rom[2310] = 25'b1111111111111111001010001;
    rom[2311] = 25'b1111111111111111001001101;
    rom[2312] = 25'b1111111111111111001001001;
    rom[2313] = 25'b1111111111111111001000110;
    rom[2314] = 25'b1111111111111111001000011;
    rom[2315] = 25'b1111111111111111000111110;
    rom[2316] = 25'b1111111111111111000111011;
    rom[2317] = 25'b1111111111111111000111000;
    rom[2318] = 25'b1111111111111111000110100;
    rom[2319] = 25'b1111111111111111000110000;
    rom[2320] = 25'b1111111111111111000101101;
    rom[2321] = 25'b1111111111111111000101001;
    rom[2322] = 25'b1111111111111111000100110;
    rom[2323] = 25'b1111111111111111000100010;
    rom[2324] = 25'b1111111111111111000011110;
    rom[2325] = 25'b1111111111111111000011011;
    rom[2326] = 25'b1111111111111111000010110;
    rom[2327] = 25'b1111111111111111000010011;
    rom[2328] = 25'b1111111111111111000010000;
    rom[2329] = 25'b1111111111111111000001100;
    rom[2330] = 25'b1111111111111111000001000;
    rom[2331] = 25'b1111111111111111000000101;
    rom[2332] = 25'b1111111111111111000000001;
    rom[2333] = 25'b1111111111111110111111110;
    rom[2334] = 25'b1111111111111110111111010;
    rom[2335] = 25'b1111111111111110111110110;
    rom[2336] = 25'b1111111111111110111110011;
    rom[2337] = 25'b1111111111111110111101110;
    rom[2338] = 25'b1111111111111110111101011;
    rom[2339] = 25'b1111111111111110111101000;
    rom[2340] = 25'b1111111111111110111100100;
    rom[2341] = 25'b1111111111111110111100000;
    rom[2342] = 25'b1111111111111110111011101;
    rom[2343] = 25'b1111111111111110111011001;
    rom[2344] = 25'b1111111111111110111010110;
    rom[2345] = 25'b1111111111111110111010010;
    rom[2346] = 25'b1111111111111110111001110;
    rom[2347] = 25'b1111111111111110111001011;
    rom[2348] = 25'b1111111111111110111000111;
    rom[2349] = 25'b1111111111111110111000011;
    rom[2350] = 25'b1111111111111110111000000;
    rom[2351] = 25'b1111111111111110110111100;
    rom[2352] = 25'b1111111111111110110111000;
    rom[2353] = 25'b1111111111111110110110101;
    rom[2354] = 25'b1111111111111110110110001;
    rom[2355] = 25'b1111111111111110110101110;
    rom[2356] = 25'b1111111111111110110101010;
    rom[2357] = 25'b1111111111111110110100110;
    rom[2358] = 25'b1111111111111110110100011;
    rom[2359] = 25'b1111111111111110110011111;
    rom[2360] = 25'b1111111111111110110011011;
    rom[2361] = 25'b1111111111111110110011000;
    rom[2362] = 25'b1111111111111110110010100;
    rom[2363] = 25'b1111111111111110110010001;
    rom[2364] = 25'b1111111111111110110001110;
    rom[2365] = 25'b1111111111111110110001001;
    rom[2366] = 25'b1111111111111110110000110;
    rom[2367] = 25'b1111111111111110110000010;
    rom[2368] = 25'b1111111111111110101111111;
    rom[2369] = 25'b1111111111111110101111011;
    rom[2370] = 25'b1111111111111110101110111;
    rom[2371] = 25'b1111111111111110101110100;
    rom[2372] = 25'b1111111111111110101110001;
    rom[2373] = 25'b1111111111111110101101101;
    rom[2374] = 25'b1111111111111110101101010;
    rom[2375] = 25'b1111111111111110101100110;
    rom[2376] = 25'b1111111111111110101100010;
    rom[2377] = 25'b1111111111111110101011111;
    rom[2378] = 25'b1111111111111110101011011;
    rom[2379] = 25'b1111111111111110101011000;
    rom[2380] = 25'b1111111111111110101010101;
    rom[2381] = 25'b1111111111111110101010001;
    rom[2382] = 25'b1111111111111110101001101;
    rom[2383] = 25'b1111111111111110101001001;
    rom[2384] = 25'b1111111111111110101000110;
    rom[2385] = 25'b1111111111111110101000011;
    rom[2386] = 25'b1111111111111110100111111;
    rom[2387] = 25'b1111111111111110100111100;
    rom[2388] = 25'b1111111111111110100111000;
    rom[2389] = 25'b1111111111111110100110101;
    rom[2390] = 25'b1111111111111110100110010;
    rom[2391] = 25'b1111111111111110100101110;
    rom[2392] = 25'b1111111111111110100101011;
    rom[2393] = 25'b1111111111111110100100111;
    rom[2394] = 25'b1111111111111110100100100;
    rom[2395] = 25'b1111111111111110100100001;
    rom[2396] = 25'b1111111111111110100011101;
    rom[2397] = 25'b1111111111111110100011010;
    rom[2398] = 25'b1111111111111110100010110;
    rom[2399] = 25'b1111111111111110100010011;
    rom[2400] = 25'b1111111111111110100010000;
    rom[2401] = 25'b1111111111111110100001100;
    rom[2402] = 25'b1111111111111110100001001;
    rom[2403] = 25'b1111111111111110100000101;
    rom[2404] = 25'b1111111111111110100000010;
    rom[2405] = 25'b1111111111111110011111111;
    rom[2406] = 25'b1111111111111110011111011;
    rom[2407] = 25'b1111111111111110011111001;
    rom[2408] = 25'b1111111111111110011110101;
    rom[2409] = 25'b1111111111111110011110010;
    rom[2410] = 25'b1111111111111110011101110;
    rom[2411] = 25'b1111111111111110011101011;
    rom[2412] = 25'b1111111111111110011101000;
    rom[2413] = 25'b1111111111111110011100101;
    rom[2414] = 25'b1111111111111110011100010;
    rom[2415] = 25'b1111111111111110011011110;
    rom[2416] = 25'b1111111111111110011011011;
    rom[2417] = 25'b1111111111111110011011000;
    rom[2418] = 25'b1111111111111110011010101;
    rom[2419] = 25'b1111111111111110011010010;
    rom[2420] = 25'b1111111111111110011001110;
    rom[2421] = 25'b1111111111111110011001100;
    rom[2422] = 25'b1111111111111110011001000;
    rom[2423] = 25'b1111111111111110011000101;
    rom[2424] = 25'b1111111111111110011000010;
    rom[2425] = 25'b1111111111111110010111111;
    rom[2426] = 25'b1111111111111110010111011;
    rom[2427] = 25'b1111111111111110010111001;
    rom[2428] = 25'b1111111111111110010110110;
    rom[2429] = 25'b1111111111111110010110011;
    rom[2430] = 25'b1111111111111110010110000;
    rom[2431] = 25'b1111111111111110010101101;
    rom[2432] = 25'b1111111111111110010101010;
    rom[2433] = 25'b1111111111111110010100111;
    rom[2434] = 25'b1111111111111110010100100;
    rom[2435] = 25'b1111111111111110010100001;
    rom[2436] = 25'b1111111111111110010011110;
    rom[2437] = 25'b1111111111111110010011011;
    rom[2438] = 25'b1111111111111110010011000;
    rom[2439] = 25'b1111111111111110010010101;
    rom[2440] = 25'b1111111111111110010010011;
    rom[2441] = 25'b1111111111111110010001111;
    rom[2442] = 25'b1111111111111110010001101;
    rom[2443] = 25'b1111111111111110010001010;
    rom[2444] = 25'b1111111111111110010000111;
    rom[2445] = 25'b1111111111111110010000100;
    rom[2446] = 25'b1111111111111110010000010;
    rom[2447] = 25'b1111111111111110001111110;
    rom[2448] = 25'b1111111111111110001111100;
    rom[2449] = 25'b1111111111111110001111001;
    rom[2450] = 25'b1111111111111110001110111;
    rom[2451] = 25'b1111111111111110001110100;
    rom[2452] = 25'b1111111111111110001110001;
    rom[2453] = 25'b1111111111111110001101110;
    rom[2454] = 25'b1111111111111110001101100;
    rom[2455] = 25'b1111111111111110001101001;
    rom[2456] = 25'b1111111111111110001100110;
    rom[2457] = 25'b1111111111111110001100100;
    rom[2458] = 25'b1111111111111110001100001;
    rom[2459] = 25'b1111111111111110001011111;
    rom[2460] = 25'b1111111111111110001011100;
    rom[2461] = 25'b1111111111111110001011010;
    rom[2462] = 25'b1111111111111110001010111;
    rom[2463] = 25'b1111111111111110001010101;
    rom[2464] = 25'b1111111111111110001010010;
    rom[2465] = 25'b1111111111111110001010000;
    rom[2466] = 25'b1111111111111110001001110;
    rom[2467] = 25'b1111111111111110001001011;
    rom[2468] = 25'b1111111111111110001001001;
    rom[2469] = 25'b1111111111111110001000110;
    rom[2470] = 25'b1111111111111110001000100;
    rom[2471] = 25'b1111111111111110001000010;
    rom[2472] = 25'b1111111111111110000111111;
    rom[2473] = 25'b1111111111111110000111110;
    rom[2474] = 25'b1111111111111110000111011;
    rom[2475] = 25'b1111111111111110000111000;
    rom[2476] = 25'b1111111111111110000110111;
    rom[2477] = 25'b1111111111111110000110100;
    rom[2478] = 25'b1111111111111110000110011;
    rom[2479] = 25'b1111111111111110000110000;
    rom[2480] = 25'b1111111111111110000101110;
    rom[2481] = 25'b1111111111111110000101100;
    rom[2482] = 25'b1111111111111110000101010;
    rom[2483] = 25'b1111111111111110000100111;
    rom[2484] = 25'b1111111111111110000100110;
    rom[2485] = 25'b1111111111111110000100100;
    rom[2486] = 25'b1111111111111110000100010;
    rom[2487] = 25'b1111111111111110000100000;
    rom[2488] = 25'b1111111111111110000011110;
    rom[2489] = 25'b1111111111111110000011100;
    rom[2490] = 25'b1111111111111110000011010;
    rom[2491] = 25'b1111111111111110000011000;
    rom[2492] = 25'b1111111111111110000010110;
    rom[2493] = 25'b1111111111111110000010101;
    rom[2494] = 25'b1111111111111110000010011;
    rom[2495] = 25'b1111111111111110000010001;
    rom[2496] = 25'b1111111111111110000001111;
    rom[2497] = 25'b1111111111111110000001101;
    rom[2498] = 25'b1111111111111110000001011;
    rom[2499] = 25'b1111111111111110000001011;
    rom[2500] = 25'b1111111111111110000001001;
    rom[2501] = 25'b1111111111111110000000111;
    rom[2502] = 25'b1111111111111110000000101;
    rom[2503] = 25'b1111111111111110000000100;
    rom[2504] = 25'b1111111111111110000000010;
    rom[2505] = 25'b1111111111111110000000000;
    rom[2506] = 25'b1111111111111110000000000;
    rom[2507] = 25'b1111111111111101111111110;
    rom[2508] = 25'b1111111111111101111111100;
    rom[2509] = 25'b1111111111111101111111011;
    rom[2510] = 25'b1111111111111101111111010;
    rom[2511] = 25'b1111111111111101111111001;
    rom[2512] = 25'b1111111111111101111110111;
    rom[2513] = 25'b1111111111111101111110101;
    rom[2514] = 25'b1111111111111101111110100;
    rom[2515] = 25'b1111111111111101111110100;
    rom[2516] = 25'b1111111111111101111110010;
    rom[2517] = 25'b1111111111111101111110001;
    rom[2518] = 25'b1111111111111101111101111;
    rom[2519] = 25'b1111111111111101111101110;
    rom[2520] = 25'b1111111111111101111101110;
    rom[2521] = 25'b1111111111111101111101101;
    rom[2522] = 25'b1111111111111101111101011;
    rom[2523] = 25'b1111111111111101111101010;
    rom[2524] = 25'b1111111111111101111101001;
    rom[2525] = 25'b1111111111111101111101001;
    rom[2526] = 25'b1111111111111101111101000;
    rom[2527] = 25'b1111111111111101111100111;
    rom[2528] = 25'b1111111111111101111100110;
    rom[2529] = 25'b1111111111111101111100101;
    rom[2530] = 25'b1111111111111101111100100;
    rom[2531] = 25'b1111111111111101111100011;
    rom[2532] = 25'b1111111111111101111100011;
    rom[2533] = 25'b1111111111111101111100011;
    rom[2534] = 25'b1111111111111101111100010;
    rom[2535] = 25'b1111111111111101111100001;
    rom[2536] = 25'b1111111111111101111100000;
    rom[2537] = 25'b1111111111111101111100000;
    rom[2538] = 25'b1111111111111101111011111;
    rom[2539] = 25'b1111111111111101111011111;
    rom[2540] = 25'b1111111111111101111011110;
    rom[2541] = 25'b1111111111111101111011101;
    rom[2542] = 25'b1111111111111101111011101;
    rom[2543] = 25'b1111111111111101111011101;
    rom[2544] = 25'b1111111111111101111011101;
    rom[2545] = 25'b1111111111111101111011101;
    rom[2546] = 25'b1111111111111101111011101;
    rom[2547] = 25'b1111111111111101111011100;
    rom[2548] = 25'b1111111111111101111011100;
    rom[2549] = 25'b1111111111111101111011100;
    rom[2550] = 25'b1111111111111101111011100;
    rom[2551] = 25'b1111111111111101111011100;
    rom[2552] = 25'b1111111111111101111011100;
    rom[2553] = 25'b1111111111111101111011100;
    rom[2554] = 25'b1111111111111101111011100;
    rom[2555] = 25'b1111111111111101111011100;
    rom[2556] = 25'b1111111111111101111011100;
    rom[2557] = 25'b1111111111111101111011100;
    rom[2558] = 25'b1111111111111101111011100;
    rom[2559] = 25'b1111111111111101111011100;
    rom[2560] = 25'b1111111111111101111011101;
    rom[2561] = 25'b1111111111111101111011101;
    rom[2562] = 25'b1111111111111101111011101;
    rom[2563] = 25'b1111111111111101111011101;
    rom[2564] = 25'b1111111111111101111011101;
    rom[2565] = 25'b1111111111111101111011101;
    rom[2566] = 25'b1111111111111101111011110;
    rom[2567] = 25'b1111111111111101111011111;
    rom[2568] = 25'b1111111111111101111011111;
    rom[2569] = 25'b1111111111111101111100000;
    rom[2570] = 25'b1111111111111101111100001;
    rom[2571] = 25'b1111111111111101111100001;
    rom[2572] = 25'b1111111111111101111100010;
    rom[2573] = 25'b1111111111111101111100011;
    rom[2574] = 25'b1111111111111101111100011;
    rom[2575] = 25'b1111111111111101111100100;
    rom[2576] = 25'b1111111111111101111100101;
    rom[2577] = 25'b1111111111111101111100110;
    rom[2578] = 25'b1111111111111101111100111;
    rom[2579] = 25'b1111111111111101111101000;
    rom[2580] = 25'b1111111111111101111101001;
    rom[2581] = 25'b1111111111111101111101001;
    rom[2582] = 25'b1111111111111101111101010;
    rom[2583] = 25'b1111111111111101111101100;
    rom[2584] = 25'b1111111111111101111101101;
    rom[2585] = 25'b1111111111111101111101110;
    rom[2586] = 25'b1111111111111101111101111;
    rom[2587] = 25'b1111111111111101111110000;
    rom[2588] = 25'b1111111111111101111110010;
    rom[2589] = 25'b1111111111111101111110011;
    rom[2590] = 25'b1111111111111101111110100;
    rom[2591] = 25'b1111111111111101111110110;
    rom[2592] = 25'b1111111111111101111110111;
    rom[2593] = 25'b1111111111111101111111001;
    rom[2594] = 25'b1111111111111101111111010;
    rom[2595] = 25'b1111111111111101111111100;
    rom[2596] = 25'b1111111111111101111111110;
    rom[2597] = 25'b1111111111111110000000000;
    rom[2598] = 25'b1111111111111110000000001;
    rom[2599] = 25'b1111111111111110000000011;
    rom[2600] = 25'b1111111111111110000000101;
    rom[2601] = 25'b1111111111111110000000110;
    rom[2602] = 25'b1111111111111110000001000;
    rom[2603] = 25'b1111111111111110000001010;
    rom[2604] = 25'b1111111111111110000001100;
    rom[2605] = 25'b1111111111111110000001110;
    rom[2606] = 25'b1111111111111110000010000;
    rom[2607] = 25'b1111111111111110000010010;
    rom[2608] = 25'b1111111111111110000010100;
    rom[2609] = 25'b1111111111111110000010110;
    rom[2610] = 25'b1111111111111110000011001;
    rom[2611] = 25'b1111111111111110000011011;
    rom[2612] = 25'b1111111111111110000011101;
    rom[2613] = 25'b1111111111111110000100000;
    rom[2614] = 25'b1111111111111110000100010;
    rom[2615] = 25'b1111111111111110000100100;
    rom[2616] = 25'b1111111111111110000100111;
    rom[2617] = 25'b1111111111111110000101001;
    rom[2618] = 25'b1111111111111110000101100;
    rom[2619] = 25'b1111111111111110000101110;
    rom[2620] = 25'b1111111111111110000110001;
    rom[2621] = 25'b1111111111111110000110100;
    rom[2622] = 25'b1111111111111110000110111;
    rom[2623] = 25'b1111111111111110000111001;
    rom[2624] = 25'b1111111111111110000111100;
    rom[2625] = 25'b1111111111111110000111111;
    rom[2626] = 25'b1111111111111110001000010;
    rom[2627] = 25'b1111111111111110001000101;
    rom[2628] = 25'b1111111111111110001001000;
    rom[2629] = 25'b1111111111111110001001011;
    rom[2630] = 25'b1111111111111110001001110;
    rom[2631] = 25'b1111111111111110001010001;
    rom[2632] = 25'b1111111111111110001010101;
    rom[2633] = 25'b1111111111111110001011000;
    rom[2634] = 25'b1111111111111110001011011;
    rom[2635] = 25'b1111111111111110001011110;
    rom[2636] = 25'b1111111111111110001100001;
    rom[2637] = 25'b1111111111111110001100101;
    rom[2638] = 25'b1111111111111110001101000;
    rom[2639] = 25'b1111111111111110001101100;
    rom[2640] = 25'b1111111111111110001110000;
    rom[2641] = 25'b1111111111111110001110011;
    rom[2642] = 25'b1111111111111110001110111;
    rom[2643] = 25'b1111111111111110001111011;
    rom[2644] = 25'b1111111111111110001111110;
    rom[2645] = 25'b1111111111111110010000010;
    rom[2646] = 25'b1111111111111110010000110;
    rom[2647] = 25'b1111111111111110010001001;
    rom[2648] = 25'b1111111111111110010001110;
    rom[2649] = 25'b1111111111111110010010010;
    rom[2650] = 25'b1111111111111110010010101;
    rom[2651] = 25'b1111111111111110010011001;
    rom[2652] = 25'b1111111111111110010011110;
    rom[2653] = 25'b1111111111111110010100010;
    rom[2654] = 25'b1111111111111110010100110;
    rom[2655] = 25'b1111111111111110010101010;
    rom[2656] = 25'b1111111111111110010101111;
    rom[2657] = 25'b1111111111111110010110011;
    rom[2658] = 25'b1111111111111110010110111;
    rom[2659] = 25'b1111111111111110010111011;
    rom[2660] = 25'b1111111111111110011000001;
    rom[2661] = 25'b1111111111111110011000101;
    rom[2662] = 25'b1111111111111110011001001;
    rom[2663] = 25'b1111111111111110011001110;
    rom[2664] = 25'b1111111111111110011010010;
    rom[2665] = 25'b1111111111111110011011000;
    rom[2666] = 25'b1111111111111110011011101;
    rom[2667] = 25'b1111111111111110011100001;
    rom[2668] = 25'b1111111111111110011100110;
    rom[2669] = 25'b1111111111111110011101011;
    rom[2670] = 25'b1111111111111110011110000;
    rom[2671] = 25'b1111111111111110011110101;
    rom[2672] = 25'b1111111111111110011111010;
    rom[2673] = 25'b1111111111111110100000000;
    rom[2674] = 25'b1111111111111110100000101;
    rom[2675] = 25'b1111111111111110100001010;
    rom[2676] = 25'b1111111111111110100001111;
    rom[2677] = 25'b1111111111111110100010100;
    rom[2678] = 25'b1111111111111110100011001;
    rom[2679] = 25'b1111111111111110100011111;
    rom[2680] = 25'b1111111111111110100100100;
    rom[2681] = 25'b1111111111111110100101010;
    rom[2682] = 25'b1111111111111110100101111;
    rom[2683] = 25'b1111111111111110100110101;
    rom[2684] = 25'b1111111111111110100111011;
    rom[2685] = 25'b1111111111111110101000000;
    rom[2686] = 25'b1111111111111110101000110;
    rom[2687] = 25'b1111111111111110101001100;
    rom[2688] = 25'b1111111111111110101010010;
    rom[2689] = 25'b1111111111111110101011000;
    rom[2690] = 25'b1111111111111110101011110;
    rom[2691] = 25'b1111111111111110101100100;
    rom[2692] = 25'b1111111111111110101101010;
    rom[2693] = 25'b1111111111111110101110000;
    rom[2694] = 25'b1111111111111110101110110;
    rom[2695] = 25'b1111111111111110101111100;
    rom[2696] = 25'b1111111111111110110000010;
    rom[2697] = 25'b1111111111111110110001000;
    rom[2698] = 25'b1111111111111110110001111;
    rom[2699] = 25'b1111111111111110110010101;
    rom[2700] = 25'b1111111111111110110011100;
    rom[2701] = 25'b1111111111111110110100010;
    rom[2702] = 25'b1111111111111110110101001;
    rom[2703] = 25'b1111111111111110110110000;
    rom[2704] = 25'b1111111111111110110110110;
    rom[2705] = 25'b1111111111111110110111101;
    rom[2706] = 25'b1111111111111110111000011;
    rom[2707] = 25'b1111111111111110111001010;
    rom[2708] = 25'b1111111111111110111010001;
    rom[2709] = 25'b1111111111111110111011000;
    rom[2710] = 25'b1111111111111110111011111;
    rom[2711] = 25'b1111111111111110111100110;
    rom[2712] = 25'b1111111111111110111101101;
    rom[2713] = 25'b1111111111111110111110100;
    rom[2714] = 25'b1111111111111110111111011;
    rom[2715] = 25'b1111111111111111000000010;
    rom[2716] = 25'b1111111111111111000001010;
    rom[2717] = 25'b1111111111111111000010001;
    rom[2718] = 25'b1111111111111111000011000;
    rom[2719] = 25'b1111111111111111000100000;
    rom[2720] = 25'b1111111111111111000100111;
    rom[2721] = 25'b1111111111111111000101110;
    rom[2722] = 25'b1111111111111111000110110;
    rom[2723] = 25'b1111111111111111000111110;
    rom[2724] = 25'b1111111111111111001000101;
    rom[2725] = 25'b1111111111111111001001101;
    rom[2726] = 25'b1111111111111111001010101;
    rom[2727] = 25'b1111111111111111001011100;
    rom[2728] = 25'b1111111111111111001100100;
    rom[2729] = 25'b1111111111111111001101100;
    rom[2730] = 25'b1111111111111111001110100;
    rom[2731] = 25'b1111111111111111001111100;
    rom[2732] = 25'b1111111111111111010000100;
    rom[2733] = 25'b1111111111111111010001100;
    rom[2734] = 25'b1111111111111111010010100;
    rom[2735] = 25'b1111111111111111010011100;
    rom[2736] = 25'b1111111111111111010100100;
    rom[2737] = 25'b1111111111111111010101101;
    rom[2738] = 25'b1111111111111111010110110;
    rom[2739] = 25'b1111111111111111010111101;
    rom[2740] = 25'b1111111111111111011000110;
    rom[2741] = 25'b1111111111111111011001110;
    rom[2742] = 25'b1111111111111111011010111;
    rom[2743] = 25'b1111111111111111011011111;
    rom[2744] = 25'b1111111111111111011101000;
    rom[2745] = 25'b1111111111111111011110001;
    rom[2746] = 25'b1111111111111111011111010;
    rom[2747] = 25'b1111111111111111100000010;
    rom[2748] = 25'b1111111111111111100001011;
    rom[2749] = 25'b1111111111111111100010100;
    rom[2750] = 25'b1111111111111111100011100;
    rom[2751] = 25'b1111111111111111100100110;
    rom[2752] = 25'b1111111111111111100101110;
    rom[2753] = 25'b1111111111111111100111000;
    rom[2754] = 25'b1111111111111111101000001;
    rom[2755] = 25'b1111111111111111101001001;
    rom[2756] = 25'b1111111111111111101010011;
    rom[2757] = 25'b1111111111111111101011100;
    rom[2758] = 25'b1111111111111111101100110;
    rom[2759] = 25'b1111111111111111101101111;
    rom[2760] = 25'b1111111111111111101111000;
    rom[2761] = 25'b1111111111111111110000010;
    rom[2762] = 25'b1111111111111111110001011;
    rom[2763] = 25'b1111111111111111110010100;
    rom[2764] = 25'b1111111111111111110011110;
    rom[2765] = 25'b1111111111111111110101000;
    rom[2766] = 25'b1111111111111111110110001;
    rom[2767] = 25'b1111111111111111110111011;
    rom[2768] = 25'b1111111111111111111000101;
    rom[2769] = 25'b1111111111111111111001110;
    rom[2770] = 25'b1111111111111111111011000;
    rom[2771] = 25'b1111111111111111111100010;
    rom[2772] = 25'b1111111111111111111101100;
    rom[2773] = 25'b1111111111111111111110110;
    rom[2774] = 25'b0000000000000000000000000;
    rom[2775] = 25'b0000000000000000000001001;
    rom[2776] = 25'b0000000000000000000010011;
    rom[2777] = 25'b0000000000000000000011101;
    rom[2778] = 25'b0000000000000000000100111;
    rom[2779] = 25'b0000000000000000000110010;
    rom[2780] = 25'b0000000000000000000111100;
    rom[2781] = 25'b0000000000000000001000110;
    rom[2782] = 25'b0000000000000000001010000;
    rom[2783] = 25'b0000000000000000001011011;
    rom[2784] = 25'b0000000000000000001100110;
    rom[2785] = 25'b0000000000000000001110000;
    rom[2786] = 25'b0000000000000000001111011;
    rom[2787] = 25'b0000000000000000010000101;
    rom[2788] = 25'b0000000000000000010001111;
    rom[2789] = 25'b0000000000000000010011010;
    rom[2790] = 25'b0000000000000000010100101;
    rom[2791] = 25'b0000000000000000010110000;
    rom[2792] = 25'b0000000000000000010111011;
    rom[2793] = 25'b0000000000000000011000110;
    rom[2794] = 25'b0000000000000000011010000;
    rom[2795] = 25'b0000000000000000011011011;
    rom[2796] = 25'b0000000000000000011100110;
    rom[2797] = 25'b0000000000000000011110001;
    rom[2798] = 25'b0000000000000000011111100;
    rom[2799] = 25'b0000000000000000100000111;
    rom[2800] = 25'b0000000000000000100010010;
    rom[2801] = 25'b0000000000000000100011101;
    rom[2802] = 25'b0000000000000000100101000;
    rom[2803] = 25'b0000000000000000100110100;
    rom[2804] = 25'b0000000000000000100111111;
    rom[2805] = 25'b0000000000000000101001010;
    rom[2806] = 25'b0000000000000000101010101;
    rom[2807] = 25'b0000000000000000101100001;
    rom[2808] = 25'b0000000000000000101101100;
    rom[2809] = 25'b0000000000000000101111000;
    rom[2810] = 25'b0000000000000000110000011;
    rom[2811] = 25'b0000000000000000110001111;
    rom[2812] = 25'b0000000000000000110011011;
    rom[2813] = 25'b0000000000000000110100110;
    rom[2814] = 25'b0000000000000000110110010;
    rom[2815] = 25'b0000000000000000110111110;
    rom[2816] = 25'b0000000000000000111001010;
    rom[2817] = 25'b0000000000000000111010101;
    rom[2818] = 25'b0000000000000000111100001;
    rom[2819] = 25'b0000000000000000111101101;
    rom[2820] = 25'b0000000000000000111111001;
    rom[2821] = 25'b0000000000000001000000101;
    rom[2822] = 25'b0000000000000001000010001;
    rom[2823] = 25'b0000000000000001000011100;
    rom[2824] = 25'b0000000000000001000101001;
    rom[2825] = 25'b0000000000000001000110101;
    rom[2826] = 25'b0000000000000001001000001;
    rom[2827] = 25'b0000000000000001001001101;
    rom[2828] = 25'b0000000000000001001011010;
    rom[2829] = 25'b0000000000000001001100110;
    rom[2830] = 25'b0000000000000001001110001;
    rom[2831] = 25'b0000000000000001001111110;
    rom[2832] = 25'b0000000000000001010001010;
    rom[2833] = 25'b0000000000000001010010111;
    rom[2834] = 25'b0000000000000001010100011;
    rom[2835] = 25'b0000000000000001010110000;
    rom[2836] = 25'b0000000000000001010111100;
    rom[2837] = 25'b0000000000000001011001000;
    rom[2838] = 25'b0000000000000001011010101;
    rom[2839] = 25'b0000000000000001011100010;
    rom[2840] = 25'b0000000000000001011101110;
    rom[2841] = 25'b0000000000000001011111010;
    rom[2842] = 25'b0000000000000001100000111;
    rom[2843] = 25'b0000000000000001100010100;
    rom[2844] = 25'b0000000000000001100100001;
    rom[2845] = 25'b0000000000000001100101101;
    rom[2846] = 25'b0000000000000001100111010;
    rom[2847] = 25'b0000000000000001101000111;
    rom[2848] = 25'b0000000000000001101010100;
    rom[2849] = 25'b0000000000000001101100000;
    rom[2850] = 25'b0000000000000001101101101;
    rom[2851] = 25'b0000000000000001101111011;
    rom[2852] = 25'b0000000000000001110001000;
    rom[2853] = 25'b0000000000000001110010100;
    rom[2854] = 25'b0000000000000001110100001;
    rom[2855] = 25'b0000000000000001110101111;
    rom[2856] = 25'b0000000000000001110111011;
    rom[2857] = 25'b0000000000000001111001000;
    rom[2858] = 25'b0000000000000001111010110;
    rom[2859] = 25'b0000000000000001111100011;
    rom[2860] = 25'b0000000000000001111110000;
    rom[2861] = 25'b0000000000000001111111101;
    rom[2862] = 25'b0000000000000010000001011;
    rom[2863] = 25'b0000000000000010000010111;
    rom[2864] = 25'b0000000000000010000100101;
    rom[2865] = 25'b0000000000000010000110010;
    rom[2866] = 25'b0000000000000010000111111;
    rom[2867] = 25'b0000000000000010001001101;
    rom[2868] = 25'b0000000000000010001011010;
    rom[2869] = 25'b0000000000000010001100111;
    rom[2870] = 25'b0000000000000010001110101;
    rom[2871] = 25'b0000000000000010010000010;
    rom[2872] = 25'b0000000000000010010001111;
    rom[2873] = 25'b0000000000000010010011101;
    rom[2874] = 25'b0000000000000010010101010;
    rom[2875] = 25'b0000000000000010010111000;
    rom[2876] = 25'b0000000000000010011000110;
    rom[2877] = 25'b0000000000000010011010011;
    rom[2878] = 25'b0000000000000010011100001;
    rom[2879] = 25'b0000000000000010011101110;
    rom[2880] = 25'b0000000000000010011111100;
    rom[2881] = 25'b0000000000000010100001010;
    rom[2882] = 25'b0000000000000010100010111;
    rom[2883] = 25'b0000000000000010100100101;
    rom[2884] = 25'b0000000000000010100110011;
    rom[2885] = 25'b0000000000000010101000000;
    rom[2886] = 25'b0000000000000010101001110;
    rom[2887] = 25'b0000000000000010101011011;
    rom[2888] = 25'b0000000000000010101101001;
    rom[2889] = 25'b0000000000000010101110111;
    rom[2890] = 25'b0000000000000010110000101;
    rom[2891] = 25'b0000000000000010110010011;
    rom[2892] = 25'b0000000000000010110100000;
    rom[2893] = 25'b0000000000000010110101110;
    rom[2894] = 25'b0000000000000010110111011;
    rom[2895] = 25'b0000000000000010111001010;
    rom[2896] = 25'b0000000000000010111011000;
    rom[2897] = 25'b0000000000000010111100101;
    rom[2898] = 25'b0000000000000010111110100;
    rom[2899] = 25'b0000000000000011000000001;
    rom[2900] = 25'b0000000000000011000001111;
    rom[2901] = 25'b0000000000000011000011101;
    rom[2902] = 25'b0000000000000011000101011;
    rom[2903] = 25'b0000000000000011000111000;
    rom[2904] = 25'b0000000000000011001000111;
    rom[2905] = 25'b0000000000000011001010101;
    rom[2906] = 25'b0000000000000011001100011;
    rom[2907] = 25'b0000000000000011001110001;
    rom[2908] = 25'b0000000000000011001111110;
    rom[2909] = 25'b0000000000000011010001101;
    rom[2910] = 25'b0000000000000011010011010;
    rom[2911] = 25'b0000000000000011010101001;
    rom[2912] = 25'b0000000000000011010110110;
    rom[2913] = 25'b0000000000000011011000101;
    rom[2914] = 25'b0000000000000011011010010;
    rom[2915] = 25'b0000000000000011011100001;
    rom[2916] = 25'b0000000000000011011101110;
    rom[2917] = 25'b0000000000000011011111101;
    rom[2918] = 25'b0000000000000011100001011;
    rom[2919] = 25'b0000000000000011100011001;
    rom[2920] = 25'b0000000000000011100100111;
    rom[2921] = 25'b0000000000000011100110101;
    rom[2922] = 25'b0000000000000011101000011;
    rom[2923] = 25'b0000000000000011101010001;
    rom[2924] = 25'b0000000000000011101011111;
    rom[2925] = 25'b0000000000000011101101101;
    rom[2926] = 25'b0000000000000011101111011;
    rom[2927] = 25'b0000000000000011110001001;
    rom[2928] = 25'b0000000000000011110010111;
    rom[2929] = 25'b0000000000000011110100101;
    rom[2930] = 25'b0000000000000011110110011;
    rom[2931] = 25'b0000000000000011111000001;
    rom[2932] = 25'b0000000000000011111001111;
    rom[2933] = 25'b0000000000000011111011101;
    rom[2934] = 25'b0000000000000011111101011;
    rom[2935] = 25'b0000000000000011111111010;
    rom[2936] = 25'b0000000000000100000000111;
    rom[2937] = 25'b0000000000000100000010101;
    rom[2938] = 25'b0000000000000100000100011;
    rom[2939] = 25'b0000000000000100000110001;
    rom[2940] = 25'b0000000000000100000111111;
    rom[2941] = 25'b0000000000000100001001101;
    rom[2942] = 25'b0000000000000100001011011;
    rom[2943] = 25'b0000000000000100001101001;
    rom[2944] = 25'b0000000000000100001110111;
    rom[2945] = 25'b0000000000000100010000101;
    rom[2946] = 25'b0000000000000100010010011;
    rom[2947] = 25'b0000000000000100010100001;
    rom[2948] = 25'b0000000000000100010101111;
    rom[2949] = 25'b0000000000000100010111100;
    rom[2950] = 25'b0000000000000100011001011;
    rom[2951] = 25'b0000000000000100011011000;
    rom[2952] = 25'b0000000000000100011100110;
    rom[2953] = 25'b0000000000000100011110100;
    rom[2954] = 25'b0000000000000100100000010;
    rom[2955] = 25'b0000000000000100100010000;
    rom[2956] = 25'b0000000000000100100011101;
    rom[2957] = 25'b0000000000000100100101100;
    rom[2958] = 25'b0000000000000100100111001;
    rom[2959] = 25'b0000000000000100101000111;
    rom[2960] = 25'b0000000000000100101010101;
    rom[2961] = 25'b0000000000000100101100010;
    rom[2962] = 25'b0000000000000100101110000;
    rom[2963] = 25'b0000000000000100101111101;
    rom[2964] = 25'b0000000000000100110001100;
    rom[2965] = 25'b0000000000000100110011001;
    rom[2966] = 25'b0000000000000100110100111;
    rom[2967] = 25'b0000000000000100110110101;
    rom[2968] = 25'b0000000000000100111000010;
    rom[2969] = 25'b0000000000000100111010000;
    rom[2970] = 25'b0000000000000100111011101;
    rom[2971] = 25'b0000000000000100111101010;
    rom[2972] = 25'b0000000000000100111111000;
    rom[2973] = 25'b0000000000000101000000101;
    rom[2974] = 25'b0000000000000101000010011;
    rom[2975] = 25'b0000000000000101000100001;
    rom[2976] = 25'b0000000000000101000101101;
    rom[2977] = 25'b0000000000000101000111011;
    rom[2978] = 25'b0000000000000101001001001;
    rom[2979] = 25'b0000000000000101001010110;
    rom[2980] = 25'b0000000000000101001100011;
    rom[2981] = 25'b0000000000000101001110001;
    rom[2982] = 25'b0000000000000101001111101;
    rom[2983] = 25'b0000000000000101010001011;
    rom[2984] = 25'b0000000000000101010011000;
    rom[2985] = 25'b0000000000000101010100101;
    rom[2986] = 25'b0000000000000101010110010;
    rom[2987] = 25'b0000000000000101011000000;
    rom[2988] = 25'b0000000000000101011001100;
    rom[2989] = 25'b0000000000000101011011001;
    rom[2990] = 25'b0000000000000101011100111;
    rom[2991] = 25'b0000000000000101011110100;
    rom[2992] = 25'b0000000000000101100000000;
    rom[2993] = 25'b0000000000000101100001101;
    rom[2994] = 25'b0000000000000101100011010;
    rom[2995] = 25'b0000000000000101100100111;
    rom[2996] = 25'b0000000000000101100110011;
    rom[2997] = 25'b0000000000000101101000000;
    rom[2998] = 25'b0000000000000101101001101;
    rom[2999] = 25'b0000000000000101101011010;
    rom[3000] = 25'b0000000000000101101100110;
    rom[3001] = 25'b0000000000000101101110011;
    rom[3002] = 25'b0000000000000101110000000;
    rom[3003] = 25'b0000000000000101110001100;
    rom[3004] = 25'b0000000000000101110011001;
    rom[3005] = 25'b0000000000000101110100100;
    rom[3006] = 25'b0000000000000101110110001;
    rom[3007] = 25'b0000000000000101110111110;
    rom[3008] = 25'b0000000000000101111001010;
    rom[3009] = 25'b0000000000000101111010110;
    rom[3010] = 25'b0000000000000101111100011;
    rom[3011] = 25'b0000000000000101111101110;
    rom[3012] = 25'b0000000000000101111111010;
    rom[3013] = 25'b0000000000000110000000110;
    rom[3014] = 25'b0000000000000110000010011;
    rom[3015] = 25'b0000000000000110000011111;
    rom[3016] = 25'b0000000000000110000101011;
    rom[3017] = 25'b0000000000000110000110111;
    rom[3018] = 25'b0000000000000110001000011;
    rom[3019] = 25'b0000000000000110001001110;
    rom[3020] = 25'b0000000000000110001011010;
    rom[3021] = 25'b0000000000000110001100110;
    rom[3022] = 25'b0000000000000110001110001;
    rom[3023] = 25'b0000000000000110001111101;
    rom[3024] = 25'b0000000000000110010001000;
    rom[3025] = 25'b0000000000000110010010011;
    rom[3026] = 25'b0000000000000110010011111;
    rom[3027] = 25'b0000000000000110010101010;
    rom[3028] = 25'b0000000000000110010110110;
    rom[3029] = 25'b0000000000000110011000001;
    rom[3030] = 25'b0000000000000110011001100;
    rom[3031] = 25'b0000000000000110011011000;
    rom[3032] = 25'b0000000000000110011100011;
    rom[3033] = 25'b0000000000000110011101101;
    rom[3034] = 25'b0000000000000110011111000;
    rom[3035] = 25'b0000000000000110100000011;
    rom[3036] = 25'b0000000000000110100001110;
    rom[3037] = 25'b0000000000000110100011001;
    rom[3038] = 25'b0000000000000110100100011;
    rom[3039] = 25'b0000000000000110100101110;
    rom[3040] = 25'b0000000000000110100111000;
    rom[3041] = 25'b0000000000000110101000011;
    rom[3042] = 25'b0000000000000110101001110;
    rom[3043] = 25'b0000000000000110101011000;
    rom[3044] = 25'b0000000000000110101100010;
    rom[3045] = 25'b0000000000000110101101100;
    rom[3046] = 25'b0000000000000110101110111;
    rom[3047] = 25'b0000000000000110110000001;
    rom[3048] = 25'b0000000000000110110001011;
    rom[3049] = 25'b0000000000000110110010100;
    rom[3050] = 25'b0000000000000110110011111;
    rom[3051] = 25'b0000000000000110110101001;
    rom[3052] = 25'b0000000000000110110110010;
    rom[3053] = 25'b0000000000000110110111100;
    rom[3054] = 25'b0000000000000110111000110;
    rom[3055] = 25'b0000000000000110111001111;
    rom[3056] = 25'b0000000000000110111011000;
    rom[3057] = 25'b0000000000000110111100010;
    rom[3058] = 25'b0000000000000110111101011;
    rom[3059] = 25'b0000000000000110111110100;
    rom[3060] = 25'b0000000000000110111111110;
    rom[3061] = 25'b0000000000000111000000111;
    rom[3062] = 25'b0000000000000111000010000;
    rom[3063] = 25'b0000000000000111000011001;
    rom[3064] = 25'b0000000000000111000100010;
    rom[3065] = 25'b0000000000000111000101011;
    rom[3066] = 25'b0000000000000111000110011;
    rom[3067] = 25'b0000000000000111000111100;
    rom[3068] = 25'b0000000000000111001000100;
    rom[3069] = 25'b0000000000000111001001101;
    rom[3070] = 25'b0000000000000111001010101;
    rom[3071] = 25'b0000000000000111001011110;
    rom[3072] = 25'b0000000000000111001100110;
    rom[3073] = 25'b0000000000000111001101110;
    rom[3074] = 25'b0000000000000111001110110;
    rom[3075] = 25'b0000000000000111001111110;
    rom[3076] = 25'b0000000000000111010000110;
    rom[3077] = 25'b0000000000000111010001110;
    rom[3078] = 25'b0000000000000111010010101;
    rom[3079] = 25'b0000000000000111010011101;
    rom[3080] = 25'b0000000000000111010100100;
    rom[3081] = 25'b0000000000000111010101100;
    rom[3082] = 25'b0000000000000111010110100;
    rom[3083] = 25'b0000000000000111010111011;
    rom[3084] = 25'b0000000000000111011000010;
    rom[3085] = 25'b0000000000000111011001001;
    rom[3086] = 25'b0000000000000111011010000;
    rom[3087] = 25'b0000000000000111011010111;
    rom[3088] = 25'b0000000000000111011011101;
    rom[3089] = 25'b0000000000000111011100100;
    rom[3090] = 25'b0000000000000111011101011;
    rom[3091] = 25'b0000000000000111011110010;
    rom[3092] = 25'b0000000000000111011111000;
    rom[3093] = 25'b0000000000000111011111111;
    rom[3094] = 25'b0000000000000111100000101;
    rom[3095] = 25'b0000000000000111100001011;
    rom[3096] = 25'b0000000000000111100010001;
    rom[3097] = 25'b0000000000000111100010110;
    rom[3098] = 25'b0000000000000111100011100;
    rom[3099] = 25'b0000000000000111100100010;
    rom[3100] = 25'b0000000000000111100101000;
    rom[3101] = 25'b0000000000000111100101101;
    rom[3102] = 25'b0000000000000111100110011;
    rom[3103] = 25'b0000000000000111100111000;
    rom[3104] = 25'b0000000000000111100111110;
    rom[3105] = 25'b0000000000000111101000011;
    rom[3106] = 25'b0000000000000111101001000;
    rom[3107] = 25'b0000000000000111101001101;
    rom[3108] = 25'b0000000000000111101010010;
    rom[3109] = 25'b0000000000000111101010110;
    rom[3110] = 25'b0000000000000111101011011;
    rom[3111] = 25'b0000000000000111101100000;
    rom[3112] = 25'b0000000000000111101100100;
    rom[3113] = 25'b0000000000000111101101000;
    rom[3114] = 25'b0000000000000111101101100;
    rom[3115] = 25'b0000000000000111101110001;
    rom[3116] = 25'b0000000000000111101110101;
    rom[3117] = 25'b0000000000000111101111000;
    rom[3118] = 25'b0000000000000111101111100;
    rom[3119] = 25'b0000000000000111110000000;
    rom[3120] = 25'b0000000000000111110000011;
    rom[3121] = 25'b0000000000000111110000111;
    rom[3122] = 25'b0000000000000111110001010;
    rom[3123] = 25'b0000000000000111110001110;
    rom[3124] = 25'b0000000000000111110010000;
    rom[3125] = 25'b0000000000000111110010011;
    rom[3126] = 25'b0000000000000111110010110;
    rom[3127] = 25'b0000000000000111110011001;
    rom[3128] = 25'b0000000000000111110011011;
    rom[3129] = 25'b0000000000000111110011110;
    rom[3130] = 25'b0000000000000111110100000;
    rom[3131] = 25'b0000000000000111110100011;
    rom[3132] = 25'b0000000000000111110100100;
    rom[3133] = 25'b0000000000000111110100111;
    rom[3134] = 25'b0000000000000111110101001;
    rom[3135] = 25'b0000000000000111110101010;
    rom[3136] = 25'b0000000000000111110101100;
    rom[3137] = 25'b0000000000000111110101110;
    rom[3138] = 25'b0000000000000111110101111;
    rom[3139] = 25'b0000000000000111110110000;
    rom[3140] = 25'b0000000000000111110110001;
    rom[3141] = 25'b0000000000000111110110010;
    rom[3142] = 25'b0000000000000111110110011;
    rom[3143] = 25'b0000000000000111110110100;
    rom[3144] = 25'b0000000000000111110110101;
    rom[3145] = 25'b0000000000000111110110110;
    rom[3146] = 25'b0000000000000111110110110;
    rom[3147] = 25'b0000000000000111110110110;
    rom[3148] = 25'b0000000000000111110110110;
    rom[3149] = 25'b0000000000000111110110110;
    rom[3150] = 25'b0000000000000111110110110;
    rom[3151] = 25'b0000000000000111110110110;
    rom[3152] = 25'b0000000000000111110110110;
    rom[3153] = 25'b0000000000000111110110101;
    rom[3154] = 25'b0000000000000111110110101;
    rom[3155] = 25'b0000000000000111110110100;
    rom[3156] = 25'b0000000000000111110110011;
    rom[3157] = 25'b0000000000000111110110010;
    rom[3158] = 25'b0000000000000111110110000;
    rom[3159] = 25'b0000000000000111110110000;
    rom[3160] = 25'b0000000000000111110101110;
    rom[3161] = 25'b0000000000000111110101100;
    rom[3162] = 25'b0000000000000111110101010;
    rom[3163] = 25'b0000000000000111110101001;
    rom[3164] = 25'b0000000000000111110100111;
    rom[3165] = 25'b0000000000000111110100100;
    rom[3166] = 25'b0000000000000111110100011;
    rom[3167] = 25'b0000000000000111110100000;
    rom[3168] = 25'b0000000000000111110011110;
    rom[3169] = 25'b0000000000000111110011011;
    rom[3170] = 25'b0000000000000111110011000;
    rom[3171] = 25'b0000000000000111110010101;
    rom[3172] = 25'b0000000000000111110010010;
    rom[3173] = 25'b0000000000000111110001111;
    rom[3174] = 25'b0000000000000111110001100;
    rom[3175] = 25'b0000000000000111110001000;
    rom[3176] = 25'b0000000000000111110000100;
    rom[3177] = 25'b0000000000000111110000001;
    rom[3178] = 25'b0000000000000111101111101;
    rom[3179] = 25'b0000000000000111101111000;
    rom[3180] = 25'b0000000000000111101110101;
    rom[3181] = 25'b0000000000000111101110000;
    rom[3182] = 25'b0000000000000111101101100;
    rom[3183] = 25'b0000000000000111101100111;
    rom[3184] = 25'b0000000000000111101100010;
    rom[3185] = 25'b0000000000000111101011101;
    rom[3186] = 25'b0000000000000111101011000;
    rom[3187] = 25'b0000000000000111101010011;
    rom[3188] = 25'b0000000000000111101001110;
    rom[3189] = 25'b0000000000000111101001000;
    rom[3190] = 25'b0000000000000111101000011;
    rom[3191] = 25'b0000000000000111100111101;
    rom[3192] = 25'b0000000000000111100110111;
    rom[3193] = 25'b0000000000000111100110000;
    rom[3194] = 25'b0000000000000111100101010;
    rom[3195] = 25'b0000000000000111100100100;
    rom[3196] = 25'b0000000000000111100011101;
    rom[3197] = 25'b0000000000000111100010110;
    rom[3198] = 25'b0000000000000111100010000;
    rom[3199] = 25'b0000000000000111100001001;
    rom[3200] = 25'b0000000000000111100000001;
    rom[3201] = 25'b0000000000000111011111010;
    rom[3202] = 25'b0000000000000111011110011;
    rom[3203] = 25'b0000000000000111011101011;
    rom[3204] = 25'b0000000000000111011100011;
    rom[3205] = 25'b0000000000000111011011011;
    rom[3206] = 25'b0000000000000111011010011;
    rom[3207] = 25'b0000000000000111011001011;
    rom[3208] = 25'b0000000000000111011000010;
    rom[3209] = 25'b0000000000000111010111010;
    rom[3210] = 25'b0000000000000111010110001;
    rom[3211] = 25'b0000000000000111010101000;
    rom[3212] = 25'b0000000000000111010011111;
    rom[3213] = 25'b0000000000000111010010110;
    rom[3214] = 25'b0000000000000111010001101;
    rom[3215] = 25'b0000000000000111010000010;
    rom[3216] = 25'b0000000000000111001111001;
    rom[3217] = 25'b0000000000000111001101111;
    rom[3218] = 25'b0000000000000111001100110;
    rom[3219] = 25'b0000000000000111001011011;
    rom[3220] = 25'b0000000000000111001010001;
    rom[3221] = 25'b0000000000000111001000110;
    rom[3222] = 25'b0000000000000111000111100;
    rom[3223] = 25'b0000000000000111000110001;
    rom[3224] = 25'b0000000000000111000100110;
    rom[3225] = 25'b0000000000000111000011011;
    rom[3226] = 25'b0000000000000111000010000;
    rom[3227] = 25'b0000000000000111000000100;
    rom[3228] = 25'b0000000000000110111111001;
    rom[3229] = 25'b0000000000000110111101101;
    rom[3230] = 25'b0000000000000110111100001;
    rom[3231] = 25'b0000000000000110111010100;
    rom[3232] = 25'b0000000000000110111001000;
    rom[3233] = 25'b0000000000000110110111011;
    rom[3234] = 25'b0000000000000110110110000;
    rom[3235] = 25'b0000000000000110110100011;
    rom[3236] = 25'b0000000000000110110010101;
    rom[3237] = 25'b0000000000000110110001000;
    rom[3238] = 25'b0000000000000110101111011;
    rom[3239] = 25'b0000000000000110101101110;
    rom[3240] = 25'b0000000000000110101100000;
    rom[3241] = 25'b0000000000000110101010010;
    rom[3242] = 25'b0000000000000110101000100;
    rom[3243] = 25'b0000000000000110100110111;
    rom[3244] = 25'b0000000000000110100101000;
    rom[3245] = 25'b0000000000000110100011010;
    rom[3246] = 25'b0000000000000110100001011;
    rom[3247] = 25'b0000000000000110011111100;
    rom[3248] = 25'b0000000000000110011101110;
    rom[3249] = 25'b0000000000000110011011110;
    rom[3250] = 25'b0000000000000110011001111;
    rom[3251] = 25'b0000000000000110011000000;
    rom[3252] = 25'b0000000000000110010110000;
    rom[3253] = 25'b0000000000000110010100000;
    rom[3254] = 25'b0000000000000110010010000;
    rom[3255] = 25'b0000000000000110010000000;
    rom[3256] = 25'b0000000000000110001110000;
    rom[3257] = 25'b0000000000000110001100000;
    rom[3258] = 25'b0000000000000110001001111;
    rom[3259] = 25'b0000000000000110000111110;
    rom[3260] = 25'b0000000000000110000101101;
    rom[3261] = 25'b0000000000000110000011100;
    rom[3262] = 25'b0000000000000110000001011;
    rom[3263] = 25'b0000000000000101111111010;
    rom[3264] = 25'b0000000000000101111101000;
    rom[3265] = 25'b0000000000000101111010110;
    rom[3266] = 25'b0000000000000101111000100;
    rom[3267] = 25'b0000000000000101110110001;
    rom[3268] = 25'b0000000000000101110011111;
    rom[3269] = 25'b0000000000000101110001101;
    rom[3270] = 25'b0000000000000101101111010;
    rom[3271] = 25'b0000000000000101101100111;
    rom[3272] = 25'b0000000000000101101010101;
    rom[3273] = 25'b0000000000000101101000001;
    rom[3274] = 25'b0000000000000101100101101;
    rom[3275] = 25'b0000000000000101100011010;
    rom[3276] = 25'b0000000000000101100000110;
    rom[3277] = 25'b0000000000000101011110011;
    rom[3278] = 25'b0000000000000101011011110;
    rom[3279] = 25'b0000000000000101011001011;
    rom[3280] = 25'b0000000000000101010110110;
    rom[3281] = 25'b0000000000000101010100001;
    rom[3282] = 25'b0000000000000101010001101;
    rom[3283] = 25'b0000000000000101001111000;
    rom[3284] = 25'b0000000000000101001100011;
    rom[3285] = 25'b0000000000000101001001110;
    rom[3286] = 25'b0000000000000101000111000;
    rom[3287] = 25'b0000000000000101000100010;
    rom[3288] = 25'b0000000000000101000001101;
    rom[3289] = 25'b0000000000000100111110111;
    rom[3290] = 25'b0000000000000100111100001;
    rom[3291] = 25'b0000000000000100111001011;
    rom[3292] = 25'b0000000000000100110110100;
    rom[3293] = 25'b0000000000000100110011110;
    rom[3294] = 25'b0000000000000100110000111;
    rom[3295] = 25'b0000000000000100101110000;
    rom[3296] = 25'b0000000000000100101011001;
    rom[3297] = 25'b0000000000000100101000001;
    rom[3298] = 25'b0000000000000100100101010;
    rom[3299] = 25'b0000000000000100100010010;
    rom[3300] = 25'b0000000000000100011111010;
    rom[3301] = 25'b0000000000000100011100011;
    rom[3302] = 25'b0000000000000100011001010;
    rom[3303] = 25'b0000000000000100010110010;
    rom[3304] = 25'b0000000000000100010011001;
    rom[3305] = 25'b0000000000000100010000001;
    rom[3306] = 25'b0000000000000100001101000;
    rom[3307] = 25'b0000000000000100001001111;
    rom[3308] = 25'b0000000000000100000110101;
    rom[3309] = 25'b0000000000000100000011100;
    rom[3310] = 25'b0000000000000100000000011;
    rom[3311] = 25'b0000000000000011111101001;
    rom[3312] = 25'b0000000000000011111001111;
    rom[3313] = 25'b0000000000000011110110101;
    rom[3314] = 25'b0000000000000011110011011;
    rom[3315] = 25'b0000000000000011110000000;
    rom[3316] = 25'b0000000000000011101100110;
    rom[3317] = 25'b0000000000000011101001011;
    rom[3318] = 25'b0000000000000011100110000;
    rom[3319] = 25'b0000000000000011100010101;
    rom[3320] = 25'b0000000000000011011111010;
    rom[3321] = 25'b0000000000000011011011110;
    rom[3322] = 25'b0000000000000011011000011;
    rom[3323] = 25'b0000000000000011010100111;
    rom[3324] = 25'b0000000000000011010001011;
    rom[3325] = 25'b0000000000000011001101111;
    rom[3326] = 25'b0000000000000011001010011;
    rom[3327] = 25'b0000000000000011000110111;
    rom[3328] = 25'b0000000000000011000011010;
    rom[3329] = 25'b0000000000000010111111101;
    rom[3330] = 25'b0000000000000010111100000;
    rom[3331] = 25'b0000000000000010111000011;
    rom[3332] = 25'b0000000000000010110100110;
    rom[3333] = 25'b0000000000000010110001000;
    rom[3334] = 25'b0000000000000010101101011;
    rom[3335] = 25'b0000000000000010101001101;
    rom[3336] = 25'b0000000000000010100101111;
    rom[3337] = 25'b0000000000000010100010001;
    rom[3338] = 25'b0000000000000010011110011;
    rom[3339] = 25'b0000000000000010011010100;
    rom[3340] = 25'b0000000000000010010110110;
    rom[3341] = 25'b0000000000000010010010111;
    rom[3342] = 25'b0000000000000010001111000;
    rom[3343] = 25'b0000000000000010001011001;
    rom[3344] = 25'b0000000000000010000111010;
    rom[3345] = 25'b0000000000000010000011011;
    rom[3346] = 25'b0000000000000001111111011;
    rom[3347] = 25'b0000000000000001111011011;
    rom[3348] = 25'b0000000000000001110111011;
    rom[3349] = 25'b0000000000000001110011011;
    rom[3350] = 25'b0000000000000001101111011;
    rom[3351] = 25'b0000000000000001101011011;
    rom[3352] = 25'b0000000000000001100111010;
    rom[3353] = 25'b0000000000000001100011010;
    rom[3354] = 25'b0000000000000001011111001;
    rom[3355] = 25'b0000000000000001011011000;
    rom[3356] = 25'b0000000000000001010110110;
    rom[3357] = 25'b0000000000000001010010101;
    rom[3358] = 25'b0000000000000001001110100;
    rom[3359] = 25'b0000000000000001001010010;
    rom[3360] = 25'b0000000000000001000110001;
    rom[3361] = 25'b0000000000000001000001111;
    rom[3362] = 25'b0000000000000000111101101;
    rom[3363] = 25'b0000000000000000111001010;
    rom[3364] = 25'b0000000000000000110101000;
    rom[3365] = 25'b0000000000000000110000101;
    rom[3366] = 25'b0000000000000000101100010;
    rom[3367] = 25'b0000000000000000100111111;
    rom[3368] = 25'b0000000000000000100011100;
    rom[3369] = 25'b0000000000000000011111010;
    rom[3370] = 25'b0000000000000000011010110;
    rom[3371] = 25'b0000000000000000010110011;
    rom[3372] = 25'b0000000000000000010001111;
    rom[3373] = 25'b0000000000000000001101100;
    rom[3374] = 25'b0000000000000000001001000;
    rom[3375] = 25'b0000000000000000000100011;
    rom[3376] = 25'b0000000000000000000000000;
    rom[3377] = 25'b1111111111111111111011100;
    rom[3378] = 25'b1111111111111111110110111;
    rom[3379] = 25'b1111111111111111110010011;
    rom[3380] = 25'b1111111111111111101101101;
    rom[3381] = 25'b1111111111111111101001001;
    rom[3382] = 25'b1111111111111111100100011;
    rom[3383] = 25'b1111111111111111011111111;
    rom[3384] = 25'b1111111111111111011011001;
    rom[3385] = 25'b1111111111111111010110100;
    rom[3386] = 25'b1111111111111111010001110;
    rom[3387] = 25'b1111111111111111001101000;
    rom[3388] = 25'b1111111111111111001000010;
    rom[3389] = 25'b1111111111111111000011100;
    rom[3390] = 25'b1111111111111110111110101;
    rom[3391] = 25'b1111111111111110111001111;
    rom[3392] = 25'b1111111111111110110101001;
    rom[3393] = 25'b1111111111111110110000010;
    rom[3394] = 25'b1111111111111110101011011;
    rom[3395] = 25'b1111111111111110100110100;
    rom[3396] = 25'b1111111111111110100001101;
    rom[3397] = 25'b1111111111111110011100110;
    rom[3398] = 25'b1111111111111110010111111;
    rom[3399] = 25'b1111111111111110010011000;
    rom[3400] = 25'b1111111111111110001110000;
    rom[3401] = 25'b1111111111111110001001000;
    rom[3402] = 25'b1111111111111110000100000;
    rom[3403] = 25'b1111111111111101111111000;
    rom[3404] = 25'b1111111111111101111010000;
    rom[3405] = 25'b1111111111111101110101000;
    rom[3406] = 25'b1111111111111101110000000;
    rom[3407] = 25'b1111111111111101101010111;
    rom[3408] = 25'b1111111111111101100101110;
    rom[3409] = 25'b1111111111111101100000101;
    rom[3410] = 25'b1111111111111101011011101;
    rom[3411] = 25'b1111111111111101010110100;
    rom[3412] = 25'b1111111111111101010001011;
    rom[3413] = 25'b1111111111111101001100001;
    rom[3414] = 25'b1111111111111101000111000;
    rom[3415] = 25'b1111111111111101000001111;
    rom[3416] = 25'b1111111111111100111100101;
    rom[3417] = 25'b1111111111111100110111011;
    rom[3418] = 25'b1111111111111100110010010;
    rom[3419] = 25'b1111111111111100101100111;
    rom[3420] = 25'b1111111111111100100111110;
    rom[3421] = 25'b1111111111111100100010011;
    rom[3422] = 25'b1111111111111100011101001;
    rom[3423] = 25'b1111111111111100010111110;
    rom[3424] = 25'b1111111111111100010010011;
    rom[3425] = 25'b1111111111111100001101001;
    rom[3426] = 25'b1111111111111100000111110;
    rom[3427] = 25'b1111111111111100000010100;
    rom[3428] = 25'b1111111111111011111101001;
    rom[3429] = 25'b1111111111111011110111101;
    rom[3430] = 25'b1111111111111011110010011;
    rom[3431] = 25'b1111111111111011101100111;
    rom[3432] = 25'b1111111111111011100111100;
    rom[3433] = 25'b1111111111111011100010001;
    rom[3434] = 25'b1111111111111011011100100;
    rom[3435] = 25'b1111111111111011010111001;
    rom[3436] = 25'b1111111111111011010001101;
    rom[3437] = 25'b1111111111111011001100001;
    rom[3438] = 25'b1111111111111011000110101;
    rom[3439] = 25'b1111111111111011000001001;
    rom[3440] = 25'b1111111111111010111011101;
    rom[3441] = 25'b1111111111111010110110000;
    rom[3442] = 25'b1111111111111010110000100;
    rom[3443] = 25'b1111111111111010101010111;
    rom[3444] = 25'b1111111111111010100101011;
    rom[3445] = 25'b1111111111111010011111111;
    rom[3446] = 25'b1111111111111010011010010;
    rom[3447] = 25'b1111111111111010010100100;
    rom[3448] = 25'b1111111111111010001110111;
    rom[3449] = 25'b1111111111111010001001010;
    rom[3450] = 25'b1111111111111010000011101;
    rom[3451] = 25'b1111111111111001111110000;
    rom[3452] = 25'b1111111111111001111000011;
    rom[3453] = 25'b1111111111111001110010101;
    rom[3454] = 25'b1111111111111001101101000;
    rom[3455] = 25'b1111111111111001100111010;
    rom[3456] = 25'b1111111111111001100001101;
    rom[3457] = 25'b1111111111111001011011111;
    rom[3458] = 25'b1111111111111001010110001;
    rom[3459] = 25'b1111111111111001010000011;
    rom[3460] = 25'b1111111111111001001010101;
    rom[3461] = 25'b1111111111111001000100111;
    rom[3462] = 25'b1111111111111000111111010;
    rom[3463] = 25'b1111111111111000111001100;
    rom[3464] = 25'b1111111111111000110011110;
    rom[3465] = 25'b1111111111111000101101111;
    rom[3466] = 25'b1111111111111000101000001;
    rom[3467] = 25'b1111111111111000100010010;
    rom[3468] = 25'b1111111111111000011100011;
    rom[3469] = 25'b1111111111111000010110110;
    rom[3470] = 25'b1111111111111000010000111;
    rom[3471] = 25'b1111111111111000001011000;
    rom[3472] = 25'b1111111111111000000101001;
    rom[3473] = 25'b1111111111110111111111010;
    rom[3474] = 25'b1111111111110111111001100;
    rom[3475] = 25'b1111111111110111110011101;
    rom[3476] = 25'b1111111111110111101101101;
    rom[3477] = 25'b1111111111110111100111110;
    rom[3478] = 25'b1111111111110111100010000;
    rom[3479] = 25'b1111111111110111011100000;
    rom[3480] = 25'b1111111111110111010110001;
    rom[3481] = 25'b1111111111110111010000010;
    rom[3482] = 25'b1111111111110111001010011;
    rom[3483] = 25'b1111111111110111000100011;
    rom[3484] = 25'b1111111111110110111110100;
    rom[3485] = 25'b1111111111110110111000101;
    rom[3486] = 25'b1111111111110110110010101;
    rom[3487] = 25'b1111111111110110101100110;
    rom[3488] = 25'b1111111111110110100110110;
    rom[3489] = 25'b1111111111110110100000110;
    rom[3490] = 25'b1111111111110110011010111;
    rom[3491] = 25'b1111111111110110010100111;
    rom[3492] = 25'b1111111111110110001110111;
    rom[3493] = 25'b1111111111110110001001000;
    rom[3494] = 25'b1111111111110110000011000;
    rom[3495] = 25'b1111111111110101111101001;
    rom[3496] = 25'b1111111111110101110111001;
    rom[3497] = 25'b1111111111110101110001000;
    rom[3498] = 25'b1111111111110101101011001;
    rom[3499] = 25'b1111111111110101100101001;
    rom[3500] = 25'b1111111111110101011111010;
    rom[3501] = 25'b1111111111110101011001001;
    rom[3502] = 25'b1111111111110101010011001;
    rom[3503] = 25'b1111111111110101001101001;
    rom[3504] = 25'b1111111111110101000111001;
    rom[3505] = 25'b1111111111110101000001010;
    rom[3506] = 25'b1111111111110100111011001;
    rom[3507] = 25'b1111111111110100110101010;
    rom[3508] = 25'b1111111111110100101111001;
    rom[3509] = 25'b1111111111110100101001001;
    rom[3510] = 25'b1111111111110100100011001;
    rom[3511] = 25'b1111111111110100011101001;
    rom[3512] = 25'b1111111111110100010111001;
    rom[3513] = 25'b1111111111110100010001001;
    rom[3514] = 25'b1111111111110100001011001;
    rom[3515] = 25'b1111111111110100000101001;
    rom[3516] = 25'b1111111111110011111111001;
    rom[3517] = 25'b1111111111110011111001001;
    rom[3518] = 25'b1111111111110011110011001;
    rom[3519] = 25'b1111111111110011101101001;
    rom[3520] = 25'b1111111111110011100111000;
    rom[3521] = 25'b1111111111110011100001001;
    rom[3522] = 25'b1111111111110011011011000;
    rom[3523] = 25'b1111111111110011010101001;
    rom[3524] = 25'b1111111111110011001111000;
    rom[3525] = 25'b1111111111110011001001001;
    rom[3526] = 25'b1111111111110011000011001;
    rom[3527] = 25'b1111111111110010111101001;
    rom[3528] = 25'b1111111111110010110111001;
    rom[3529] = 25'b1111111111110010110001001;
    rom[3530] = 25'b1111111111110010101011001;
    rom[3531] = 25'b1111111111110010100101001;
    rom[3532] = 25'b1111111111110010011111010;
    rom[3533] = 25'b1111111111110010011001010;
    rom[3534] = 25'b1111111111110010010011001;
    rom[3535] = 25'b1111111111110010001101010;
    rom[3536] = 25'b1111111111110010000111010;
    rom[3537] = 25'b1111111111110010000001011;
    rom[3538] = 25'b1111111111110001111011011;
    rom[3539] = 25'b1111111111110001110101011;
    rom[3540] = 25'b1111111111110001101111100;
    rom[3541] = 25'b1111111111110001101001100;
    rom[3542] = 25'b1111111111110001100011101;
    rom[3543] = 25'b1111111111110001011101110;
    rom[3544] = 25'b1111111111110001010111110;
    rom[3545] = 25'b1111111111110001010001111;
    rom[3546] = 25'b1111111111110001001100000;
    rom[3547] = 25'b1111111111110001000110000;
    rom[3548] = 25'b1111111111110001000000001;
    rom[3549] = 25'b1111111111110000111010010;
    rom[3550] = 25'b1111111111110000110100011;
    rom[3551] = 25'b1111111111110000101110100;
    rom[3552] = 25'b1111111111110000101000101;
    rom[3553] = 25'b1111111111110000100010110;
    rom[3554] = 25'b1111111111110000011101000;
    rom[3555] = 25'b1111111111110000010111001;
    rom[3556] = 25'b1111111111110000010001010;
    rom[3557] = 25'b1111111111110000001011011;
    rom[3558] = 25'b1111111111110000000101101;
    rom[3559] = 25'b1111111111101111111111111;
    rom[3560] = 25'b1111111111101111111010000;
    rom[3561] = 25'b1111111111101111110100010;
    rom[3562] = 25'b1111111111101111101110011;
    rom[3563] = 25'b1111111111101111101000101;
    rom[3564] = 25'b1111111111101111100010111;
    rom[3565] = 25'b1111111111101111011101001;
    rom[3566] = 25'b1111111111101111010111011;
    rom[3567] = 25'b1111111111101111010001110;
    rom[3568] = 25'b1111111111101111001100000;
    rom[3569] = 25'b1111111111101111000110010;
    rom[3570] = 25'b1111111111101111000000101;
    rom[3571] = 25'b1111111111101110111010111;
    rom[3572] = 25'b1111111111101110110101010;
    rom[3573] = 25'b1111111111101110101111101;
    rom[3574] = 25'b1111111111101110101001111;
    rom[3575] = 25'b1111111111101110100100010;
    rom[3576] = 25'b1111111111101110011110101;
    rom[3577] = 25'b1111111111101110011001000;
    rom[3578] = 25'b1111111111101110010011011;
    rom[3579] = 25'b1111111111101110001101111;
    rom[3580] = 25'b1111111111101110001000011;
    rom[3581] = 25'b1111111111101110000010110;
    rom[3582] = 25'b1111111111101101111101001;
    rom[3583] = 25'b1111111111101101110111101;
    rom[3584] = 25'b1111111111101101110010001;
    rom[3585] = 25'b1111111111101101101100110;
    rom[3586] = 25'b1111111111101101100111001;
    rom[3587] = 25'b1111111111101101100001110;
    rom[3588] = 25'b1111111111101101011100011;
    rom[3589] = 25'b1111111111101101010110111;
    rom[3590] = 25'b1111111111101101010001100;
    rom[3591] = 25'b1111111111101101001100000;
    rom[3592] = 25'b1111111111101101000110101;
    rom[3593] = 25'b1111111111101101000001011;
    rom[3594] = 25'b1111111111101100111011111;
    rom[3595] = 25'b1111111111101100110110101;
    rom[3596] = 25'b1111111111101100110001010;
    rom[3597] = 25'b1111111111101100101100000;
    rom[3598] = 25'b1111111111101100100110110;
    rom[3599] = 25'b1111111111101100100001011;
    rom[3600] = 25'b1111111111101100011100010;
    rom[3601] = 25'b1111111111101100010111000;
    rom[3602] = 25'b1111111111101100010001110;
    rom[3603] = 25'b1111111111101100001100101;
    rom[3604] = 25'b1111111111101100000111100;
    rom[3605] = 25'b1111111111101100000010010;
    rom[3606] = 25'b1111111111101011111101001;
    rom[3607] = 25'b1111111111101011111000001;
    rom[3608] = 25'b1111111111101011110011000;
    rom[3609] = 25'b1111111111101011101110000;
    rom[3610] = 25'b1111111111101011101000111;
    rom[3611] = 25'b1111111111101011100011111;
    rom[3612] = 25'b1111111111101011011110111;
    rom[3613] = 25'b1111111111101011011001111;
    rom[3614] = 25'b1111111111101011010101000;
    rom[3615] = 25'b1111111111101011010000000;
    rom[3616] = 25'b1111111111101011001011001;
    rom[3617] = 25'b1111111111101011000110010;
    rom[3618] = 25'b1111111111101011000001011;
    rom[3619] = 25'b1111111111101010111100100;
    rom[3620] = 25'b1111111111101010110111110;
    rom[3621] = 25'b1111111111101010110010111;
    rom[3622] = 25'b1111111111101010101110001;
    rom[3623] = 25'b1111111111101010101001011;
    rom[3624] = 25'b1111111111101010100100110;
    rom[3625] = 25'b1111111111101010100000000;
    rom[3626] = 25'b1111111111101010011011010;
    rom[3627] = 25'b1111111111101010010110110;
    rom[3628] = 25'b1111111111101010010010000;
    rom[3629] = 25'b1111111111101010001101100;
    rom[3630] = 25'b1111111111101010001000111;
    rom[3631] = 25'b1111111111101010000100010;
    rom[3632] = 25'b1111111111101001111111111;
    rom[3633] = 25'b1111111111101001111011011;
    rom[3634] = 25'b1111111111101001110110111;
    rom[3635] = 25'b1111111111101001110010011;
    rom[3636] = 25'b1111111111101001101110000;
    rom[3637] = 25'b1111111111101001101001101;
    rom[3638] = 25'b1111111111101001100101010;
    rom[3639] = 25'b1111111111101001100000111;
    rom[3640] = 25'b1111111111101001011100101;
    rom[3641] = 25'b1111111111101001011000011;
    rom[3642] = 25'b1111111111101001010100001;
    rom[3643] = 25'b1111111111101001001111111;
    rom[3644] = 25'b1111111111101001001011110;
    rom[3645] = 25'b1111111111101001000111101;
    rom[3646] = 25'b1111111111101001000011100;
    rom[3647] = 25'b1111111111101000111111011;
    rom[3648] = 25'b1111111111101000111011010;
    rom[3649] = 25'b1111111111101000110111011;
    rom[3650] = 25'b1111111111101000110011010;
    rom[3651] = 25'b1111111111101000101111011;
    rom[3652] = 25'b1111111111101000101011011;
    rom[3653] = 25'b1111111111101000100111100;
    rom[3654] = 25'b1111111111101000100011100;
    rom[3655] = 25'b1111111111101000011111110;
    rom[3656] = 25'b1111111111101000011011111;
    rom[3657] = 25'b1111111111101000011000001;
    rom[3658] = 25'b1111111111101000010100011;
    rom[3659] = 25'b1111111111101000010000110;
    rom[3660] = 25'b1111111111101000001101000;
    rom[3661] = 25'b1111111111101000001001011;
    rom[3662] = 25'b1111111111101000000101110;
    rom[3663] = 25'b1111111111101000000010001;
    rom[3664] = 25'b1111111111100111111110101;
    rom[3665] = 25'b1111111111100111111011001;
    rom[3666] = 25'b1111111111100111110111101;
    rom[3667] = 25'b1111111111100111110100010;
    rom[3668] = 25'b1111111111100111110000111;
    rom[3669] = 25'b1111111111100111101101100;
    rom[3670] = 25'b1111111111100111101010001;
    rom[3671] = 25'b1111111111100111100110110;
    rom[3672] = 25'b1111111111100111100011100;
    rom[3673] = 25'b1111111111100111100000010;
    rom[3674] = 25'b1111111111100111011101001;
    rom[3675] = 25'b1111111111100111011010000;
    rom[3676] = 25'b1111111111100111010110111;
    rom[3677] = 25'b1111111111100111010011111;
    rom[3678] = 25'b1111111111100111010000110;
    rom[3679] = 25'b1111111111100111001101110;
    rom[3680] = 25'b1111111111100111001010110;
    rom[3681] = 25'b1111111111100111000111110;
    rom[3682] = 25'b1111111111100111000100111;
    rom[3683] = 25'b1111111111100111000010001;
    rom[3684] = 25'b1111111111100110111111010;
    rom[3685] = 25'b1111111111100110111100100;
    rom[3686] = 25'b1111111111100110111001110;
    rom[3687] = 25'b1111111111100110110111001;
    rom[3688] = 25'b1111111111100110110100100;
    rom[3689] = 25'b1111111111100110110001111;
    rom[3690] = 25'b1111111111100110101111010;
    rom[3691] = 25'b1111111111100110101100110;
    rom[3692] = 25'b1111111111100110101010010;
    rom[3693] = 25'b1111111111100110100111110;
    rom[3694] = 25'b1111111111100110100101100;
    rom[3695] = 25'b1111111111100110100011000;
    rom[3696] = 25'b1111111111100110100000101;
    rom[3697] = 25'b1111111111100110011110100;
    rom[3698] = 25'b1111111111100110011100010;
    rom[3699] = 25'b1111111111100110011010000;
    rom[3700] = 25'b1111111111100110010111111;
    rom[3701] = 25'b1111111111100110010101110;
    rom[3702] = 25'b1111111111100110010011110;
    rom[3703] = 25'b1111111111100110010001110;
    rom[3704] = 25'b1111111111100110001111101;
    rom[3705] = 25'b1111111111100110001101110;
    rom[3706] = 25'b1111111111100110001011111;
    rom[3707] = 25'b1111111111100110001010000;
    rom[3708] = 25'b1111111111100110001000010;
    rom[3709] = 25'b1111111111100110000110100;
    rom[3710] = 25'b1111111111100110000100110;
    rom[3711] = 25'b1111111111100110000011001;
    rom[3712] = 25'b1111111111100110000001100;
    rom[3713] = 25'b1111111111100110000000000;
    rom[3714] = 25'b1111111111100101111110011;
    rom[3715] = 25'b1111111111100101111100111;
    rom[3716] = 25'b1111111111100101111011100;
    rom[3717] = 25'b1111111111100101111010001;
    rom[3718] = 25'b1111111111100101111000110;
    rom[3719] = 25'b1111111111100101110111011;
    rom[3720] = 25'b1111111111100101110110001;
    rom[3721] = 25'b1111111111100101110101000;
    rom[3722] = 25'b1111111111100101110011111;
    rom[3723] = 25'b1111111111100101110010110;
    rom[3724] = 25'b1111111111100101110001110;
    rom[3725] = 25'b1111111111100101110000110;
    rom[3726] = 25'b1111111111100101101111110;
    rom[3727] = 25'b1111111111100101101110111;
    rom[3728] = 25'b1111111111100101101110000;
    rom[3729] = 25'b1111111111100101101101001;
    rom[3730] = 25'b1111111111100101101100011;
    rom[3731] = 25'b1111111111100101101011110;
    rom[3732] = 25'b1111111111100101101011000;
    rom[3733] = 25'b1111111111100101101010100;
    rom[3734] = 25'b1111111111100101101001111;
    rom[3735] = 25'b1111111111100101101001011;
    rom[3736] = 25'b1111111111100101101000111;
    rom[3737] = 25'b1111111111100101101000100;
    rom[3738] = 25'b1111111111100101101000001;
    rom[3739] = 25'b1111111111100101100111110;
    rom[3740] = 25'b1111111111100101100111101;
    rom[3741] = 25'b1111111111100101100111011;
    rom[3742] = 25'b1111111111100101100111010;
    rom[3743] = 25'b1111111111100101100111001;
    rom[3744] = 25'b1111111111100101100111000;
    rom[3745] = 25'b1111111111100101100111000;
    rom[3746] = 25'b1111111111100101100111001;
    rom[3747] = 25'b1111111111100101100111010;
    rom[3748] = 25'b1111111111100101100111100;
    rom[3749] = 25'b1111111111100101100111110;
    rom[3750] = 25'b1111111111100101100111111;
    rom[3751] = 25'b1111111111100101101000010;
    rom[3752] = 25'b1111111111100101101000101;
    rom[3753] = 25'b1111111111100101101001001;
    rom[3754] = 25'b1111111111100101101001101;
    rom[3755] = 25'b1111111111100101101010001;
    rom[3756] = 25'b1111111111100101101010101;
    rom[3757] = 25'b1111111111100101101011011;
    rom[3758] = 25'b1111111111100101101100000;
    rom[3759] = 25'b1111111111100101101100110;
    rom[3760] = 25'b1111111111100101101101101;
    rom[3761] = 25'b1111111111100101101110100;
    rom[3762] = 25'b1111111111100101101111100;
    rom[3763] = 25'b1111111111100101110000100;
    rom[3764] = 25'b1111111111100101110001100;
    rom[3765] = 25'b1111111111100101110010101;
    rom[3766] = 25'b1111111111100101110011111;
    rom[3767] = 25'b1111111111100101110101000;
    rom[3768] = 25'b1111111111100101110110010;
    rom[3769] = 25'b1111111111100101110111101;
    rom[3770] = 25'b1111111111100101111001000;
    rom[3771] = 25'b1111111111100101111010011;
    rom[3772] = 25'b1111111111100101111011111;
    rom[3773] = 25'b1111111111100101111101100;
    rom[3774] = 25'b1111111111100101111111001;
    rom[3775] = 25'b1111111111100110000000110;
    rom[3776] = 25'b1111111111100110000010100;
    rom[3777] = 25'b1111111111100110000100010;
    rom[3778] = 25'b1111111111100110000110010;
    rom[3779] = 25'b1111111111100110001000001;
    rom[3780] = 25'b1111111111100110001010000;
    rom[3781] = 25'b1111111111100110001100000;
    rom[3782] = 25'b1111111111100110001110001;
    rom[3783] = 25'b1111111111100110010000010;
    rom[3784] = 25'b1111111111100110010010100;
    rom[3785] = 25'b1111111111100110010100110;
    rom[3786] = 25'b1111111111100110010111001;
    rom[3787] = 25'b1111111111100110011001100;
    rom[3788] = 25'b1111111111100110011100000;
    rom[3789] = 25'b1111111111100110011110100;
    rom[3790] = 25'b1111111111100110100001000;
    rom[3791] = 25'b1111111111100110100011101;
    rom[3792] = 25'b1111111111100110100110011;
    rom[3793] = 25'b1111111111100110101001001;
    rom[3794] = 25'b1111111111100110101100000;
    rom[3795] = 25'b1111111111100110101110111;
    rom[3796] = 25'b1111111111100110110001110;
    rom[3797] = 25'b1111111111100110110100110;
    rom[3798] = 25'b1111111111100110110111110;
    rom[3799] = 25'b1111111111100110111011000;
    rom[3800] = 25'b1111111111100110111110001;
    rom[3801] = 25'b1111111111100111000001011;
    rom[3802] = 25'b1111111111100111000100101;
    rom[3803] = 25'b1111111111100111001000000;
    rom[3804] = 25'b1111111111100111001011011;
    rom[3805] = 25'b1111111111100111001110111;
    rom[3806] = 25'b1111111111100111010010100;
    rom[3807] = 25'b1111111111100111010110001;
    rom[3808] = 25'b1111111111100111011001110;
    rom[3809] = 25'b1111111111100111011101100;
    rom[3810] = 25'b1111111111100111100001011;
    rom[3811] = 25'b1111111111100111100101010;
    rom[3812] = 25'b1111111111100111101001001;
    rom[3813] = 25'b1111111111100111101101001;
    rom[3814] = 25'b1111111111100111110001010;
    rom[3815] = 25'b1111111111100111110101010;
    rom[3816] = 25'b1111111111100111111001100;
    rom[3817] = 25'b1111111111100111111101110;
    rom[3818] = 25'b1111111111101000000010001;
    rom[3819] = 25'b1111111111101000000110100;
    rom[3820] = 25'b1111111111101000001010111;
    rom[3821] = 25'b1111111111101000001111100;
    rom[3822] = 25'b1111111111101000010100000;
    rom[3823] = 25'b1111111111101000011000110;
    rom[3824] = 25'b1111111111101000011101011;
    rom[3825] = 25'b1111111111101000100010001;
    rom[3826] = 25'b1111111111101000100111000;
    rom[3827] = 25'b1111111111101000101011111;
    rom[3828] = 25'b1111111111101000110000111;
    rom[3829] = 25'b1111111111101000110101111;
    rom[3830] = 25'b1111111111101000111011000;
    rom[3831] = 25'b1111111111101001000000001;
    rom[3832] = 25'b1111111111101001000101011;
    rom[3833] = 25'b1111111111101001001010101;
    rom[3834] = 25'b1111111111101001010000000;
    rom[3835] = 25'b1111111111101001010101011;
    rom[3836] = 25'b1111111111101001011011000;
    rom[3837] = 25'b1111111111101001100000100;
    rom[3838] = 25'b1111111111101001100110001;
    rom[3839] = 25'b1111111111101001101011110;
    rom[3840] = 25'b1111111111101001110001100;
    rom[3841] = 25'b1111111111101001110111011;
    rom[3842] = 25'b1111111111101001111101001;
    rom[3843] = 25'b1111111111101010000011001;
    rom[3844] = 25'b1111111111101010001001001;
    rom[3845] = 25'b1111111111101010001111010;
    rom[3846] = 25'b1111111111101010010101011;
    rom[3847] = 25'b1111111111101010011011101;
    rom[3848] = 25'b1111111111101010100001111;
    rom[3849] = 25'b1111111111101010101000010;
    rom[3850] = 25'b1111111111101010101110101;
    rom[3851] = 25'b1111111111101010110101001;
    rom[3852] = 25'b1111111111101010111011101;
    rom[3853] = 25'b1111111111101011000010010;
    rom[3854] = 25'b1111111111101011001001000;
    rom[3855] = 25'b1111111111101011001111110;
    rom[3856] = 25'b1111111111101011010110101;
    rom[3857] = 25'b1111111111101011011101011;
    rom[3858] = 25'b1111111111101011100100011;
    rom[3859] = 25'b1111111111101011101011011;
    rom[3860] = 25'b1111111111101011110010011;
    rom[3861] = 25'b1111111111101011111001101;
    rom[3862] = 25'b1111111111101100000000110;
    rom[3863] = 25'b1111111111101100001000001;
    rom[3864] = 25'b1111111111101100001111100;
    rom[3865] = 25'b1111111111101100010110111;
    rom[3866] = 25'b1111111111101100011110011;
    rom[3867] = 25'b1111111111101100100101111;
    rom[3868] = 25'b1111111111101100101101100;
    rom[3869] = 25'b1111111111101100110101010;
    rom[3870] = 25'b1111111111101100111101000;
    rom[3871] = 25'b1111111111101101000100110;
    rom[3872] = 25'b1111111111101101001100110;
    rom[3873] = 25'b1111111111101101010100100;
    rom[3874] = 25'b1111111111101101011100101;
    rom[3875] = 25'b1111111111101101100100110;
    rom[3876] = 25'b1111111111101101101100111;
    rom[3877] = 25'b1111111111101101110101001;
    rom[3878] = 25'b1111111111101101111101011;
    rom[3879] = 25'b1111111111101110000101101;
    rom[3880] = 25'b1111111111101110001110001;
    rom[3881] = 25'b1111111111101110010110101;
    rom[3882] = 25'b1111111111101110011111010;
    rom[3883] = 25'b1111111111101110100111110;
    rom[3884] = 25'b1111111111101110110000100;
    rom[3885] = 25'b1111111111101110111001010;
    rom[3886] = 25'b1111111111101111000010001;
    rom[3887] = 25'b1111111111101111001011000;
    rom[3888] = 25'b1111111111101111010011111;
    rom[3889] = 25'b1111111111101111011101000;
    rom[3890] = 25'b1111111111101111100110000;
    rom[3891] = 25'b1111111111101111101111001;
    rom[3892] = 25'b1111111111101111111000011;
    rom[3893] = 25'b1111111111110000000001110;
    rom[3894] = 25'b1111111111110000001011001;
    rom[3895] = 25'b1111111111110000010100100;
    rom[3896] = 25'b1111111111110000011101111;
    rom[3897] = 25'b1111111111110000100111100;
    rom[3898] = 25'b1111111111110000110001001;
    rom[3899] = 25'b1111111111110000111010111;
    rom[3900] = 25'b1111111111110001000100101;
    rom[3901] = 25'b1111111111110001001110011;
    rom[3902] = 25'b1111111111110001011000010;
    rom[3903] = 25'b1111111111110001100010001;
    rom[3904] = 25'b1111111111110001101100010;
    rom[3905] = 25'b1111111111110001110110011;
    rom[3906] = 25'b1111111111110010000000100;
    rom[3907] = 25'b1111111111110010001010101;
    rom[3908] = 25'b1111111111110010010101000;
    rom[3909] = 25'b1111111111110010011111010;
    rom[3910] = 25'b1111111111110010101001110;
    rom[3911] = 25'b1111111111110010110100010;
    rom[3912] = 25'b1111111111110010111110110;
    rom[3913] = 25'b1111111111110011001001010;
    rom[3914] = 25'b1111111111110011010100000;
    rom[3915] = 25'b1111111111110011011110110;
    rom[3916] = 25'b1111111111110011101001100;
    rom[3917] = 25'b1111111111110011110100100;
    rom[3918] = 25'b1111111111110011111111010;
    rom[3919] = 25'b1111111111110100001010011;
    rom[3920] = 25'b1111111111110100010101011;
    rom[3921] = 25'b1111111111110100100000100;
    rom[3922] = 25'b1111111111110100101011110;
    rom[3923] = 25'b1111111111110100110111000;
    rom[3924] = 25'b1111111111110101000010010;
    rom[3925] = 25'b1111111111110101001101101;
    rom[3926] = 25'b1111111111110101011001001;
    rom[3927] = 25'b1111111111110101100100101;
    rom[3928] = 25'b1111111111110101110000010;
    rom[3929] = 25'b1111111111110101111011110;
    rom[3930] = 25'b1111111111110110000111100;
    rom[3931] = 25'b1111111111110110010011010;
    rom[3932] = 25'b1111111111110110011111001;
    rom[3933] = 25'b1111111111110110101011000;
    rom[3934] = 25'b1111111111110110110110111;
    rom[3935] = 25'b1111111111110111000010111;
    rom[3936] = 25'b1111111111110111001111000;
    rom[3937] = 25'b1111111111110111011011001;
    rom[3938] = 25'b1111111111110111100111011;
    rom[3939] = 25'b1111111111110111110011101;
    rom[3940] = 25'b1111111111111000000000000;
    rom[3941] = 25'b1111111111111000001100010;
    rom[3942] = 25'b1111111111111000011000110;
    rom[3943] = 25'b1111111111111000100101010;
    rom[3944] = 25'b1111111111111000110001110;
    rom[3945] = 25'b1111111111111000111110100;
    rom[3946] = 25'b1111111111111001001011001;
    rom[3947] = 25'b1111111111111001010111111;
    rom[3948] = 25'b1111111111111001100100110;
    rom[3949] = 25'b1111111111111001110001101;
    rom[3950] = 25'b1111111111111001111110100;
    rom[3951] = 25'b1111111111111010001011011;
    rom[3952] = 25'b1111111111111010011000100;
    rom[3953] = 25'b1111111111111010100101101;
    rom[3954] = 25'b1111111111111010110010110;
    rom[3955] = 25'b1111111111111011000000000;
    rom[3956] = 25'b1111111111111011001101011;
    rom[3957] = 25'b1111111111111011011010101;
    rom[3958] = 25'b1111111111111011101000000;
    rom[3959] = 25'b1111111111111011110101100;
    rom[3960] = 25'b1111111111111100000011000;
    rom[3961] = 25'b1111111111111100010000101;
    rom[3962] = 25'b1111111111111100011110010;
    rom[3963] = 25'b1111111111111100101100000;
    rom[3964] = 25'b1111111111111100111001101;
    rom[3965] = 25'b1111111111111101000111100;
    rom[3966] = 25'b1111111111111101010101010;
    rom[3967] = 25'b1111111111111101100011010;
    rom[3968] = 25'b1111111111111101110001010;
    rom[3969] = 25'b1111111111111101111111010;
    rom[3970] = 25'b1111111111111110001101011;
    rom[3971] = 25'b1111111111111110011011100;
    rom[3972] = 25'b1111111111111110101001110;
    rom[3973] = 25'b1111111111111110111000000;
    rom[3974] = 25'b1111111111111111000110010;
    rom[3975] = 25'b1111111111111111010100100;
    rom[3976] = 25'b1111111111111111100011000;
    rom[3977] = 25'b1111111111111111110001100;
    rom[3978] = 25'b0000000000000000000000000;
    rom[3979] = 25'b0000000000000000001110100;
    rom[3980] = 25'b0000000000000000011101001;
    rom[3981] = 25'b0000000000000000101011110;
    rom[3982] = 25'b0000000000000000111010100;
    rom[3983] = 25'b0000000000000001001001010;
    rom[3984] = 25'b0000000000000001011000001;
    rom[3985] = 25'b0000000000000001100111000;
    rom[3986] = 25'b0000000000000001110110000;
    rom[3987] = 25'b0000000000000010000100111;
    rom[3988] = 25'b0000000000000010010100000;
    rom[3989] = 25'b0000000000000010100011001;
    rom[3990] = 25'b0000000000000010110010010;
    rom[3991] = 25'b0000000000000011000001011;
    rom[3992] = 25'b0000000000000011010000101;
    rom[3993] = 25'b0000000000000011011111111;
    rom[3994] = 25'b0000000000000011101111011;
    rom[3995] = 25'b0000000000000011111110101;
    rom[3996] = 25'b0000000000000100001110001;
    rom[3997] = 25'b0000000000000100011101101;
    rom[3998] = 25'b0000000000000100101101001;
    rom[3999] = 25'b0000000000000100111100110;
    rom[4000] = 25'b0000000000000101001100011;
    rom[4001] = 25'b0000000000000101011100001;
    rom[4002] = 25'b0000000000000101101011111;
    rom[4003] = 25'b0000000000000101111011101;
    rom[4004] = 25'b0000000000000110001011011;
    rom[4005] = 25'b0000000000000110011011010;
    rom[4006] = 25'b0000000000000110101011010;
    rom[4007] = 25'b0000000000000110111011001;
    rom[4008] = 25'b0000000000000111001011001;
    rom[4009] = 25'b0000000000000111011011001;
    rom[4010] = 25'b0000000000000111101011010;
    rom[4011] = 25'b0000000000000111111011011;
    rom[4012] = 25'b0000000000001000001011100;
    rom[4013] = 25'b0000000000001000011011110;
    rom[4014] = 25'b0000000000001000101100000;
    rom[4015] = 25'b0000000000001000111100011;
    rom[4016] = 25'b0000000000001001001100110;
    rom[4017] = 25'b0000000000001001011101001;
    rom[4018] = 25'b0000000000001001101101100;
    rom[4019] = 25'b0000000000001001111101111;
    rom[4020] = 25'b0000000000001010001110100;
    rom[4021] = 25'b0000000000001010011111000;
    rom[4022] = 25'b0000000000001010101111101;
    rom[4023] = 25'b0000000000001011000000010;
    rom[4024] = 25'b0000000000001011010001000;
    rom[4025] = 25'b0000000000001011100001101;
    rom[4026] = 25'b0000000000001011110010011;
    rom[4027] = 25'b0000000000001100000011001;
    rom[4028] = 25'b0000000000001100010011111;
    rom[4029] = 25'b0000000000001100100100111;
    rom[4030] = 25'b0000000000001100110101110;
    rom[4031] = 25'b0000000000001101000110101;
    rom[4032] = 25'b0000000000001101010111100;
    rom[4033] = 25'b0000000000001101101000100;
    rom[4034] = 25'b0000000000001101111001101;
    rom[4035] = 25'b0000000000001110001010101;
    rom[4036] = 25'b0000000000001110011011110;
    rom[4037] = 25'b0000000000001110101100111;
    rom[4038] = 25'b0000000000001110111110001;
    rom[4039] = 25'b0000000000001111001111010;
    rom[4040] = 25'b0000000000001111100000101;
    rom[4041] = 25'b0000000000001111110001110;
    rom[4042] = 25'b0000000000010000000011001;
    rom[4043] = 25'b0000000000010000010100100;
    rom[4044] = 25'b0000000000010000100101110;
    rom[4045] = 25'b0000000000010000110111010;
    rom[4046] = 25'b0000000000010001001000101;
    rom[4047] = 25'b0000000000010001011010001;
    rom[4048] = 25'b0000000000010001101011100;
    rom[4049] = 25'b0000000000010001111101001;
    rom[4050] = 25'b0000000000010010001110101;
    rom[4051] = 25'b0000000000010010100000001;
    rom[4052] = 25'b0000000000010010110001110;
    rom[4053] = 25'b0000000000010011000011011;
    rom[4054] = 25'b0000000000010011010101000;
    rom[4055] = 25'b0000000000010011100110101;
    rom[4056] = 25'b0000000000010011111000011;
    rom[4057] = 25'b0000000000010100001010000;
    rom[4058] = 25'b0000000000010100011011110;
    rom[4059] = 25'b0000000000010100101101100;
    rom[4060] = 25'b0000000000010100111111011;
    rom[4061] = 25'b0000000000010101010001001;
    rom[4062] = 25'b0000000000010101100011000;
    rom[4063] = 25'b0000000000010101110100111;
    rom[4064] = 25'b0000000000010110000110110;
    rom[4065] = 25'b0000000000010110011000110;
    rom[4066] = 25'b0000000000010110101010101;
    rom[4067] = 25'b0000000000010110111100100;
    rom[4068] = 25'b0000000000010111001110100;
    rom[4069] = 25'b0000000000010111100000100;
    rom[4070] = 25'b0000000000010111110010100;
    rom[4071] = 25'b0000000000011000000100100;
    rom[4072] = 25'b0000000000011000010110101;
    rom[4073] = 25'b0000000000011000101000101;
    rom[4074] = 25'b0000000000011000111010110;
    rom[4075] = 25'b0000000000011001001100110;
    rom[4076] = 25'b0000000000011001011110111;
    rom[4077] = 25'b0000000000011001110001000;
    rom[4078] = 25'b0000000000011010000011001;
    rom[4079] = 25'b0000000000011010010101010;
    rom[4080] = 25'b0000000000011010100111100;
    rom[4081] = 25'b0000000000011010111001100;
    rom[4082] = 25'b0000000000011011001011111;
    rom[4083] = 25'b0000000000011011011110000;
    rom[4084] = 25'b0000000000011011110000010;
    rom[4085] = 25'b0000000000011100000010011;
    rom[4086] = 25'b0000000000011100010100101;
    rom[4087] = 25'b0000000000011100100110111;
    rom[4088] = 25'b0000000000011100111001001;
    rom[4089] = 25'b0000000000011101001011011;
    rom[4090] = 25'b0000000000011101011101110;
    rom[4091] = 25'b0000000000011101110000000;
    rom[4092] = 25'b0000000000011110000010010;
    rom[4093] = 25'b0000000000011110010100100;
    rom[4094] = 25'b0000000000011110100110111;
    rom[4095] = 25'b0000000000011110111001001;
    rom[4096] = 25'b0000000000011111001011011;
    rom[4097] = 25'b0000000000011111011101110;
    rom[4098] = 25'b0000000000011111110000000;
    rom[4099] = 25'b0000000000100000000010011;
    rom[4100] = 25'b0000000000100000010100101;
    rom[4101] = 25'b0000000000100000100111000;
    rom[4102] = 25'b0000000000100000111001011;
    rom[4103] = 25'b0000000000100001001011101;
    rom[4104] = 25'b0000000000100001011110000;
    rom[4105] = 25'b0000000000100001110000010;
    rom[4106] = 25'b0000000000100010000010101;
    rom[4107] = 25'b0000000000100010010101000;
    rom[4108] = 25'b0000000000100010100111010;
    rom[4109] = 25'b0000000000100010111001100;
    rom[4110] = 25'b0000000000100011001100000;
    rom[4111] = 25'b0000000000100011011110010;
    rom[4112] = 25'b0000000000100011110000100;
    rom[4113] = 25'b0000000000100100000010110;
    rom[4114] = 25'b0000000000100100010101001;
    rom[4115] = 25'b0000000000100100100111011;
    rom[4116] = 25'b0000000000100100111001101;
    rom[4117] = 25'b0000000000100101001100000;
    rom[4118] = 25'b0000000000100101011110010;
    rom[4119] = 25'b0000000000100101110000100;
    rom[4120] = 25'b0000000000100110000010110;
    rom[4121] = 25'b0000000000100110010101000;
    rom[4122] = 25'b0000000000100110100111010;
    rom[4123] = 25'b0000000000100110111001100;
    rom[4124] = 25'b0000000000100111001011101;
    rom[4125] = 25'b0000000000100111011101111;
    rom[4126] = 25'b0000000000100111110000001;
    rom[4127] = 25'b0000000000101000000010010;
    rom[4128] = 25'b0000000000101000010100011;
    rom[4129] = 25'b0000000000101000100110100;
    rom[4130] = 25'b0000000000101000111000110;
    rom[4131] = 25'b0000000000101001001010110;
    rom[4132] = 25'b0000000000101001011100111;
    rom[4133] = 25'b0000000000101001101110111;
    rom[4134] = 25'b0000000000101010000001000;
    rom[4135] = 25'b0000000000101010010011001;
    rom[4136] = 25'b0000000000101010100101001;
    rom[4137] = 25'b0000000000101010110111001;
    rom[4138] = 25'b0000000000101011001001001;
    rom[4139] = 25'b0000000000101011011011000;
    rom[4140] = 25'b0000000000101011101101000;
    rom[4141] = 25'b0000000000101011111111000;
    rom[4142] = 25'b0000000000101100010000111;
    rom[4143] = 25'b0000000000101100100010110;
    rom[4144] = 25'b0000000000101100110100100;
    rom[4145] = 25'b0000000000101101000110011;
    rom[4146] = 25'b0000000000101101011000001;
    rom[4147] = 25'b0000000000101101101010000;
    rom[4148] = 25'b0000000000101101111011110;
    rom[4149] = 25'b0000000000101110001101100;
    rom[4150] = 25'b0000000000101110011111010;
    rom[4151] = 25'b0000000000101110110000111;
    rom[4152] = 25'b0000000000101111000010100;
    rom[4153] = 25'b0000000000101111010100001;
    rom[4154] = 25'b0000000000101111100101101;
    rom[4155] = 25'b0000000000101111110111010;
    rom[4156] = 25'b0000000000110000001000110;
    rom[4157] = 25'b0000000000110000011010010;
    rom[4158] = 25'b0000000000110000101011101;
    rom[4159] = 25'b0000000000110000111101001;
    rom[4160] = 25'b0000000000110001001110100;
    rom[4161] = 25'b0000000000110001011111111;
    rom[4162] = 25'b0000000000110001110001001;
    rom[4163] = 25'b0000000000110010000010011;
    rom[4164] = 25'b0000000000110010010011101;
    rom[4165] = 25'b0000000000110010100100111;
    rom[4166] = 25'b0000000000110010110110000;
    rom[4167] = 25'b0000000000110011000111001;
    rom[4168] = 25'b0000000000110011011000001;
    rom[4169] = 25'b0000000000110011101001010;
    rom[4170] = 25'b0000000000110011111010010;
    rom[4171] = 25'b0000000000110100001011010;
    rom[4172] = 25'b0000000000110100011100001;
    rom[4173] = 25'b0000000000110100101101000;
    rom[4174] = 25'b0000000000110100111101111;
    rom[4175] = 25'b0000000000110101001110101;
    rom[4176] = 25'b0000000000110101011111011;
    rom[4177] = 25'b0000000000110101110000001;
    rom[4178] = 25'b0000000000110110000000110;
    rom[4179] = 25'b0000000000110110010001011;
    rom[4180] = 25'b0000000000110110100010000;
    rom[4181] = 25'b0000000000110110110010011;
    rom[4182] = 25'b0000000000110111000010111;
    rom[4183] = 25'b0000000000110111010011010;
    rom[4184] = 25'b0000000000110111100011101;
    rom[4185] = 25'b0000000000110111110011111;
    rom[4186] = 25'b0000000000111000000100010;
    rom[4187] = 25'b0000000000111000010100100;
    rom[4188] = 25'b0000000000111000100100100;
    rom[4189] = 25'b0000000000111000110100101;
    rom[4190] = 25'b0000000000111001000100110;
    rom[4191] = 25'b0000000000111001010100101;
    rom[4192] = 25'b0000000000111001100100101;
    rom[4193] = 25'b0000000000111001110100100;
    rom[4194] = 25'b0000000000111010000100010;
    rom[4195] = 25'b0000000000111010010100000;
    rom[4196] = 25'b0000000000111010100011110;
    rom[4197] = 25'b0000000000111010110011011;
    rom[4198] = 25'b0000000000111011000010111;
    rom[4199] = 25'b0000000000111011010010011;
    rom[4200] = 25'b0000000000111011100010000;
    rom[4201] = 25'b0000000000111011110001011;
    rom[4202] = 25'b0000000000111100000000101;
    rom[4203] = 25'b0000000000111100001111111;
    rom[4204] = 25'b0000000000111100011111001;
    rom[4205] = 25'b0000000000111100101110010;
    rom[4206] = 25'b0000000000111100111101010;
    rom[4207] = 25'b0000000000111101001100011;
    rom[4208] = 25'b0000000000111101011011010;
    rom[4209] = 25'b0000000000111101101010001;
    rom[4210] = 25'b0000000000111101111000111;
    rom[4211] = 25'b0000000000111110000111110;
    rom[4212] = 25'b0000000000111110010110011;
    rom[4213] = 25'b0000000000111110100100111;
    rom[4214] = 25'b0000000000111110110011011;
    rom[4215] = 25'b0000000000111111000001111;
    rom[4216] = 25'b0000000000111111010000010;
    rom[4217] = 25'b0000000000111111011110100;
    rom[4218] = 25'b0000000000111111101100110;
    rom[4219] = 25'b0000000000111111111011000;
    rom[4220] = 25'b0000000001000000001001000;
    rom[4221] = 25'b0000000001000000010111000;
    rom[4222] = 25'b0000000001000000100100111;
    rom[4223] = 25'b0000000001000000110010110;
    rom[4224] = 25'b0000000001000001000000101;
    rom[4225] = 25'b0000000001000001001110001;
    rom[4226] = 25'b0000000001000001011011110;
    rom[4227] = 25'b0000000001000001101001010;
    rom[4228] = 25'b0000000001000001110110110;
    rom[4229] = 25'b0000000001000010000100010;
    rom[4230] = 25'b0000000001000010010001011;
    rom[4231] = 25'b0000000001000010011110101;
    rom[4232] = 25'b0000000001000010101011110;
    rom[4233] = 25'b0000000001000010111000110;
    rom[4234] = 25'b0000000001000011000101101;
    rom[4235] = 25'b0000000001000011010010100;
    rom[4236] = 25'b0000000001000011011111010;
    rom[4237] = 25'b0000000001000011101100000;
    rom[4238] = 25'b0000000001000011111000101;
    rom[4239] = 25'b0000000001000100000101000;
    rom[4240] = 25'b0000000001000100010001100;
    rom[4241] = 25'b0000000001000100011101110;
    rom[4242] = 25'b0000000001000100101010000;
    rom[4243] = 25'b0000000001000100110110001;
    rom[4244] = 25'b0000000001000101000010010;
    rom[4245] = 25'b0000000001000101001110001;
    rom[4246] = 25'b0000000001000101011010001;
    rom[4247] = 25'b0000000001000101100101110;
    rom[4248] = 25'b0000000001000101110001100;
    rom[4249] = 25'b0000000001000101111101001;
    rom[4250] = 25'b0000000001000110001000100;
    rom[4251] = 25'b0000000001000110010011111;
    rom[4252] = 25'b0000000001000110011111010;
    rom[4253] = 25'b0000000001000110101010011;
    rom[4254] = 25'b0000000001000110110101011;
    rom[4255] = 25'b0000000001000111000000100;
    rom[4256] = 25'b0000000001000111001011010;
    rom[4257] = 25'b0000000001000111010110000;
    rom[4258] = 25'b0000000001000111100000110;
    rom[4259] = 25'b0000000001000111101011010;
    rom[4260] = 25'b0000000001000111110101111;
    rom[4261] = 25'b0000000001001000000000001;
    rom[4262] = 25'b0000000001001000001010100;
    rom[4263] = 25'b0000000001001000010100100;
    rom[4264] = 25'b0000000001001000011110101;
    rom[4265] = 25'b0000000001001000101000101;
    rom[4266] = 25'b0000000001001000110010011;
    rom[4267] = 25'b0000000001001000111100010;
    rom[4268] = 25'b0000000001001001000101110;
    rom[4269] = 25'b0000000001001001001111010;
    rom[4270] = 25'b0000000001001001011000110;
    rom[4271] = 25'b0000000001001001100010000;
    rom[4272] = 25'b0000000001001001101011010;
    rom[4273] = 25'b0000000001001001110100010;
    rom[4274] = 25'b0000000001001001111101001;
    rom[4275] = 25'b0000000001001010000110000;
    rom[4276] = 25'b0000000001001010001110110;
    rom[4277] = 25'b0000000001001010010111011;
    rom[4278] = 25'b0000000001001010011111111;
    rom[4279] = 25'b0000000001001010101000010;
    rom[4280] = 25'b0000000001001010110000011;
    rom[4281] = 25'b0000000001001010111000101;
    rom[4282] = 25'b0000000001001011000000101;
    rom[4283] = 25'b0000000001001011001000100;
    rom[4284] = 25'b0000000001001011010000010;
    rom[4285] = 25'b0000000001001011011000000;
    rom[4286] = 25'b0000000001001011011111100;
    rom[4287] = 25'b0000000001001011100111000;
    rom[4288] = 25'b0000000001001011101110001;
    rom[4289] = 25'b0000000001001011110101011;
    rom[4290] = 25'b0000000001001011111100011;
    rom[4291] = 25'b0000000001001100000011011;
    rom[4292] = 25'b0000000001001100001010001;
    rom[4293] = 25'b0000000001001100010000111;
    rom[4294] = 25'b0000000001001100010111011;
    rom[4295] = 25'b0000000001001100011101110;
    rom[4296] = 25'b0000000001001100100100001;
    rom[4297] = 25'b0000000001001100101010010;
    rom[4298] = 25'b0000000001001100110000010;
    rom[4299] = 25'b0000000001001100110110001;
    rom[4300] = 25'b0000000001001100111100000;
    rom[4301] = 25'b0000000001001101000001101;
    rom[4302] = 25'b0000000001001101000111001;
    rom[4303] = 25'b0000000001001101001100100;
    rom[4304] = 25'b0000000001001101010001110;
    rom[4305] = 25'b0000000001001101010110111;
    rom[4306] = 25'b0000000001001101011011111;
    rom[4307] = 25'b0000000001001101100000110;
    rom[4308] = 25'b0000000001001101100101100;
    rom[4309] = 25'b0000000001001101101010000;
    rom[4310] = 25'b0000000001001101101110100;
    rom[4311] = 25'b0000000001001101110010110;
    rom[4312] = 25'b0000000001001101110111000;
    rom[4313] = 25'b0000000001001101111011000;
    rom[4314] = 25'b0000000001001101111110111;
    rom[4315] = 25'b0000000001001110000010101;
    rom[4316] = 25'b0000000001001110000110010;
    rom[4317] = 25'b0000000001001110001001110;
    rom[4318] = 25'b0000000001001110001101000;
    rom[4319] = 25'b0000000001001110010000010;
    rom[4320] = 25'b0000000001001110010011010;
    rom[4321] = 25'b0000000001001110010110001;
    rom[4322] = 25'b0000000001001110011000111;
    rom[4323] = 25'b0000000001001110011011101;
    rom[4324] = 25'b0000000001001110011110000;
    rom[4325] = 25'b0000000001001110100000011;
    rom[4326] = 25'b0000000001001110100010101;
    rom[4327] = 25'b0000000001001110100100101;
    rom[4328] = 25'b0000000001001110100110100;
    rom[4329] = 25'b0000000001001110101000010;
    rom[4330] = 25'b0000000001001110101001111;
    rom[4331] = 25'b0000000001001110101011010;
    rom[4332] = 25'b0000000001001110101100101;
    rom[4333] = 25'b0000000001001110101101110;
    rom[4334] = 25'b0000000001001110101110110;
    rom[4335] = 25'b0000000001001110101111101;
    rom[4336] = 25'b0000000001001110110000010;
    rom[4337] = 25'b0000000001001110110000111;
    rom[4338] = 25'b0000000001001110110001010;
    rom[4339] = 25'b0000000001001110110001100;
    rom[4340] = 25'b0000000001001110110001101;
    rom[4341] = 25'b0000000001001110110001100;
    rom[4342] = 25'b0000000001001110110001010;
    rom[4343] = 25'b0000000001001110110000111;
    rom[4344] = 25'b0000000001001110110000010;
    rom[4345] = 25'b0000000001001110101111101;
    rom[4346] = 25'b0000000001001110101110111;
    rom[4347] = 25'b0000000001001110101101111;
    rom[4348] = 25'b0000000001001110101100110;
    rom[4349] = 25'b0000000001001110101011010;
    rom[4350] = 25'b0000000001001110101001111;
    rom[4351] = 25'b0000000001001110101000010;
    rom[4352] = 25'b0000000001001110100110011;
    rom[4353] = 25'b0000000001001110100100100;
    rom[4354] = 25'b0000000001001110100010011;
    rom[4355] = 25'b0000000001001110100000001;
    rom[4356] = 25'b0000000001001110011101110;
    rom[4357] = 25'b0000000001001110011011000;
    rom[4358] = 25'b0000000001001110011000010;
    rom[4359] = 25'b0000000001001110010101011;
    rom[4360] = 25'b0000000001001110010010011;
    rom[4361] = 25'b0000000001001110001111000;
    rom[4362] = 25'b0000000001001110001011101;
    rom[4363] = 25'b0000000001001110001000001;
    rom[4364] = 25'b0000000001001110000100011;
    rom[4365] = 25'b0000000001001110000000100;
    rom[4366] = 25'b0000000001001101111100011;
    rom[4367] = 25'b0000000001001101111000001;
    rom[4368] = 25'b0000000001001101110011110;
    rom[4369] = 25'b0000000001001101101111001;
    rom[4370] = 25'b0000000001001101101010100;
    rom[4371] = 25'b0000000001001101100101100;
    rom[4372] = 25'b0000000001001101100000100;
    rom[4373] = 25'b0000000001001101011011001;
    rom[4374] = 25'b0000000001001101010101110;
    rom[4375] = 25'b0000000001001101010000010;
    rom[4376] = 25'b0000000001001101001010100;
    rom[4377] = 25'b0000000001001101000100100;
    rom[4378] = 25'b0000000001001100111110100;
    rom[4379] = 25'b0000000001001100111000001;
    rom[4380] = 25'b0000000001001100110001110;
    rom[4381] = 25'b0000000001001100101011001;
    rom[4382] = 25'b0000000001001100100100010;
    rom[4383] = 25'b0000000001001100011101011;
    rom[4384] = 25'b0000000001001100010110010;
    rom[4385] = 25'b0000000001001100001110111;
    rom[4386] = 25'b0000000001001100000111100;
    rom[4387] = 25'b0000000001001011111111111;
    rom[4388] = 25'b0000000001001011111000000;
    rom[4389] = 25'b0000000001001011110000000;
    rom[4390] = 25'b0000000001001011100111110;
    rom[4391] = 25'b0000000001001011011111011;
    rom[4392] = 25'b0000000001001011010110111;
    rom[4393] = 25'b0000000001001011001110001;
    rom[4394] = 25'b0000000001001011000101011;
    rom[4395] = 25'b0000000001001010111100011;
    rom[4396] = 25'b0000000001001010110011001;
    rom[4397] = 25'b0000000001001010101001101;
    rom[4398] = 25'b0000000001001010100000000;
    rom[4399] = 25'b0000000001001010010110010;
    rom[4400] = 25'b0000000001001010001100011;
    rom[4401] = 25'b0000000001001010000010001;
    rom[4402] = 25'b0000000001001001110111111;
    rom[4403] = 25'b0000000001001001101101100;
    rom[4404] = 25'b0000000001001001100010110;
    rom[4405] = 25'b0000000001001001011000000;
    rom[4406] = 25'b0000000001001001001100111;
    rom[4407] = 25'b0000000001001001000001101;
    rom[4408] = 25'b0000000001001000110110010;
    rom[4409] = 25'b0000000001001000101010110;
    rom[4410] = 25'b0000000001001000011111000;
    rom[4411] = 25'b0000000001001000010011001;
    rom[4412] = 25'b0000000001001000000111000;
    rom[4413] = 25'b0000000001000111111010101;
    rom[4414] = 25'b0000000001000111101110001;
    rom[4415] = 25'b0000000001000111100001100;
    rom[4416] = 25'b0000000001000111010100101;
    rom[4417] = 25'b0000000001000111000111110;
    rom[4418] = 25'b0000000001000110111010100;
    rom[4419] = 25'b0000000001000110101101001;
    rom[4420] = 25'b0000000001000110011111100;
    rom[4421] = 25'b0000000001000110010001110;
    rom[4422] = 25'b0000000001000110000011111;
    rom[4423] = 25'b0000000001000101110101110;
    rom[4424] = 25'b0000000001000101100111011;
    rom[4425] = 25'b0000000001000101011000111;
    rom[4426] = 25'b0000000001000101001010010;
    rom[4427] = 25'b0000000001000100111011011;
    rom[4428] = 25'b0000000001000100101100011;
    rom[4429] = 25'b0000000001000100011101001;
    rom[4430] = 25'b0000000001000100001101101;
    rom[4431] = 25'b0000000001000011111110001;
    rom[4432] = 25'b0000000001000011101110010;
    rom[4433] = 25'b0000000001000011011110011;
    rom[4434] = 25'b0000000001000011001110001;
    rom[4435] = 25'b0000000001000010111101110;
    rom[4436] = 25'b0000000001000010101101011;
    rom[4437] = 25'b0000000001000010011100101;
    rom[4438] = 25'b0000000001000010001011110;
    rom[4439] = 25'b0000000001000001111010101;
    rom[4440] = 25'b0000000001000001101001010;
    rom[4441] = 25'b0000000001000001010111111;
    rom[4442] = 25'b0000000001000001000110010;
    rom[4443] = 25'b0000000001000000110100011;
    rom[4444] = 25'b0000000001000000100010011;
    rom[4445] = 25'b0000000001000000010000010;
    rom[4446] = 25'b0000000000111111111101110;
    rom[4447] = 25'b0000000000111111101011010;
    rom[4448] = 25'b0000000000111111011000011;
    rom[4449] = 25'b0000000000111111000101100;
    rom[4450] = 25'b0000000000111110110010011;
    rom[4451] = 25'b0000000000111110011111000;
    rom[4452] = 25'b0000000000111110001011100;
    rom[4453] = 25'b0000000000111101110111110;
    rom[4454] = 25'b0000000000111101100011111;
    rom[4455] = 25'b0000000000111101001111110;
    rom[4456] = 25'b0000000000111100111011101;
    rom[4457] = 25'b0000000000111100100111000;
    rom[4458] = 25'b0000000000111100010010011;
    rom[4459] = 25'b0000000000111011111101101;
    rom[4460] = 25'b0000000000111011101000101;
    rom[4461] = 25'b0000000000111011010011011;
    rom[4462] = 25'b0000000000111010111110000;
    rom[4463] = 25'b0000000000111010101000100;
    rom[4464] = 25'b0000000000111010010010110;
    rom[4465] = 25'b0000000000111001111100110;
    rom[4466] = 25'b0000000000111001100110101;
    rom[4467] = 25'b0000000000111001010000010;
    rom[4468] = 25'b0000000000111000111001110;
    rom[4469] = 25'b0000000000111000100011001;
    rom[4470] = 25'b0000000000111000001100010;
    rom[4471] = 25'b0000000000110111110101010;
    rom[4472] = 25'b0000000000110111011101111;
    rom[4473] = 25'b0000000000110111000110011;
    rom[4474] = 25'b0000000000110110101110111;
    rom[4475] = 25'b0000000000110110010111000;
    rom[4476] = 25'b0000000000110101111111000;
    rom[4477] = 25'b0000000000110101100110111;
    rom[4478] = 25'b0000000000110101001110100;
    rom[4479] = 25'b0000000000110100110110000;
    rom[4480] = 25'b0000000000110100011101001;
    rom[4481] = 25'b0000000000110100000100010;
    rom[4482] = 25'b0000000000110011101011001;
    rom[4483] = 25'b0000000000110011010001110;
    rom[4484] = 25'b0000000000110010111000011;
    rom[4485] = 25'b0000000000110010011110101;
    rom[4486] = 25'b0000000000110010000100111;
    rom[4487] = 25'b0000000000110001101010110;
    rom[4488] = 25'b0000000000110001010000101;
    rom[4489] = 25'b0000000000110000110110001;
    rom[4490] = 25'b0000000000110000011011101;
    rom[4491] = 25'b0000000000110000000000111;
    rom[4492] = 25'b0000000000101111100101111;
    rom[4493] = 25'b0000000000101111001010110;
    rom[4494] = 25'b0000000000101110101111100;
    rom[4495] = 25'b0000000000101110010011111;
    rom[4496] = 25'b0000000000101101111000010;
    rom[4497] = 25'b0000000000101101011100011;
    rom[4498] = 25'b0000000000101101000000011;
    rom[4499] = 25'b0000000000101100100100001;
    rom[4500] = 25'b0000000000101100000111110;
    rom[4501] = 25'b0000000000101011101011001;
    rom[4502] = 25'b0000000000101011001110010;
    rom[4503] = 25'b0000000000101010110001011;
    rom[4504] = 25'b0000000000101010010100010;
    rom[4505] = 25'b0000000000101001110110111;
    rom[4506] = 25'b0000000000101001011001100;
    rom[4507] = 25'b0000000000101000111011110;
    rom[4508] = 25'b0000000000101000011101111;
    rom[4509] = 25'b0000000000100111111111111;
    rom[4510] = 25'b0000000000100111100001110;
    rom[4511] = 25'b0000000000100111000011011;
    rom[4512] = 25'b0000000000100110100100110;
    rom[4513] = 25'b0000000000100110000110000;
    rom[4514] = 25'b0000000000100101100111000;
    rom[4515] = 25'b0000000000100101001000000;
    rom[4516] = 25'b0000000000100100101000110;
    rom[4517] = 25'b0000000000100100001001010;
    rom[4518] = 25'b0000000000100011101001110;
    rom[4519] = 25'b0000000000100011001001111;
    rom[4520] = 25'b0000000000100010101001111;
    rom[4521] = 25'b0000000000100010001001111;
    rom[4522] = 25'b0000000000100001101001100;
    rom[4523] = 25'b0000000000100001001001000;
    rom[4524] = 25'b0000000000100000101000011;
    rom[4525] = 25'b0000000000100000000111100;
    rom[4526] = 25'b0000000000011111100110011;
    rom[4527] = 25'b0000000000011111000101010;
    rom[4528] = 25'b0000000000011110100100000;
    rom[4529] = 25'b0000000000011110000010011;
    rom[4530] = 25'b0000000000011101100000101;
    rom[4531] = 25'b0000000000011100111110111;
    rom[4532] = 25'b0000000000011100011100111;
    rom[4533] = 25'b0000000000011011111010101;
    rom[4534] = 25'b0000000000011011011000010;
    rom[4535] = 25'b0000000000011010110101110;
    rom[4536] = 25'b0000000000011010010011001;
    rom[4537] = 25'b0000000000011001110000010;
    rom[4538] = 25'b0000000000011001001101001;
    rom[4539] = 25'b0000000000011000101001111;
    rom[4540] = 25'b0000000000011000000110101;
    rom[4541] = 25'b0000000000010111100011000;
    rom[4542] = 25'b0000000000010110111111011;
    rom[4543] = 25'b0000000000010110011011100;
    rom[4544] = 25'b0000000000010101110111100;
    rom[4545] = 25'b0000000000010101010011010;
    rom[4546] = 25'b0000000000010100101111000;
    rom[4547] = 25'b0000000000010100001010100;
    rom[4548] = 25'b0000000000010011100101110;
    rom[4549] = 25'b0000000000010011000001000;
    rom[4550] = 25'b0000000000010010011100000;
    rom[4551] = 25'b0000000000010001110110111;
    rom[4552] = 25'b0000000000010001010001101;
    rom[4553] = 25'b0000000000010000101100001;
    rom[4554] = 25'b0000000000010000000110100;
    rom[4555] = 25'b0000000000001111100000110;
    rom[4556] = 25'b0000000000001110111010111;
    rom[4557] = 25'b0000000000001110010100110;
    rom[4558] = 25'b0000000000001101101110100;
    rom[4559] = 25'b0000000000001101001000001;
    rom[4560] = 25'b0000000000001100100001101;
    rom[4561] = 25'b0000000000001011111011000;
    rom[4562] = 25'b0000000000001011010100000;
    rom[4563] = 25'b0000000000001010101101001;
    rom[4564] = 25'b0000000000001010000101111;
    rom[4565] = 25'b0000000000001001011110101;
    rom[4566] = 25'b0000000000001000110111010;
    rom[4567] = 25'b0000000000001000001111101;
    rom[4568] = 25'b0000000000000111100111111;
    rom[4569] = 25'b0000000000000111000000000;
    rom[4570] = 25'b0000000000000110011000000;
    rom[4571] = 25'b0000000000000101101111110;
    rom[4572] = 25'b0000000000000101000111100;
    rom[4573] = 25'b0000000000000100011111000;
    rom[4574] = 25'b0000000000000011110110100;
    rom[4575] = 25'b0000000000000011001101101;
    rom[4576] = 25'b0000000000000010100100111;
    rom[4577] = 25'b0000000000000001111011110;
    rom[4578] = 25'b0000000000000001010010101;
    rom[4579] = 25'b0000000000000000101001010;
    rom[4580] = 25'b0000000000000000000000000;
    rom[4581] = 25'b1111111111111111010110011;
    rom[4582] = 25'b1111111111111110101100110;
    rom[4583] = 25'b1111111111111110000010110;
    rom[4584] = 25'b1111111111111101011000111;
    rom[4585] = 25'b1111111111111100101110110;
    rom[4586] = 25'b1111111111111100000100100;
    rom[4587] = 25'b1111111111111011011010001;
    rom[4588] = 25'b1111111111111010101111101;
    rom[4589] = 25'b1111111111111010000101000;
    rom[4590] = 25'b1111111111111001011010010;
    rom[4591] = 25'b1111111111111000101111011;
    rom[4592] = 25'b1111111111111000000100010;
    rom[4593] = 25'b1111111111110111011001001;
    rom[4594] = 25'b1111111111110110101101111;
    rom[4595] = 25'b1111111111110110000010100;
    rom[4596] = 25'b1111111111110101010111000;
    rom[4597] = 25'b1111111111110100101011011;
    rom[4598] = 25'b1111111111110011111111100;
    rom[4599] = 25'b1111111111110011010011101;
    rom[4600] = 25'b1111111111110010100111110;
    rom[4601] = 25'b1111111111110001111011100;
    rom[4602] = 25'b1111111111110001001111010;
    rom[4603] = 25'b1111111111110000100010111;
    rom[4604] = 25'b1111111111101111110110100;
    rom[4605] = 25'b1111111111101111001001111;
    rom[4606] = 25'b1111111111101110011101001;
    rom[4607] = 25'b1111111111101101110000010;
    rom[4608] = 25'b1111111111101101000011011;
    rom[4609] = 25'b1111111111101100010110011;
    rom[4610] = 25'b1111111111101011101001001;
    rom[4611] = 25'b1111111111101010111011111;
    rom[4612] = 25'b1111111111101010001110101;
    rom[4613] = 25'b1111111111101001100001001;
    rom[4614] = 25'b1111111111101000110011100;
    rom[4615] = 25'b1111111111101000000101110;
    rom[4616] = 25'b1111111111100111011000001;
    rom[4617] = 25'b1111111111100110101010001;
    rom[4618] = 25'b1111111111100101111100001;
    rom[4619] = 25'b1111111111100101001110001;
    rom[4620] = 25'b1111111111100100011111111;
    rom[4621] = 25'b1111111111100011110001101;
    rom[4622] = 25'b1111111111100011000011010;
    rom[4623] = 25'b1111111111100010010100101;
    rom[4624] = 25'b1111111111100001100110001;
    rom[4625] = 25'b1111111111100000110111011;
    rom[4626] = 25'b1111111111100000001000101;
    rom[4627] = 25'b1111111111011111011001111;
    rom[4628] = 25'b1111111111011110101010111;
    rom[4629] = 25'b1111111111011101111011111;
    rom[4630] = 25'b1111111111011101001100110;
    rom[4631] = 25'b1111111111011100011101100;
    rom[4632] = 25'b1111111111011011101110001;
    rom[4633] = 25'b1111111111011010111110111;
    rom[4634] = 25'b1111111111011010001111011;
    rom[4635] = 25'b1111111111011001011111111;
    rom[4636] = 25'b1111111111011000110000010;
    rom[4637] = 25'b1111111111011000000000100;
    rom[4638] = 25'b1111111111010111010000110;
    rom[4639] = 25'b1111111111010110100000111;
    rom[4640] = 25'b1111111111010101110001000;
    rom[4641] = 25'b1111111111010101000000111;
    rom[4642] = 25'b1111111111010100010000111;
    rom[4643] = 25'b1111111111010011100000101;
    rom[4644] = 25'b1111111111010010110000011;
    rom[4645] = 25'b1111111111010010000000001;
    rom[4646] = 25'b1111111111010001001111110;
    rom[4647] = 25'b1111111111010000011111010;
    rom[4648] = 25'b1111111111001111101110111;
    rom[4649] = 25'b1111111111001110111110010;
    rom[4650] = 25'b1111111111001110001101101;
    rom[4651] = 25'b1111111111001101011101000;
    rom[4652] = 25'b1111111111001100101100001;
    rom[4653] = 25'b1111111111001011111011011;
    rom[4654] = 25'b1111111111001011001010101;
    rom[4655] = 25'b1111111111001010011001100;
    rom[4656] = 25'b1111111111001001101000101;
    rom[4657] = 25'b1111111111001000110111100;
    rom[4658] = 25'b1111111111001000000110100;
    rom[4659] = 25'b1111111111000111010101010;
    rom[4660] = 25'b1111111111000110100100010;
    rom[4661] = 25'b1111111111000101110011000;
    rom[4662] = 25'b1111111111000101000001101;
    rom[4663] = 25'b1111111111000100010000010;
    rom[4664] = 25'b1111111111000011011110111;
    rom[4665] = 25'b1111111111000010101101100;
    rom[4666] = 25'b1111111111000001111100000;
    rom[4667] = 25'b1111111111000001001010101;
    rom[4668] = 25'b1111111111000000011001000;
    rom[4669] = 25'b1111111110111111100111011;
    rom[4670] = 25'b1111111110111110110101110;
    rom[4671] = 25'b1111111110111110000100001;
    rom[4672] = 25'b1111111110111101010010011;
    rom[4673] = 25'b1111111110111100100000101;
    rom[4674] = 25'b1111111110111011101110111;
    rom[4675] = 25'b1111111110111010111101001;
    rom[4676] = 25'b1111111110111010001011011;
    rom[4677] = 25'b1111111110111001011001100;
    rom[4678] = 25'b1111111110111000100111110;
    rom[4679] = 25'b1111111110110111110101111;
    rom[4680] = 25'b1111111110110111000011111;
    rom[4681] = 25'b1111111110110110010010000;
    rom[4682] = 25'b1111111110110101100000000;
    rom[4683] = 25'b1111111110110100101110001;
    rom[4684] = 25'b1111111110110011111100001;
    rom[4685] = 25'b1111111110110011001010000;
    rom[4686] = 25'b1111111110110010011000001;
    rom[4687] = 25'b1111111110110001100110000;
    rom[4688] = 25'b1111111110110000110100000;
    rom[4689] = 25'b1111111110110000000010000;
    rom[4690] = 25'b1111111110101111001111111;
    rom[4691] = 25'b1111111110101110011101111;
    rom[4692] = 25'b1111111110101101101011111;
    rom[4693] = 25'b1111111110101100111001110;
    rom[4694] = 25'b1111111110101100000111110;
    rom[4695] = 25'b1111111110101011010101101;
    rom[4696] = 25'b1111111110101010100011100;
    rom[4697] = 25'b1111111110101001110001100;
    rom[4698] = 25'b1111111110101000111111100;
    rom[4699] = 25'b1111111110101000001101100;
    rom[4700] = 25'b1111111110100111011011011;
    rom[4701] = 25'b1111111110100110101001011;
    rom[4702] = 25'b1111111110100101110111011;
    rom[4703] = 25'b1111111110100101000101011;
    rom[4704] = 25'b1111111110100100010011011;
    rom[4705] = 25'b1111111110100011100001011;
    rom[4706] = 25'b1111111110100010101111100;
    rom[4707] = 25'b1111111110100001111101100;
    rom[4708] = 25'b1111111110100001001011100;
    rom[4709] = 25'b1111111110100000011001101;
    rom[4710] = 25'b1111111110011111100111110;
    rom[4711] = 25'b1111111110011110110110000;
    rom[4712] = 25'b1111111110011110000100001;
    rom[4713] = 25'b1111111110011101010010011;
    rom[4714] = 25'b1111111110011100100000101;
    rom[4715] = 25'b1111111110011011101110111;
    rom[4716] = 25'b1111111110011010111101001;
    rom[4717] = 25'b1111111110011010001011100;
    rom[4718] = 25'b1111111110011001011001111;
    rom[4719] = 25'b1111111110011000101000010;
    rom[4720] = 25'b1111111110010111110110110;
    rom[4721] = 25'b1111111110010111000101010;
    rom[4722] = 25'b1111111110010110010011111;
    rom[4723] = 25'b1111111110010101100010011;
    rom[4724] = 25'b1111111110010100110001000;
    rom[4725] = 25'b1111111110010011111111101;
    rom[4726] = 25'b1111111110010011001110011;
    rom[4727] = 25'b1111111110010010011101001;
    rom[4728] = 25'b1111111110010001101100000;
    rom[4729] = 25'b1111111110010000111011000;
    rom[4730] = 25'b1111111110010000001001111;
    rom[4731] = 25'b1111111110001111011000111;
    rom[4732] = 25'b1111111110001110100111111;
    rom[4733] = 25'b1111111110001101110111000;
    rom[4734] = 25'b1111111110001101000110010;
    rom[4735] = 25'b1111111110001100010101100;
    rom[4736] = 25'b1111111110001011100100111;
    rom[4737] = 25'b1111111110001010110100001;
    rom[4738] = 25'b1111111110001010000011101;
    rom[4739] = 25'b1111111110001001010011001;
    rom[4740] = 25'b1111111110001000100010110;
    rom[4741] = 25'b1111111110000111110010100;
    rom[4742] = 25'b1111111110000111000010001;
    rom[4743] = 25'b1111111110000110010010000;
    rom[4744] = 25'b1111111110000101100010000;
    rom[4745] = 25'b1111111110000100110010000;
    rom[4746] = 25'b1111111110000100000010001;
    rom[4747] = 25'b1111111110000011010010010;
    rom[4748] = 25'b1111111110000010100010100;
    rom[4749] = 25'b1111111110000001110010110;
    rom[4750] = 25'b1111111110000001000011010;
    rom[4751] = 25'b1111111110000000010011111;
    rom[4752] = 25'b1111111101111111100100011;
    rom[4753] = 25'b1111111101111110110101001;
    rom[4754] = 25'b1111111101111110000101111;
    rom[4755] = 25'b1111111101111101010110110;
    rom[4756] = 25'b1111111101111100100111110;
    rom[4757] = 25'b1111111101111011111001000;
    rom[4758] = 25'b1111111101111011001010010;
    rom[4759] = 25'b1111111101111010011011101;
    rom[4760] = 25'b1111111101111001101101000;
    rom[4761] = 25'b1111111101111000111110100;
    rom[4762] = 25'b1111111101111000010000010;
    rom[4763] = 25'b1111111101110111100010000;
    rom[4764] = 25'b1111111101110110110011111;
    rom[4765] = 25'b1111111101110110000101111;
    rom[4766] = 25'b1111111101110101011000000;
    rom[4767] = 25'b1111111101110100101010010;
    rom[4768] = 25'b1111111101110011111100101;
    rom[4769] = 25'b1111111101110011001111001;
    rom[4770] = 25'b1111111101110010100001110;
    rom[4771] = 25'b1111111101110001110100100;
    rom[4772] = 25'b1111111101110001000111011;
    rom[4773] = 25'b1111111101110000011010011;
    rom[4774] = 25'b1111111101101111101101100;
    rom[4775] = 25'b1111111101101111000000110;
    rom[4776] = 25'b1111111101101110010100010;
    rom[4777] = 25'b1111111101101101100111110;
    rom[4778] = 25'b1111111101101100111011100;
    rom[4779] = 25'b1111111101101100001111010;
    rom[4780] = 25'b1111111101101011100011010;
    rom[4781] = 25'b1111111101101010110111011;
    rom[4782] = 25'b1111111101101010001011101;
    rom[4783] = 25'b1111111101101001100000000;
    rom[4784] = 25'b1111111101101000110100101;
    rom[4785] = 25'b1111111101101000001001011;
    rom[4786] = 25'b1111111101100111011110010;
    rom[4787] = 25'b1111111101100110110011010;
    rom[4788] = 25'b1111111101100110001000100;
    rom[4789] = 25'b1111111101100101011101111;
    rom[4790] = 25'b1111111101100100110011011;
    rom[4791] = 25'b1111111101100100001001001;
    rom[4792] = 25'b1111111101100011011111000;
    rom[4793] = 25'b1111111101100010110101000;
    rom[4794] = 25'b1111111101100010001011001;
    rom[4795] = 25'b1111111101100001100001100;
    rom[4796] = 25'b1111111101100000111000001;
    rom[4797] = 25'b1111111101100000001110110;
    rom[4798] = 25'b1111111101011111100101101;
    rom[4799] = 25'b1111111101011110111100110;
    rom[4800] = 25'b1111111101011110010011111;
    rom[4801] = 25'b1111111101011101101011011;
    rom[4802] = 25'b1111111101011101000011000;
    rom[4803] = 25'b1111111101011100011010110;
    rom[4804] = 25'b1111111101011011110010110;
    rom[4805] = 25'b1111111101011011001010111;
    rom[4806] = 25'b1111111101011010100011010;
    rom[4807] = 25'b1111111101011001111011110;
    rom[4808] = 25'b1111111101011001010100101;
    rom[4809] = 25'b1111111101011000101101100;
    rom[4810] = 25'b1111111101011000000110101;
    rom[4811] = 25'b1111111101010111100000000;
    rom[4812] = 25'b1111111101010110111001100;
    rom[4813] = 25'b1111111101010110010011010;
    rom[4814] = 25'b1111111101010101101101010;
    rom[4815] = 25'b1111111101010101000111100;
    rom[4816] = 25'b1111111101010100100001111;
    rom[4817] = 25'b1111111101010011111100011;
    rom[4818] = 25'b1111111101010011010111010;
    rom[4819] = 25'b1111111101010010110010010;
    rom[4820] = 25'b1111111101010010001101100;
    rom[4821] = 25'b1111111101010001101000111;
    rom[4822] = 25'b1111111101010001000100100;
    rom[4823] = 25'b1111111101010000100000100;
    rom[4824] = 25'b1111111101001111111100100;
    rom[4825] = 25'b1111111101001111011000111;
    rom[4826] = 25'b1111111101001110110101011;
    rom[4827] = 25'b1111111101001110010010010;
    rom[4828] = 25'b1111111101001101101111010;
    rom[4829] = 25'b1111111101001101001100100;
    rom[4830] = 25'b1111111101001100101010000;
    rom[4831] = 25'b1111111101001100000111110;
    rom[4832] = 25'b1111111101001011100101101;
    rom[4833] = 25'b1111111101001011000011111;
    rom[4834] = 25'b1111111101001010100010011;
    rom[4835] = 25'b1111111101001010000001000;
    rom[4836] = 25'b1111111101001001100000000;
    rom[4837] = 25'b1111111101001000111111001;
    rom[4838] = 25'b1111111101001000011110100;
    rom[4839] = 25'b1111111101000111111110010;
    rom[4840] = 25'b1111111101000111011110001;
    rom[4841] = 25'b1111111101000110111110011;
    rom[4842] = 25'b1111111101000110011110110;
    rom[4843] = 25'b1111111101000101111111100;
    rom[4844] = 25'b1111111101000101100000100;
    rom[4845] = 25'b1111111101000101000001101;
    rom[4846] = 25'b1111111101000100100011001;
    rom[4847] = 25'b1111111101000100000101000;
    rom[4848] = 25'b1111111101000011100111000;
    rom[4849] = 25'b1111111101000011001001010;
    rom[4850] = 25'b1111111101000010101011110;
    rom[4851] = 25'b1111111101000010001110101;
    rom[4852] = 25'b1111111101000001110001110;
    rom[4853] = 25'b1111111101000001010101000;
    rom[4854] = 25'b1111111101000000111000110;
    rom[4855] = 25'b1111111101000000011100101;
    rom[4856] = 25'b1111111101000000000000110;
    rom[4857] = 25'b1111111100111111100101010;
    rom[4858] = 25'b1111111100111111001010000;
    rom[4859] = 25'b1111111100111110101111001;
    rom[4860] = 25'b1111111100111110010100100;
    rom[4861] = 25'b1111111100111101111010001;
    rom[4862] = 25'b1111111100111101100000000;
    rom[4863] = 25'b1111111100111101000110010;
    rom[4864] = 25'b1111111100111100101100110;
    rom[4865] = 25'b1111111100111100010011100;
    rom[4866] = 25'b1111111100111011111010101;
    rom[4867] = 25'b1111111100111011100010000;
    rom[4868] = 25'b1111111100111011001001110;
    rom[4869] = 25'b1111111100111010110001110;
    rom[4870] = 25'b1111111100111010011010000;
    rom[4871] = 25'b1111111100111010000010101;
    rom[4872] = 25'b1111111100111001101011100;
    rom[4873] = 25'b1111111100111001010100101;
    rom[4874] = 25'b1111111100111000111110010;
    rom[4875] = 25'b1111111100111000101000001;
    rom[4876] = 25'b1111111100111000010010010;
    rom[4877] = 25'b1111111100110111111100110;
    rom[4878] = 25'b1111111100110111100111100;
    rom[4879] = 25'b1111111100110111010010101;
    rom[4880] = 25'b1111111100110110111110000;
    rom[4881] = 25'b1111111100110110101001111;
    rom[4882] = 25'b1111111100110110010101111;
    rom[4883] = 25'b1111111100110110000010010;
    rom[4884] = 25'b1111111100110101101111000;
    rom[4885] = 25'b1111111100110101011100000;
    rom[4886] = 25'b1111111100110101001001011;
    rom[4887] = 25'b1111111100110100110111001;
    rom[4888] = 25'b1111111100110100100101001;
    rom[4889] = 25'b1111111100110100010011101;
    rom[4890] = 25'b1111111100110100000010010;
    rom[4891] = 25'b1111111100110011110001011;
    rom[4892] = 25'b1111111100110011100000110;
    rom[4893] = 25'b1111111100110011010000100;
    rom[4894] = 25'b1111111100110011000000101;
    rom[4895] = 25'b1111111100110010110001000;
    rom[4896] = 25'b1111111100110010100001110;
    rom[4897] = 25'b1111111100110010010010111;
    rom[4898] = 25'b1111111100110010000100010;
    rom[4899] = 25'b1111111100110001110110001;
    rom[4900] = 25'b1111111100110001101000011;
    rom[4901] = 25'b1111111100110001011010111;
    rom[4902] = 25'b1111111100110001001101101;
    rom[4903] = 25'b1111111100110001000000111;
    rom[4904] = 25'b1111111100110000110100100;
    rom[4905] = 25'b1111111100110000101000100;
    rom[4906] = 25'b1111111100110000011100110;
    rom[4907] = 25'b1111111100110000010001011;
    rom[4908] = 25'b1111111100110000000110011;
    rom[4909] = 25'b1111111100101111111011110;
    rom[4910] = 25'b1111111100101111110001101;
    rom[4911] = 25'b1111111100101111100111110;
    rom[4912] = 25'b1111111100101111011110010;
    rom[4913] = 25'b1111111100101111010101001;
    rom[4914] = 25'b1111111100101111001100010;
    rom[4915] = 25'b1111111100101111000011111;
    rom[4916] = 25'b1111111100101110111011111;
    rom[4917] = 25'b1111111100101110110100010;
    rom[4918] = 25'b1111111100101110101101000;
    rom[4919] = 25'b1111111100101110100110001;
    rom[4920] = 25'b1111111100101110011111101;
    rom[4921] = 25'b1111111100101110011001101;
    rom[4922] = 25'b1111111100101110010011111;
    rom[4923] = 25'b1111111100101110001110011;
    rom[4924] = 25'b1111111100101110001001011;
    rom[4925] = 25'b1111111100101110000100111;
    rom[4926] = 25'b1111111100101110000000101;
    rom[4927] = 25'b1111111100101101111100111;
    rom[4928] = 25'b1111111100101101111001100;
    rom[4929] = 25'b1111111100101101110110100;
    rom[4930] = 25'b1111111100101101110011111;
    rom[4931] = 25'b1111111100101101110001101;
    rom[4932] = 25'b1111111100101101101111110;
    rom[4933] = 25'b1111111100101101101110010;
    rom[4934] = 25'b1111111100101101101101010;
    rom[4935] = 25'b1111111100101101101100101;
    rom[4936] = 25'b1111111100101101101100011;
    rom[4937] = 25'b1111111100101101101100101;
    rom[4938] = 25'b1111111100101101101101001;
    rom[4939] = 25'b1111111100101101101110001;
    rom[4940] = 25'b1111111100101101101111100;
    rom[4941] = 25'b1111111100101101110001010;
    rom[4942] = 25'b1111111100101101110011100;
    rom[4943] = 25'b1111111100101101110110000;
    rom[4944] = 25'b1111111100101101111001001;
    rom[4945] = 25'b1111111100101101111100100;
    rom[4946] = 25'b1111111100101110000000011;
    rom[4947] = 25'b1111111100101110000100101;
    rom[4948] = 25'b1111111100101110001001010;
    rom[4949] = 25'b1111111100101110001110011;
    rom[4950] = 25'b1111111100101110010011111;
    rom[4951] = 25'b1111111100101110011001110;
    rom[4952] = 25'b1111111100101110100000001;
    rom[4953] = 25'b1111111100101110100110111;
    rom[4954] = 25'b1111111100101110101110001;
    rom[4955] = 25'b1111111100101110110101101;
    rom[4956] = 25'b1111111100101110111101110;
    rom[4957] = 25'b1111111100101111000110010;
    rom[4958] = 25'b1111111100101111001111000;
    rom[4959] = 25'b1111111100101111011000011;
    rom[4960] = 25'b1111111100101111100010001;
    rom[4961] = 25'b1111111100101111101100010;
    rom[4962] = 25'b1111111100101111110110111;
    rom[4963] = 25'b1111111100110000000001111;
    rom[4964] = 25'b1111111100110000001101011;
    rom[4965] = 25'b1111111100110000011001010;
    rom[4966] = 25'b1111111100110000100101101;
    rom[4967] = 25'b1111111100110000110010011;
    rom[4968] = 25'b1111111100110000111111100;
    rom[4969] = 25'b1111111100110001001101001;
    rom[4970] = 25'b1111111100110001011011010;
    rom[4971] = 25'b1111111100110001101001110;
    rom[4972] = 25'b1111111100110001111000110;
    rom[4973] = 25'b1111111100110010001000001;
    rom[4974] = 25'b1111111100110010011000000;
    rom[4975] = 25'b1111111100110010101000010;
    rom[4976] = 25'b1111111100110010111000111;
    rom[4977] = 25'b1111111100110011001010001;
    rom[4978] = 25'b1111111100110011011011110;
    rom[4979] = 25'b1111111100110011101101110;
    rom[4980] = 25'b1111111100110100000000010;
    rom[4981] = 25'b1111111100110100010011001;
    rom[4982] = 25'b1111111100110100100110101;
    rom[4983] = 25'b1111111100110100111010011;
    rom[4984] = 25'b1111111100110101001110110;
    rom[4985] = 25'b1111111100110101100011100;
    rom[4986] = 25'b1111111100110101111000110;
    rom[4987] = 25'b1111111100110110001110010;
    rom[4988] = 25'b1111111100110110100100011;
    rom[4989] = 25'b1111111100110110111011000;
    rom[4990] = 25'b1111111100110111010010000;
    rom[4991] = 25'b1111111100110111101001011;
    rom[4992] = 25'b1111111100111000000001011;
    rom[4993] = 25'b1111111100111000011001101;
    rom[4994] = 25'b1111111100111000110010100;
    rom[4995] = 25'b1111111100111001001011111;
    rom[4996] = 25'b1111111100111001100101101;
    rom[4997] = 25'b1111111100111001111111110;
    rom[4998] = 25'b1111111100111010011010011;
    rom[4999] = 25'b1111111100111010110101100;
    rom[5000] = 25'b1111111100111011010001001;
    rom[5001] = 25'b1111111100111011101101001;
    rom[5002] = 25'b1111111100111100001001101;
    rom[5003] = 25'b1111111100111100100110101;
    rom[5004] = 25'b1111111100111101000100001;
    rom[5005] = 25'b1111111100111101100010000;
    rom[5006] = 25'b1111111100111110000000010;
    rom[5007] = 25'b1111111100111110011111001;
    rom[5008] = 25'b1111111100111110111110011;
    rom[5009] = 25'b1111111100111111011110001;
    rom[5010] = 25'b1111111100111111111110011;
    rom[5011] = 25'b1111111101000000011111000;
    rom[5012] = 25'b1111111101000001000000001;
    rom[5013] = 25'b1111111101000001100001110;
    rom[5014] = 25'b1111111101000010000011110;
    rom[5015] = 25'b1111111101000010100110011;
    rom[5016] = 25'b1111111101000011001001010;
    rom[5017] = 25'b1111111101000011101100110;
    rom[5018] = 25'b1111111101000100010000110;
    rom[5019] = 25'b1111111101000100110101010;
    rom[5020] = 25'b1111111101000101011010000;
    rom[5021] = 25'b1111111101000101111111011;
    rom[5022] = 25'b1111111101000110100101001;
    rom[5023] = 25'b1111111101000111001011100;
    rom[5024] = 25'b1111111101000111110010010;
    rom[5025] = 25'b1111111101001000011001100;
    rom[5026] = 25'b1111111101001001000001001;
    rom[5027] = 25'b1111111101001001101001010;
    rom[5028] = 25'b1111111101001010010001111;
    rom[5029] = 25'b1111111101001010111011000;
    rom[5030] = 25'b1111111101001011100100101;
    rom[5031] = 25'b1111111101001100001110110;
    rom[5032] = 25'b1111111101001100111001010;
    rom[5033] = 25'b1111111101001101100100010;
    rom[5034] = 25'b1111111101001110001111101;
    rom[5035] = 25'b1111111101001110111011101;
    rom[5036] = 25'b1111111101001111101000000;
    rom[5037] = 25'b1111111101010000010100111;
    rom[5038] = 25'b1111111101010001000010001;
    rom[5039] = 25'b1111111101010001110000000;
    rom[5040] = 25'b1111111101010010011110011;
    rom[5041] = 25'b1111111101010011001101001;
    rom[5042] = 25'b1111111101010011111100011;
    rom[5043] = 25'b1111111101010100101100000;
    rom[5044] = 25'b1111111101010101011100010;
    rom[5045] = 25'b1111111101010110001100111;
    rom[5046] = 25'b1111111101010110111110000;
    rom[5047] = 25'b1111111101010111101111101;
    rom[5048] = 25'b1111111101011000100001101;
    rom[5049] = 25'b1111111101011001010100001;
    rom[5050] = 25'b1111111101011010000111001;
    rom[5051] = 25'b1111111101011010111010110;
    rom[5052] = 25'b1111111101011011101110101;
    rom[5053] = 25'b1111111101011100100011000;
    rom[5054] = 25'b1111111101011101011000000;
    rom[5055] = 25'b1111111101011110001101011;
    rom[5056] = 25'b1111111101011111000011001;
    rom[5057] = 25'b1111111101011111111001100;
    rom[5058] = 25'b1111111101100000110000010;
    rom[5059] = 25'b1111111101100001100111100;
    rom[5060] = 25'b1111111101100010011111010;
    rom[5061] = 25'b1111111101100011010111011;
    rom[5062] = 25'b1111111101100100010000000;
    rom[5063] = 25'b1111111101100101001001001;
    rom[5064] = 25'b1111111101100110000010110;
    rom[5065] = 25'b1111111101100110111100110;
    rom[5066] = 25'b1111111101100111110111011;
    rom[5067] = 25'b1111111101101000110010011;
    rom[5068] = 25'b1111111101101001101101110;
    rom[5069] = 25'b1111111101101010101001101;
    rom[5070] = 25'b1111111101101011100110000;
    rom[5071] = 25'b1111111101101100100010111;
    rom[5072] = 25'b1111111101101101100000010;
    rom[5073] = 25'b1111111101101110011110000;
    rom[5074] = 25'b1111111101101111011100010;
    rom[5075] = 25'b1111111101110000011011000;
    rom[5076] = 25'b1111111101110001011010001;
    rom[5077] = 25'b1111111101110010011001110;
    rom[5078] = 25'b1111111101110011011001111;
    rom[5079] = 25'b1111111101110100011010011;
    rom[5080] = 25'b1111111101110101011011100;
    rom[5081] = 25'b1111111101110110011101000;
    rom[5082] = 25'b1111111101110111011110111;
    rom[5083] = 25'b1111111101111000100001010;
    rom[5084] = 25'b1111111101111001100100001;
    rom[5085] = 25'b1111111101111010100111011;
    rom[5086] = 25'b1111111101111011101011010;
    rom[5087] = 25'b1111111101111100101111100;
    rom[5088] = 25'b1111111101111101110100001;
    rom[5089] = 25'b1111111101111110111001010;
    rom[5090] = 25'b1111111101111111111110110;
    rom[5091] = 25'b1111111110000001000100111;
    rom[5092] = 25'b1111111110000010001011011;
    rom[5093] = 25'b1111111110000011010010011;
    rom[5094] = 25'b1111111110000100011001101;
    rom[5095] = 25'b1111111110000101100001100;
    rom[5096] = 25'b1111111110000110101001111;
    rom[5097] = 25'b1111111110000111110010101;
    rom[5098] = 25'b1111111110001000111011110;
    rom[5099] = 25'b1111111110001010000101100;
    rom[5100] = 25'b1111111110001011001111101;
    rom[5101] = 25'b1111111110001100011010001;
    rom[5102] = 25'b1111111110001101100101000;
    rom[5103] = 25'b1111111110001110110000011;
    rom[5104] = 25'b1111111110001111111100011;
    rom[5105] = 25'b1111111110010001001000100;
    rom[5106] = 25'b1111111110010010010101010;
    rom[5107] = 25'b1111111110010011100010100;
    rom[5108] = 25'b1111111110010100110000001;
    rom[5109] = 25'b1111111110010101111110010;
    rom[5110] = 25'b1111111110010111001100110;
    rom[5111] = 25'b1111111110011000011011101;
    rom[5112] = 25'b1111111110011001101011000;
    rom[5113] = 25'b1111111110011010111010110;
    rom[5114] = 25'b1111111110011100001011000;
    rom[5115] = 25'b1111111110011101011011101;
    rom[5116] = 25'b1111111110011110101100110;
    rom[5117] = 25'b1111111110011111111110010;
    rom[5118] = 25'b1111111110100001010000010;
    rom[5119] = 25'b1111111110100010100010100;
    rom[5120] = 25'b1111111110100011110101010;
    rom[5121] = 25'b1111111110100101001000100;
    rom[5122] = 25'b1111111110100110011100001;
    rom[5123] = 25'b1111111110100111110000010;
    rom[5124] = 25'b1111111110101001000100110;
    rom[5125] = 25'b1111111110101010011001100;
    rom[5126] = 25'b1111111110101011101110111;
    rom[5127] = 25'b1111111110101101000100101;
    rom[5128] = 25'b1111111110101110011010110;
    rom[5129] = 25'b1111111110101111110001010;
    rom[5130] = 25'b1111111110110001001000010;
    rom[5131] = 25'b1111111110110010011111101;
    rom[5132] = 25'b1111111110110011110111011;
    rom[5133] = 25'b1111111110110101001111101;
    rom[5134] = 25'b1111111110110110101000001;
    rom[5135] = 25'b1111111110111000000001001;
    rom[5136] = 25'b1111111110111001011010100;
    rom[5137] = 25'b1111111110111010110100011;
    rom[5138] = 25'b1111111110111100001110100;
    rom[5139] = 25'b1111111110111101101001001;
    rom[5140] = 25'b1111111110111111000100001;
    rom[5141] = 25'b1111111111000000011111011;
    rom[5142] = 25'b1111111111000001111011010;
    rom[5143] = 25'b1111111111000011010111011;
    rom[5144] = 25'b1111111111000100110011111;
    rom[5145] = 25'b1111111111000110010001000;
    rom[5146] = 25'b1111111111000111101110001;
    rom[5147] = 25'b1111111111001001001100000;
    rom[5148] = 25'b1111111111001010101010000;
    rom[5149] = 25'b1111111111001100001000100;
    rom[5150] = 25'b1111111111001101100111011;
    rom[5151] = 25'b1111111111001111000110101;
    rom[5152] = 25'b1111111111010000100110010;
    rom[5153] = 25'b1111111111010010000110010;
    rom[5154] = 25'b1111111111010011100110100;
    rom[5155] = 25'b1111111111010101000111010;
    rom[5156] = 25'b1111111111010110101000100;
    rom[5157] = 25'b1111111111011000001001111;
    rom[5158] = 25'b1111111111011001101011110;
    rom[5159] = 25'b1111111111011011001101111;
    rom[5160] = 25'b1111111111011100110000011;
    rom[5161] = 25'b1111111111011110010011011;
    rom[5162] = 25'b1111111111011111110110101;
    rom[5163] = 25'b1111111111100001011010010;
    rom[5164] = 25'b1111111111100010111110010;
    rom[5165] = 25'b1111111111100100100010101;
    rom[5166] = 25'b1111111111100110000111010;
    rom[5167] = 25'b1111111111100111101100010;
    rom[5168] = 25'b1111111111101001010001110;
    rom[5169] = 25'b1111111111101010110111011;
    rom[5170] = 25'b1111111111101100011101011;
    rom[5171] = 25'b1111111111101110000011111;
    rom[5172] = 25'b1111111111101111101010101;
    rom[5173] = 25'b1111111111110001010001101;
    rom[5174] = 25'b1111111111110010111001000;
    rom[5175] = 25'b1111111111110100100000110;
    rom[5176] = 25'b1111111111110110001000111;
    rom[5177] = 25'b1111111111110111110001010;
    rom[5178] = 25'b1111111111111001011010000;
    rom[5179] = 25'b1111111111111011000011000;
    rom[5180] = 25'b1111111111111100101100011;
    rom[5181] = 25'b1111111111111110010110000;
    rom[5182] = 25'b0000000000000000000000000;
    rom[5183] = 25'b0000000000000001101010001;
    rom[5184] = 25'b0000000000000011010100110;
    rom[5185] = 25'b0000000000000100111111110;
    rom[5186] = 25'b0000000000000110101011000;
    rom[5187] = 25'b0000000000001000010110100;
    rom[5188] = 25'b0000000000001010000010010;
    rom[5189] = 25'b0000000000001011101110100;
    rom[5190] = 25'b0000000000001101011010111;
    rom[5191] = 25'b0000000000001111000111101;
    rom[5192] = 25'b0000000000010000110100101;
    rom[5193] = 25'b0000000000010010100010000;
    rom[5194] = 25'b0000000000010100001111101;
    rom[5195] = 25'b0000000000010101111101011;
    rom[5196] = 25'b0000000000010111101011100;
    rom[5197] = 25'b0000000000011001011010000;
    rom[5198] = 25'b0000000000011011001000101;
    rom[5199] = 25'b0000000000011100110111101;
    rom[5200] = 25'b0000000000011110100111000;
    rom[5201] = 25'b0000000000100000010110100;
    rom[5202] = 25'b0000000000100010000110011;
    rom[5203] = 25'b0000000000100011110110011;
    rom[5204] = 25'b0000000000100101100110101;
    rom[5205] = 25'b0000000000100111010111010;
    rom[5206] = 25'b0000000000101001001000001;
    rom[5207] = 25'b0000000000101010111001001;
    rom[5208] = 25'b0000000000101100101010101;
    rom[5209] = 25'b0000000000101110011100001;
    rom[5210] = 25'b0000000000110000001110000;
    rom[5211] = 25'b0000000000110010000000000;
    rom[5212] = 25'b0000000000110011110010011;
    rom[5213] = 25'b0000000000110101100100111;
    rom[5214] = 25'b0000000000110111010111110;
    rom[5215] = 25'b0000000000111001001010110;
    rom[5216] = 25'b0000000000111010111110000;
    rom[5217] = 25'b0000000000111100110001100;
    rom[5218] = 25'b0000000000111110100101001;
    rom[5219] = 25'b0000000001000000011001001;
    rom[5220] = 25'b0000000001000010001101010;
    rom[5221] = 25'b0000000001000100000001101;
    rom[5222] = 25'b0000000001000101110110001;
    rom[5223] = 25'b0000000001000111101011000;
    rom[5224] = 25'b0000000001001001011111111;
    rom[5225] = 25'b0000000001001011010101001;
    rom[5226] = 25'b0000000001001101001010100;
    rom[5227] = 25'b0000000001001111000000000;
    rom[5228] = 25'b0000000001010000110101111;
    rom[5229] = 25'b0000000001010010101011111;
    rom[5230] = 25'b0000000001010100100010000;
    rom[5231] = 25'b0000000001010110011000011;
    rom[5232] = 25'b0000000001011000001110111;
    rom[5233] = 25'b0000000001011010000101101;
    rom[5234] = 25'b0000000001011011111100011;
    rom[5235] = 25'b0000000001011101110011100;
    rom[5236] = 25'b0000000001011111101010110;
    rom[5237] = 25'b0000000001100001100010001;
    rom[5238] = 25'b0000000001100011011001101;
    rom[5239] = 25'b0000000001100101010001011;
    rom[5240] = 25'b0000000001100111001001010;
    rom[5241] = 25'b0000000001101001000001011;
    rom[5242] = 25'b0000000001101010111001100;
    rom[5243] = 25'b0000000001101100110001110;
    rom[5244] = 25'b0000000001101110101010011;
    rom[5245] = 25'b0000000001110000100010111;
    rom[5246] = 25'b0000000001110010011011101;
    rom[5247] = 25'b0000000001110100010100100;
    rom[5248] = 25'b0000000001110110001101100;
    rom[5249] = 25'b0000000001111000000110110;
    rom[5250] = 25'b0000000001111010000000000;
    rom[5251] = 25'b0000000001111011111001100;
    rom[5252] = 25'b0000000001111101110011000;
    rom[5253] = 25'b0000000001111111101100101;
    rom[5254] = 25'b0000000010000001100110011;
    rom[5255] = 25'b0000000010000011100000001;
    rom[5256] = 25'b0000000010000101011010001;
    rom[5257] = 25'b0000000010000111010100010;
    rom[5258] = 25'b0000000010001001001110011;
    rom[5259] = 25'b0000000010001011001000101;
    rom[5260] = 25'b0000000010001101000011000;
    rom[5261] = 25'b0000000010001110111101011;
    rom[5262] = 25'b0000000010010000111000000;
    rom[5263] = 25'b0000000010010010110010100;
    rom[5264] = 25'b0000000010010100101101010;
    rom[5265] = 25'b0000000010010110101000000;
    rom[5266] = 25'b0000000010011000100010110;
    rom[5267] = 25'b0000000010011010011101110;
    rom[5268] = 25'b0000000010011100011000110;
    rom[5269] = 25'b0000000010011110010011110;
    rom[5270] = 25'b0000000010100000001110111;
    rom[5271] = 25'b0000000010100010001001111;
    rom[5272] = 25'b0000000010100100000101000;
    rom[5273] = 25'b0000000010100110000000011;
    rom[5274] = 25'b0000000010100111111011101;
    rom[5275] = 25'b0000000010101001110110111;
    rom[5276] = 25'b0000000010101011110010010;
    rom[5277] = 25'b0000000010101101101101101;
    rom[5278] = 25'b0000000010101111101001001;
    rom[5279] = 25'b0000000010110001100100100;
    rom[5280] = 25'b0000000010110011011111111;
    rom[5281] = 25'b0000000010110101011011011;
    rom[5282] = 25'b0000000010110111010110111;
    rom[5283] = 25'b0000000010111001010010011;
    rom[5284] = 25'b0000000010111011001101111;
    rom[5285] = 25'b0000000010111101001001011;
    rom[5286] = 25'b0000000010111111000100111;
    rom[5287] = 25'b0000000011000001000000100;
    rom[5288] = 25'b0000000011000010111011111;
    rom[5289] = 25'b0000000011000100110111011;
    rom[5290] = 25'b0000000011000110110010111;
    rom[5291] = 25'b0000000011001000101110010;
    rom[5292] = 25'b0000000011001010101001110;
    rom[5293] = 25'b0000000011001100100101001;
    rom[5294] = 25'b0000000011001110100000100;
    rom[5295] = 25'b0000000011010000011011111;
    rom[5296] = 25'b0000000011010010010111001;
    rom[5297] = 25'b0000000011010100010010011;
    rom[5298] = 25'b0000000011010110001101101;
    rom[5299] = 25'b0000000011011000001000110;
    rom[5300] = 25'b0000000011011010000011111;
    rom[5301] = 25'b0000000011011011111110111;
    rom[5302] = 25'b0000000011011101111001111;
    rom[5303] = 25'b0000000011011111110100110;
    rom[5304] = 25'b0000000011100001101111101;
    rom[5305] = 25'b0000000011100011101010100;
    rom[5306] = 25'b0000000011100101100101001;
    rom[5307] = 25'b0000000011100111011111111;
    rom[5308] = 25'b0000000011101001011010010;
    rom[5309] = 25'b0000000011101011010100110;
    rom[5310] = 25'b0000000011101101001111001;
    rom[5311] = 25'b0000000011101111001001011;
    rom[5312] = 25'b0000000011110001000011100;
    rom[5313] = 25'b0000000011110010111101101;
    rom[5314] = 25'b0000000011110100110111100;
    rom[5315] = 25'b0000000011110110110001011;
    rom[5316] = 25'b0000000011111000101011001;
    rom[5317] = 25'b0000000011111010100100110;
    rom[5318] = 25'b0000000011111100011110001;
    rom[5319] = 25'b0000000011111110010111100;
    rom[5320] = 25'b0000000100000000010000110;
    rom[5321] = 25'b0000000100000010001001111;
    rom[5322] = 25'b0000000100000100000010110;
    rom[5323] = 25'b0000000100000101111011100;
    rom[5324] = 25'b0000000100000111110100001;
    rom[5325] = 25'b0000000100001001101100110;
    rom[5326] = 25'b0000000100001011100100111;
    rom[5327] = 25'b0000000100001101011101001;
    rom[5328] = 25'b0000000100001111010101010;
    rom[5329] = 25'b0000000100010001001101000;
    rom[5330] = 25'b0000000100010011000100101;
    rom[5331] = 25'b0000000100010100111100001;
    rom[5332] = 25'b0000000100010110110011100;
    rom[5333] = 25'b0000000100011000101010101;
    rom[5334] = 25'b0000000100011010100001100;
    rom[5335] = 25'b0000000100011100011000010;
    rom[5336] = 25'b0000000100011110001110111;
    rom[5337] = 25'b0000000100100000000101001;
    rom[5338] = 25'b0000000100100001111011010;
    rom[5339] = 25'b0000000100100011110001010;
    rom[5340] = 25'b0000000100100101100111000;
    rom[5341] = 25'b0000000100100111011100011;
    rom[5342] = 25'b0000000100101001010001101;
    rom[5343] = 25'b0000000100101011000110110;
    rom[5344] = 25'b0000000100101100111011101;
    rom[5345] = 25'b0000000100101110110000001;
    rom[5346] = 25'b0000000100110000100100100;
    rom[5347] = 25'b0000000100110010011000101;
    rom[5348] = 25'b0000000100110100001100100;
    rom[5349] = 25'b0000000100110110000000000;
    rom[5350] = 25'b0000000100110111110011011;
    rom[5351] = 25'b0000000100111001100110011;
    rom[5352] = 25'b0000000100111011011001010;
    rom[5353] = 25'b0000000100111101001011111;
    rom[5354] = 25'b0000000100111110111110001;
    rom[5355] = 25'b0000000101000000110000001;
    rom[5356] = 25'b0000000101000010100001111;
    rom[5357] = 25'b0000000101000100010011010;
    rom[5358] = 25'b0000000101000110000100011;
    rom[5359] = 25'b0000000101000111110101010;
    rom[5360] = 25'b0000000101001001100101111;
    rom[5361] = 25'b0000000101001011010110001;
    rom[5362] = 25'b0000000101001101000110001;
    rom[5363] = 25'b0000000101001110110101110;
    rom[5364] = 25'b0000000101010000100101000;
    rom[5365] = 25'b0000000101010010010100000;
    rom[5366] = 25'b0000000101010100000010110;
    rom[5367] = 25'b0000000101010101110001000;
    rom[5368] = 25'b0000000101010111011111001;
    rom[5369] = 25'b0000000101011001001100110;
    rom[5370] = 25'b0000000101011010111010010;
    rom[5371] = 25'b0000000101011100100111001;
    rom[5372] = 25'b0000000101011110010011110;
    rom[5373] = 25'b0000000101100000000000001;
    rom[5374] = 25'b0000000101100001101100000;
    rom[5375] = 25'b0000000101100011010111101;
    rom[5376] = 25'b0000000101100101000010111;
    rom[5377] = 25'b0000000101100110101101110;
    rom[5378] = 25'b0000000101101000011000001;
    rom[5379] = 25'b0000000101101010000010010;
    rom[5380] = 25'b0000000101101011101100000;
    rom[5381] = 25'b0000000101101101010101011;
    rom[5382] = 25'b0000000101101110111110011;
    rom[5383] = 25'b0000000101110000100110111;
    rom[5384] = 25'b0000000101110010001111000;
    rom[5385] = 25'b0000000101110011110110101;
    rom[5386] = 25'b0000000101110101011110000;
    rom[5387] = 25'b0000000101110111000101000;
    rom[5388] = 25'b0000000101111000101011100;
    rom[5389] = 25'b0000000101111010010001101;
    rom[5390] = 25'b0000000101111011110111010;
    rom[5391] = 25'b0000000101111101011100100;
    rom[5392] = 25'b0000000101111111000001011;
    rom[5393] = 25'b0000000110000000100101101;
    rom[5394] = 25'b0000000110000010001001101;
    rom[5395] = 25'b0000000110000011101101000;
    rom[5396] = 25'b0000000110000101010000001;
    rom[5397] = 25'b0000000110000110110010101;
    rom[5398] = 25'b0000000110001000010100110;
    rom[5399] = 25'b0000000110001001110110011;
    rom[5400] = 25'b0000000110001011010111100;
    rom[5401] = 25'b0000000110001100111000010;
    rom[5402] = 25'b0000000110001110011000100;
    rom[5403] = 25'b0000000110001111111000010;
    rom[5404] = 25'b0000000110010001010111100;
    rom[5405] = 25'b0000000110010010110110010;
    rom[5406] = 25'b0000000110010100010100100;
    rom[5407] = 25'b0000000110010101110010011;
    rom[5408] = 25'b0000000110010111001111101;
    rom[5409] = 25'b0000000110011000101100100;
    rom[5410] = 25'b0000000110011010001000110;
    rom[5411] = 25'b0000000110011011100100100;
    rom[5412] = 25'b0000000110011100111111110;
    rom[5413] = 25'b0000000110011110011010100;
    rom[5414] = 25'b0000000110011111110100101;
    rom[5415] = 25'b0000000110100001001110011;
    rom[5416] = 25'b0000000110100010100111100;
    rom[5417] = 25'b0000000110100100000000000;
    rom[5418] = 25'b0000000110100101011000001;
    rom[5419] = 25'b0000000110100110101111101;
    rom[5420] = 25'b0000000110101000000110100;
    rom[5421] = 25'b0000000110101001011101000;
    rom[5422] = 25'b0000000110101010110010111;
    rom[5423] = 25'b0000000110101100001000001;
    rom[5424] = 25'b0000000110101101011100110;
    rom[5425] = 25'b0000000110101110110001000;
    rom[5426] = 25'b0000000110110000000100100;
    rom[5427] = 25'b0000000110110001010111011;
    rom[5428] = 25'b0000000110110010101001111;
    rom[5429] = 25'b0000000110110011111011101;
    rom[5430] = 25'b0000000110110101001100111;
    rom[5431] = 25'b0000000110110110011101100;
    rom[5432] = 25'b0000000110110111101101100;
    rom[5433] = 25'b0000000110111000111101000;
    rom[5434] = 25'b0000000110111010001011110;
    rom[5435] = 25'b0000000110111011011010000;
    rom[5436] = 25'b0000000110111100100111100;
    rom[5437] = 25'b0000000110111101110100100;
    rom[5438] = 25'b0000000110111111000000110;
    rom[5439] = 25'b0000000111000000001100100;
    rom[5440] = 25'b0000000111000001010111100;
    rom[5441] = 25'b0000000111000010100010000;
    rom[5442] = 25'b0000000111000011101011111;
    rom[5443] = 25'b0000000111000100110101000;
    rom[5444] = 25'b0000000111000101111101100;
    rom[5445] = 25'b0000000111000111000101010;
    rom[5446] = 25'b0000000111001000001100100;
    rom[5447] = 25'b0000000111001001010011000;
    rom[5448] = 25'b0000000111001010011000110;
    rom[5449] = 25'b0000000111001011011110000;
    rom[5450] = 25'b0000000111001100100010101;
    rom[5451] = 25'b0000000111001101100110011;
    rom[5452] = 25'b0000000111001110101001101;
    rom[5453] = 25'b0000000111001111101100000;
    rom[5454] = 25'b0000000111010000101101111;
    rom[5455] = 25'b0000000111010001101110111;
    rom[5456] = 25'b0000000111010010101111011;
    rom[5457] = 25'b0000000111010011101111000;
    rom[5458] = 25'b0000000111010100101110001;
    rom[5459] = 25'b0000000111010101101100011;
    rom[5460] = 25'b0000000111010110101001111;
    rom[5461] = 25'b0000000111010111100110111;
    rom[5462] = 25'b0000000111011000100010111;
    rom[5463] = 25'b0000000111011001011110011;
    rom[5464] = 25'b0000000111011010011001000;
    rom[5465] = 25'b0000000111011011010011001;
    rom[5466] = 25'b0000000111011100001100010;
    rom[5467] = 25'b0000000111011101000100110;
    rom[5468] = 25'b0000000111011101111100100;
    rom[5469] = 25'b0000000111011110110011100;
    rom[5470] = 25'b0000000111011111101001111;
    rom[5471] = 25'b0000000111100000011111010;
    rom[5472] = 25'b0000000111100001010100000;
    rom[5473] = 25'b0000000111100010001000000;
    rom[5474] = 25'b0000000111100010111011010;
    rom[5475] = 25'b0000000111100011101101110;
    rom[5476] = 25'b0000000111100100011111011;
    rom[5477] = 25'b0000000111100101010000010;
    rom[5478] = 25'b0000000111100110000000100;
    rom[5479] = 25'b0000000111100110101111110;
    rom[5480] = 25'b0000000111100111011110011;
    rom[5481] = 25'b0000000111101000001100001;
    rom[5482] = 25'b0000000111101000111001001;
    rom[5483] = 25'b0000000111101001100101011;
    rom[5484] = 25'b0000000111101010010000110;
    rom[5485] = 25'b0000000111101010111011010;
    rom[5486] = 25'b0000000111101011100101000;
    rom[5487] = 25'b0000000111101100001110001;
    rom[5488] = 25'b0000000111101100110110001;
    rom[5489] = 25'b0000000111101101011101100;
    rom[5490] = 25'b0000000111101110000100001;
    rom[5491] = 25'b0000000111101110101001110;
    rom[5492] = 25'b0000000111101111001110101;
    rom[5493] = 25'b0000000111101111110010101;
    rom[5494] = 25'b0000000111110000010101111;
    rom[5495] = 25'b0000000111110000111000001;
    rom[5496] = 25'b0000000111110001011001101;
    rom[5497] = 25'b0000000111110001111010011;
    rom[5498] = 25'b0000000111110010011010010;
    rom[5499] = 25'b0000000111110010111001010;
    rom[5500] = 25'b0000000111110011010111011;
    rom[5501] = 25'b0000000111110011110100100;
    rom[5502] = 25'b0000000111110100010001000;
    rom[5503] = 25'b0000000111110100101100100;
    rom[5504] = 25'b0000000111110101000111001;
    rom[5505] = 25'b0000000111110101100001000;
    rom[5506] = 25'b0000000111110101111010000;
    rom[5507] = 25'b0000000111110110010010000;
    rom[5508] = 25'b0000000111110110101001001;
    rom[5509] = 25'b0000000111110110111111100;
    rom[5510] = 25'b0000000111110111010100111;
    rom[5511] = 25'b0000000111110111101001011;
    rom[5512] = 25'b0000000111110111111101000;
    rom[5513] = 25'b0000000111111000001111110;
    rom[5514] = 25'b0000000111111000100001100;
    rom[5515] = 25'b0000000111111000110010100;
    rom[5516] = 25'b0000000111111001000010100;
    rom[5517] = 25'b0000000111111001010001101;
    rom[5518] = 25'b0000000111111001011111111;
    rom[5519] = 25'b0000000111111001101101001;
    rom[5520] = 25'b0000000111111001111001100;
    rom[5521] = 25'b0000000111111010000101000;
    rom[5522] = 25'b0000000111111010001111100;
    rom[5523] = 25'b0000000111111010011001001;
    rom[5524] = 25'b0000000111111010100001111;
    rom[5525] = 25'b0000000111111010101001101;
    rom[5526] = 25'b0000000111111010110000011;
    rom[5527] = 25'b0000000111111010110110011;
    rom[5528] = 25'b0000000111111010111011010;
    rom[5529] = 25'b0000000111111010111111010;
    rom[5530] = 25'b0000000111111011000010011;
    rom[5531] = 25'b0000000111111011000100100;
    rom[5532] = 25'b0000000111111011000101101;
    rom[5533] = 25'b0000000111111011000101111;
    rom[5534] = 25'b0000000111111011000101001;
    rom[5535] = 25'b0000000111111011000011011;
    rom[5536] = 25'b0000000111111011000000110;
    rom[5537] = 25'b0000000111111010111101001;
    rom[5538] = 25'b0000000111111010111000101;
    rom[5539] = 25'b0000000111111010110011000;
    rom[5540] = 25'b0000000111111010101100100;
    rom[5541] = 25'b0000000111111010100101000;
    rom[5542] = 25'b0000000111111010011100100;
    rom[5543] = 25'b0000000111111010010011001;
    rom[5544] = 25'b0000000111111010001000101;
    rom[5545] = 25'b0000000111111001111101010;
    rom[5546] = 25'b0000000111111001110000111;
    rom[5547] = 25'b0000000111111001100011100;
    rom[5548] = 25'b0000000111111001010101001;
    rom[5549] = 25'b0000000111111001000101110;
    rom[5550] = 25'b0000000111111000110101011;
    rom[5551] = 25'b0000000111111000100100001;
    rom[5552] = 25'b0000000111111000010001110;
    rom[5553] = 25'b0000000111110111111110100;
    rom[5554] = 25'b0000000111110111101010000;
    rom[5555] = 25'b0000000111110111010100101;
    rom[5556] = 25'b0000000111110110111110011;
    rom[5557] = 25'b0000000111110110100111000;
    rom[5558] = 25'b0000000111110110001110101;
    rom[5559] = 25'b0000000111110101110101010;
    rom[5560] = 25'b0000000111110101011010111;
    rom[5561] = 25'b0000000111110100111111011;
    rom[5562] = 25'b0000000111110100100010111;
    rom[5563] = 25'b0000000111110100000101100;
    rom[5564] = 25'b0000000111110011100111000;
    rom[5565] = 25'b0000000111110011000111100;
    rom[5566] = 25'b0000000111110010100111000;
    rom[5567] = 25'b0000000111110010000101100;
    rom[5568] = 25'b0000000111110001100010110;
    rom[5569] = 25'b0000000111110000111111001;
    rom[5570] = 25'b0000000111110000011010100;
    rom[5571] = 25'b0000000111101111110100111;
    rom[5572] = 25'b0000000111101111001110001;
    rom[5573] = 25'b0000000111101110100110010;
    rom[5574] = 25'b0000000111101101111101101;
    rom[5575] = 25'b0000000111101101010011110;
    rom[5576] = 25'b0000000111101100101000111;
    rom[5577] = 25'b0000000111101011111100111;
    rom[5578] = 25'b0000000111101011001111111;
    rom[5579] = 25'b0000000111101010100001111;
    rom[5580] = 25'b0000000111101001110010110;
    rom[5581] = 25'b0000000111101001000010110;
    rom[5582] = 25'b0000000111101000010001100;
    rom[5583] = 25'b0000000111100111011111001;
    rom[5584] = 25'b0000000111100110101100000;
    rom[5585] = 25'b0000000111100101110111100;
    rom[5586] = 25'b0000000111100101000010001;
    rom[5587] = 25'b0000000111100100001011110;
    rom[5588] = 25'b0000000111100011010100001;
    rom[5589] = 25'b0000000111100010011011101;
    rom[5590] = 25'b0000000111100001100010000;
    rom[5591] = 25'b0000000111100000100111001;
    rom[5592] = 25'b0000000111011111101011011;
    rom[5593] = 25'b0000000111011110101110101;
    rom[5594] = 25'b0000000111011101110000101;
    rom[5595] = 25'b0000000111011100110001101;
    rom[5596] = 25'b0000000111011011110001101;
    rom[5597] = 25'b0000000111011010110000100;
    rom[5598] = 25'b0000000111011001101110010;
    rom[5599] = 25'b0000000111011000101011000;
    rom[5600] = 25'b0000000111010111100110101;
    rom[5601] = 25'b0000000111010110100001010;
    rom[5602] = 25'b0000000111010101011010110;
    rom[5603] = 25'b0000000111010100010011001;
    rom[5604] = 25'b0000000111010011001010100;
    rom[5605] = 25'b0000000111010010000000110;
    rom[5606] = 25'b0000000111010000110110000;
    rom[5607] = 25'b0000000111001111101010001;
    rom[5608] = 25'b0000000111001110011101001;
    rom[5609] = 25'b0000000111001101001111001;
    rom[5610] = 25'b0000000111001100000000000;
    rom[5611] = 25'b0000000111001010101111111;
    rom[5612] = 25'b0000000111001001011110100;
    rom[5613] = 25'b0000000111001000001100001;
    rom[5614] = 25'b0000000111000110111000110;
    rom[5615] = 25'b0000000111000101100100001;
    rom[5616] = 25'b0000000111000100001110101;
    rom[5617] = 25'b0000000111000010110111111;
    rom[5618] = 25'b0000000111000001100000001;
    rom[5619] = 25'b0000000111000000000111010;
    rom[5620] = 25'b0000000110111110101101010;
    rom[5621] = 25'b0000000110111101010010010;
    rom[5622] = 25'b0000000110111011110110000;
    rom[5623] = 25'b0000000110111010011000111;
    rom[5624] = 25'b0000000110111000111010101;
    rom[5625] = 25'b0000000110110111011011001;
    rom[5626] = 25'b0000000110110101111010110;
    rom[5627] = 25'b0000000110110100011001001;
    rom[5628] = 25'b0000000110110010110110101;
    rom[5629] = 25'b0000000110110001010010110;
    rom[5630] = 25'b0000000110101111101110000;
    rom[5631] = 25'b0000000110101110001000001;
    rom[5632] = 25'b0000000110101100100001001;
    rom[5633] = 25'b0000000110101010111001000;
    rom[5634] = 25'b0000000110101001001111111;
    rom[5635] = 25'b0000000110100111100101101;
    rom[5636] = 25'b0000000110100101111010010;
    rom[5637] = 25'b0000000110100100001101111;
    rom[5638] = 25'b0000000110100010100000011;
    rom[5639] = 25'b0000000110100000110001110;
    rom[5640] = 25'b0000000110011111000010000;
    rom[5641] = 25'b0000000110011101010001011;
    rom[5642] = 25'b0000000110011011011111100;
    rom[5643] = 25'b0000000110011001101100101;
    rom[5644] = 25'b0000000110010111111000101;
    rom[5645] = 25'b0000000110010110000011100;
    rom[5646] = 25'b0000000110010100001101011;
    rom[5647] = 25'b0000000110010010010110000;
    rom[5648] = 25'b0000000110010000011101110;
    rom[5649] = 25'b0000000110001110100100010;
    rom[5650] = 25'b0000000110001100101001111;
    rom[5651] = 25'b0000000110001010101110010;
    rom[5652] = 25'b0000000110001000110001101;
    rom[5653] = 25'b0000000110000110110011111;
    rom[5654] = 25'b0000000110000100110101001;
    rom[5655] = 25'b0000000110000010110101010;
    rom[5656] = 25'b0000000110000000110100010;
    rom[5657] = 25'b0000000101111110110010010;
    rom[5658] = 25'b0000000101111100101111001;
    rom[5659] = 25'b0000000101111010101011000;
    rom[5660] = 25'b0000000101111000100101110;
    rom[5661] = 25'b0000000101110110011111100;
    rom[5662] = 25'b0000000101110100011000001;
    rom[5663] = 25'b0000000101110010001111101;
    rom[5664] = 25'b0000000101110000000110010;
    rom[5665] = 25'b0000000101101101111011101;
    rom[5666] = 25'b0000000101101011110000000;
    rom[5667] = 25'b0000000101101001100011011;
    rom[5668] = 25'b0000000101100111010101100;
    rom[5669] = 25'b0000000101100101000110110;
    rom[5670] = 25'b0000000101100010110110111;
    rom[5671] = 25'b0000000101100000100110000;
    rom[5672] = 25'b0000000101011110010011111;
    rom[5673] = 25'b0000000101011100000000111;
    rom[5674] = 25'b0000000101011001101100111;
    rom[5675] = 25'b0000000101010111010111110;
    rom[5676] = 25'b0000000101010101000001100;
    rom[5677] = 25'b0000000101010010101010011;
    rom[5678] = 25'b0000000101010000010010000;
    rom[5679] = 25'b0000000101001101111000110;
    rom[5680] = 25'b0000000101001011011110011;
    rom[5681] = 25'b0000000101001001000011000;
    rom[5682] = 25'b0000000101000110100110100;
    rom[5683] = 25'b0000000101000100001001001;
    rom[5684] = 25'b0000000101000001101010101;
    rom[5685] = 25'b0000000100111111001011000;
    rom[5686] = 25'b0000000100111100101010100;
    rom[5687] = 25'b0000000100111010001000111;
    rom[5688] = 25'b0000000100110111100110010;
    rom[5689] = 25'b0000000100110101000010101;
    rom[5690] = 25'b0000000100110010011101111;
    rom[5691] = 25'b0000000100101111111000010;
    rom[5692] = 25'b0000000100101101010001101;
    rom[5693] = 25'b0000000100101010101001111;
    rom[5694] = 25'b0000000100101000000001001;
    rom[5695] = 25'b0000000100100101010111011;
    rom[5696] = 25'b0000000100100010101100101;
    rom[5697] = 25'b0000000100100000000000110;
    rom[5698] = 25'b0000000100011101010100000;
    rom[5699] = 25'b0000000100011010100110010;
    rom[5700] = 25'b0000000100010111110111100;
    rom[5701] = 25'b0000000100010101000111110;
    rom[5702] = 25'b0000000100010010010111000;
    rom[5703] = 25'b0000000100001111100101010;
    rom[5704] = 25'b0000000100001100110010100;
    rom[5705] = 25'b0000000100001001111110110;
    rom[5706] = 25'b0000000100000111001010000;
    rom[5707] = 25'b0000000100000100010100011;
    rom[5708] = 25'b0000000100000001011101110;
    rom[5709] = 25'b0000000011111110100110001;
    rom[5710] = 25'b0000000011111011101101011;
    rom[5711] = 25'b0000000011111000110011111;
    rom[5712] = 25'b0000000011110101111001011;
    rom[5713] = 25'b0000000011110010111101110;
    rom[5714] = 25'b0000000011110000000001011;
    rom[5715] = 25'b0000000011101101000100000;
    rom[5716] = 25'b0000000011101010000101101;
    rom[5717] = 25'b0000000011100111000110010;
    rom[5718] = 25'b0000000011100100000101111;
    rom[5719] = 25'b0000000011100001000100110;
    rom[5720] = 25'b0000000011011110000010100;
    rom[5721] = 25'b0000000011011010111111011;
    rom[5722] = 25'b0000000011010111111011011;
    rom[5723] = 25'b0000000011010100110110011;
    rom[5724] = 25'b0000000011010001110000100;
    rom[5725] = 25'b0000000011001110101001110;
    rom[5726] = 25'b0000000011001011100010000;
    rom[5727] = 25'b0000000011001000011001010;
    rom[5728] = 25'b0000000011000101001111101;
    rom[5729] = 25'b0000000011000010000101001;
    rom[5730] = 25'b0000000010111110111001110;
    rom[5731] = 25'b0000000010111011101101011;
    rom[5732] = 25'b0000000010111000100000010;
    rom[5733] = 25'b0000000010110101010010001;
    rom[5734] = 25'b0000000010110010000011001;
    rom[5735] = 25'b0000000010101110110011010;
    rom[5736] = 25'b0000000010101011100010100;
    rom[5737] = 25'b0000000010101000010000111;
    rom[5738] = 25'b0000000010100100111110011;
    rom[5739] = 25'b0000000010100001101010111;
    rom[5740] = 25'b0000000010011110010110101;
    rom[5741] = 25'b0000000010011011000001100;
    rom[5742] = 25'b0000000010010111101011100;
    rom[5743] = 25'b0000000010010100010100101;
    rom[5744] = 25'b0000000010010000111101000;
    rom[5745] = 25'b0000000010001101100100011;
    rom[5746] = 25'b0000000010001010001011000;
    rom[5747] = 25'b0000000010000110110000110;
    rom[5748] = 25'b0000000010000011010101101;
    rom[5749] = 25'b0000000001111111111001110;
    rom[5750] = 25'b0000000001111100011101000;
    rom[5751] = 25'b0000000001111000111111011;
    rom[5752] = 25'b0000000001110101100001000;
    rom[5753] = 25'b0000000001110010000001111;
    rom[5754] = 25'b0000000001101110100001110;
    rom[5755] = 25'b0000000001101011000001000;
    rom[5756] = 25'b0000000001100111011111010;
    rom[5757] = 25'b0000000001100011111101000;
    rom[5758] = 25'b0000000001100000011001101;
    rom[5759] = 25'b0000000001011100110101110;
    rom[5760] = 25'b0000000001011001010001000;
    rom[5761] = 25'b0000000001010101101011011;
    rom[5762] = 25'b0000000001010010000101000;
    rom[5763] = 25'b0000000001001110011101111;
    rom[5764] = 25'b0000000001001010110110000;
    rom[5765] = 25'b0000000001000111001101100;
    rom[5766] = 25'b0000000001000011100100001;
    rom[5767] = 25'b0000000000111111111001111;
    rom[5768] = 25'b0000000000111100001111000;
    rom[5769] = 25'b0000000000111000100011100;
    rom[5770] = 25'b0000000000110100110111001;
    rom[5771] = 25'b0000000000110001001001111;
    rom[5772] = 25'b0000000000101101011100010;
    rom[5773] = 25'b0000000000101001101101101;
    rom[5774] = 25'b0000000000100101111110100;
    rom[5775] = 25'b0000000000100010001110100;
    rom[5776] = 25'b0000000000011110011101110;
    rom[5777] = 25'b0000000000011010101100100;
    rom[5778] = 25'b0000000000010110111010011;
    rom[5779] = 25'b0000000000010011000111110;
    rom[5780] = 25'b0000000000001111010100010;
    rom[5781] = 25'b0000000000001011100000001;
    rom[5782] = 25'b0000000000000111101011011;
    rom[5783] = 25'b0000000000000011110110000;
    rom[5784] = 25'b0000000000000000000000000;
    rom[5785] = 25'b1111111111111100001001010;
    rom[5786] = 25'b1111111111111000010001110;
    rom[5787] = 25'b1111111111110100011001110;
    rom[5788] = 25'b1111111111110000100001001;
    rom[5789] = 25'b1111111111101100100111110;
    rom[5790] = 25'b1111111111101000101101111;
    rom[5791] = 25'b1111111111100100110011010;
    rom[5792] = 25'b1111111111100000111000001;
    rom[5793] = 25'b1111111111011100111100011;
    rom[5794] = 25'b1111111111011001000000000;
    rom[5795] = 25'b1111111111010101000011000;
    rom[5796] = 25'b1111111111010001000101011;
    rom[5797] = 25'b1111111111001101000111010;
    rom[5798] = 25'b1111111111001001001000100;
    rom[5799] = 25'b1111111111000101001001010;
    rom[5800] = 25'b1111111111000001001001010;
    rom[5801] = 25'b1111111110111101001000111;
    rom[5802] = 25'b1111111110111001000111110;
    rom[5803] = 25'b1111111110110101000110011;
    rom[5804] = 25'b1111111110110001000100010;
    rom[5805] = 25'b1111111110101101000001100;
    rom[5806] = 25'b1111111110101000111110100;
    rom[5807] = 25'b1111111110100100111010110;
    rom[5808] = 25'b1111111110100000110110100;
    rom[5809] = 25'b1111111110011100110001110;
    rom[5810] = 25'b1111111110011000101100101;
    rom[5811] = 25'b1111111110010100100110111;
    rom[5812] = 25'b1111111110010000100000101;
    rom[5813] = 25'b1111111110001100011001111;
    rom[5814] = 25'b1111111110001000010010110;
    rom[5815] = 25'b1111111110000100001011001;
    rom[5816] = 25'b1111111110000000000010111;
    rom[5817] = 25'b1111111101111011111010010;
    rom[5818] = 25'b1111111101110111110001010;
    rom[5819] = 25'b1111111101110011100111110;
    rom[5820] = 25'b1111111101101111011101111;
    rom[5821] = 25'b1111111101101011010011100;
    rom[5822] = 25'b1111111101100111001000110;
    rom[5823] = 25'b1111111101100010111101100;
    rom[5824] = 25'b1111111101011110110001111;
    rom[5825] = 25'b1111111101011010100101111;
    rom[5826] = 25'b1111111101010110011001100;
    rom[5827] = 25'b1111111101010010001100101;
    rom[5828] = 25'b1111111101001101111111011;
    rom[5829] = 25'b1111111101001001110001110;
    rom[5830] = 25'b1111111101000101100011111;
    rom[5831] = 25'b1111111101000001010101100;
    rom[5832] = 25'b1111111100111101000110111;
    rom[5833] = 25'b1111111100111000110111111;
    rom[5834] = 25'b1111111100110100101000100;
    rom[5835] = 25'b1111111100110000011000110;
    rom[5836] = 25'b1111111100101100001000101;
    rom[5837] = 25'b1111111100100111111000011;
    rom[5838] = 25'b1111111100100011100111110;
    rom[5839] = 25'b1111111100011111010110110;
    rom[5840] = 25'b1111111100011011000101011;
    rom[5841] = 25'b1111111100010110110011111;
    rom[5842] = 25'b1111111100010010100010000;
    rom[5843] = 25'b1111111100001110001111110;
    rom[5844] = 25'b1111111100001001111101011;
    rom[5845] = 25'b1111111100000101101010101;
    rom[5846] = 25'b1111111100000001010111110;
    rom[5847] = 25'b1111111011111101000100100;
    rom[5848] = 25'b1111111011111000110001001;
    rom[5849] = 25'b1111111011110100011101100;
    rom[5850] = 25'b1111111011110000001001101;
    rom[5851] = 25'b1111111011101011110101011;
    rom[5852] = 25'b1111111011100111100001001;
    rom[5853] = 25'b1111111011100011001100101;
    rom[5854] = 25'b1111111011011110110111111;
    rom[5855] = 25'b1111111011011010100011000;
    rom[5856] = 25'b1111111011010110001101111;
    rom[5857] = 25'b1111111011010001111000101;
    rom[5858] = 25'b1111111011001101100011010;
    rom[5859] = 25'b1111111011001001001101101;
    rom[5860] = 25'b1111111011000100110111111;
    rom[5861] = 25'b1111111011000000100010000;
    rom[5862] = 25'b1111111010111100001100000;
    rom[5863] = 25'b1111111010110111110101111;
    rom[5864] = 25'b1111111010110011011111101;
    rom[5865] = 25'b1111111010101111001001010;
    rom[5866] = 25'b1111111010101010110010110;
    rom[5867] = 25'b1111111010100110011100010;
    rom[5868] = 25'b1111111010100010000101101;
    rom[5869] = 25'b1111111010011101101110111;
    rom[5870] = 25'b1111111010011001011000000;
    rom[5871] = 25'b1111111010010101000001001;
    rom[5872] = 25'b1111111010010000101010010;
    rom[5873] = 25'b1111111010001100010011010;
    rom[5874] = 25'b1111111010000111111100010;
    rom[5875] = 25'b1111111010000011100101001;
    rom[5876] = 25'b1111111001111111001110010;
    rom[5877] = 25'b1111111001111010110111001;
    rom[5878] = 25'b1111111001110110100000000;
    rom[5879] = 25'b1111111001110010001000111;
    rom[5880] = 25'b1111111001101101110001111;
    rom[5881] = 25'b1111111001101001011010111;
    rom[5882] = 25'b1111111001100101000011110;
    rom[5883] = 25'b1111111001100000101100110;
    rom[5884] = 25'b1111111001011100010101111;
    rom[5885] = 25'b1111111001010111111111000;
    rom[5886] = 25'b1111111001010011101000001;
    rom[5887] = 25'b1111111001001111010001011;
    rom[5888] = 25'b1111111001001010111010110;
    rom[5889] = 25'b1111111001000110100100001;
    rom[5890] = 25'b1111111001000010001101101;
    rom[5891] = 25'b1111111000111101110111010;
    rom[5892] = 25'b1111111000111001100001000;
    rom[5893] = 25'b1111111000110101001010110;
    rom[5894] = 25'b1111111000110000110100110;
    rom[5895] = 25'b1111111000101100011110111;
    rom[5896] = 25'b1111111000101000001001001;
    rom[5897] = 25'b1111111000100011110011100;
    rom[5898] = 25'b1111111000011111011110000;
    rom[5899] = 25'b1111111000011011001000110;
    rom[5900] = 25'b1111111000010110110011110;
    rom[5901] = 25'b1111111000010010011110110;
    rom[5902] = 25'b1111111000001110001010000;
    rom[5903] = 25'b1111111000001001110101101;
    rom[5904] = 25'b1111111000000101100001011;
    rom[5905] = 25'b1111111000000001001101010;
    rom[5906] = 25'b1111110111111100111001100;
    rom[5907] = 25'b1111110111111000100101110;
    rom[5908] = 25'b1111110111110100010010100;
    rom[5909] = 25'b1111110111101111111111011;
    rom[5910] = 25'b1111110111101011101100101;
    rom[5911] = 25'b1111110111100111011010001;
    rom[5912] = 25'b1111110111100011000111111;
    rom[5913] = 25'b1111110111011110110101111;
    rom[5914] = 25'b1111110111011010100100010;
    rom[5915] = 25'b1111110111010110010010111;
    rom[5916] = 25'b1111110111010010000001111;
    rom[5917] = 25'b1111110111001101110001001;
    rom[5918] = 25'b1111110111001001100000110;
    rom[5919] = 25'b1111110111000101010000110;
    rom[5920] = 25'b1111110111000001000001001;
    rom[5921] = 25'b1111110110111100110001110;
    rom[5922] = 25'b1111110110111000100010111;
    rom[5923] = 25'b1111110110110100010100011;
    rom[5924] = 25'b1111110110110000000110001;
    rom[5925] = 25'b1111110110101011111000011;
    rom[5926] = 25'b1111110110100111101011001;
    rom[5927] = 25'b1111110110100011011110001;
    rom[5928] = 25'b1111110110011111010001110;
    rom[5929] = 25'b1111110110011011000101101;
    rom[5930] = 25'b1111110110010110111010000;
    rom[5931] = 25'b1111110110010010101110111;
    rom[5932] = 25'b1111110110001110100100001;
    rom[5933] = 25'b1111110110001010011001111;
    rom[5934] = 25'b1111110110000110010000001;
    rom[5935] = 25'b1111110110000010000110111;
    rom[5936] = 25'b1111110101111101111110001;
    rom[5937] = 25'b1111110101111001110101111;
    rom[5938] = 25'b1111110101110101101110010;
    rom[5939] = 25'b1111110101110001100111000;
    rom[5940] = 25'b1111110101101101100000010;
    rom[5941] = 25'b1111110101101001011010010;
    rom[5942] = 25'b1111110101100101010100101;
    rom[5943] = 25'b1111110101100001001111101;
    rom[5944] = 25'b1111110101011101001011001;
    rom[5945] = 25'b1111110101011001000111010;
    rom[5946] = 25'b1111110101010101000100001;
    rom[5947] = 25'b1111110101010001000001011;
    rom[5948] = 25'b1111110101001100111111010;
    rom[5949] = 25'b1111110101001000111101111;
    rom[5950] = 25'b1111110101000100111101001;
    rom[5951] = 25'b1111110101000000111100111;
    rom[5952] = 25'b1111110100111100111101011;
    rom[5953] = 25'b1111110100111000111110101;
    rom[5954] = 25'b1111110100110101000000010;
    rom[5955] = 25'b1111110100110001000010111;
    rom[5956] = 25'b1111110100101101000101111;
    rom[5957] = 25'b1111110100101001001001110;
    rom[5958] = 25'b1111110100100101001110010;
    rom[5959] = 25'b1111110100100001010011100;
    rom[5960] = 25'b1111110100011101011001101;
    rom[5961] = 25'b1111110100011001100000010;
    rom[5962] = 25'b1111110100010101100111110;
    rom[5963] = 25'b1111110100010001101111111;
    rom[5964] = 25'b1111110100001101111000111;
    rom[5965] = 25'b1111110100001010000010100;
    rom[5966] = 25'b1111110100000110001100111;
    rom[5967] = 25'b1111110100000010011000010;
    rom[5968] = 25'b1111110011111110100100010;
    rom[5969] = 25'b1111110011111010110001001;
    rom[5970] = 25'b1111110011110110111110110;
    rom[5971] = 25'b1111110011110011001101011;
    rom[5972] = 25'b1111110011101111011100101;
    rom[5973] = 25'b1111110011101011101100111;
    rom[5974] = 25'b1111110011100111111101111;
    rom[5975] = 25'b1111110011100100001111101;
    rom[5976] = 25'b1111110011100000100010011;
    rom[5977] = 25'b1111110011011100110110000;
    rom[5978] = 25'b1111110011011001001010100;
    rom[5979] = 25'b1111110011010101011111111;
    rom[5980] = 25'b1111110011010001110110001;
    rom[5981] = 25'b1111110011001110001101011;
    rom[5982] = 25'b1111110011001010100101100;
    rom[5983] = 25'b1111110011000110111110100;
    rom[5984] = 25'b1111110011000011011000100;
    rom[5985] = 25'b1111110010111111110011011;
    rom[5986] = 25'b1111110010111100001111011;
    rom[5987] = 25'b1111110010111000101100001;
    rom[5988] = 25'b1111110010110101001010000;
    rom[5989] = 25'b1111110010110001101000111;
    rom[5990] = 25'b1111110010101110001000101;
    rom[5991] = 25'b1111110010101010101001100;
    rom[5992] = 25'b1111110010100111001011011;
    rom[5993] = 25'b1111110010100011101110010;
    rom[5994] = 25'b1111110010100000010010001;
    rom[5995] = 25'b1111110010011100110111000;
    rom[5996] = 25'b1111110010011001011101001;
    rom[5997] = 25'b1111110010010110000100001;
    rom[5998] = 25'b1111110010010010101100001;
    rom[5999] = 25'b1111110010001111010101011;
    rom[6000] = 25'b1111110010001011111111101;
    rom[6001] = 25'b1111110010001000101011000;
    rom[6002] = 25'b1111110010000101010111100;
    rom[6003] = 25'b1111110010000010000101000;
    rom[6004] = 25'b1111110001111110110011111;
    rom[6005] = 25'b1111110001111011100011101;
    rom[6006] = 25'b1111110001111000010100101;
    rom[6007] = 25'b1111110001110101000110110;
    rom[6008] = 25'b1111110001110001111010001;
    rom[6009] = 25'b1111110001101110101110100;
    rom[6010] = 25'b1111110001101011100100001;
    rom[6011] = 25'b1111110001101000011011000;
    rom[6012] = 25'b1111110001100101010011000;
    rom[6013] = 25'b1111110001100010001100001;
    rom[6014] = 25'b1111110001011111000110101;
    rom[6015] = 25'b1111110001011100000010010;
    rom[6016] = 25'b1111110001011000111111001;
    rom[6017] = 25'b1111110001010101111101010;
    rom[6018] = 25'b1111110001010010111100101;
    rom[6019] = 25'b1111110001001111111101010;
    rom[6020] = 25'b1111110001001100111111001;
    rom[6021] = 25'b1111110001001010000010010;
    rom[6022] = 25'b1111110001000111000110110;
    rom[6023] = 25'b1111110001000100001100100;
    rom[6024] = 25'b1111110001000001010011100;
    rom[6025] = 25'b1111110000111110011011110;
    rom[6026] = 25'b1111110000111011100101100;
    rom[6027] = 25'b1111110000111000110000011;
    rom[6028] = 25'b1111110000110101111100110;
    rom[6029] = 25'b1111110000110011001010100;
    rom[6030] = 25'b1111110000110000011001100;
    rom[6031] = 25'b1111110000101101101001111;
    rom[6032] = 25'b1111110000101010111011101;
    rom[6033] = 25'b1111110000101000001110110;
    rom[6034] = 25'b1111110000100101100011010;
    rom[6035] = 25'b1111110000100010111001001;
    rom[6036] = 25'b1111110000100000010000011;
    rom[6037] = 25'b1111110000011101101001010;
    rom[6038] = 25'b1111110000011011000011011;
    rom[6039] = 25'b1111110000011000011110111;
    rom[6040] = 25'b1111110000010101111011111;
    rom[6041] = 25'b1111110000010011011010011;
    rom[6042] = 25'b1111110000010000111010011;
    rom[6043] = 25'b1111110000001110011011110;
    rom[6044] = 25'b1111110000001011111110101;
    rom[6045] = 25'b1111110000001001100010111;
    rom[6046] = 25'b1111110000000111001000101;
    rom[6047] = 25'b1111110000000100110000000;
    rom[6048] = 25'b1111110000000010011000111;
    rom[6049] = 25'b1111110000000000000011001;
    rom[6050] = 25'b1111101111111101101111000;
    rom[6051] = 25'b1111101111111011011100100;
    rom[6052] = 25'b1111101111111001001011011;
    rom[6053] = 25'b1111101111110110111011110;
    rom[6054] = 25'b1111101111110100101101110;
    rom[6055] = 25'b1111101111110010100001100;
    rom[6056] = 25'b1111101111110000010110101;
    rom[6057] = 25'b1111101111101110001101010;
    rom[6058] = 25'b1111101111101100000101101;
    rom[6059] = 25'b1111101111101001111111100;
    rom[6060] = 25'b1111101111100111111011001;
    rom[6061] = 25'b1111101111100101111000010;
    rom[6062] = 25'b1111101111100011110110111;
    rom[6063] = 25'b1111101111100001110111010;
    rom[6064] = 25'b1111101111011111111001010;
    rom[6065] = 25'b1111101111011101111101000;
    rom[6066] = 25'b1111101111011100000010010;
    rom[6067] = 25'b1111101111011010001001010;
    rom[6068] = 25'b1111101111011000010001111;
    rom[6069] = 25'b1111101111010110011100001;
    rom[6070] = 25'b1111101111010100101000000;
    rom[6071] = 25'b1111101111010010110101110;
    rom[6072] = 25'b1111101111010001000101000;
    rom[6073] = 25'b1111101111001111010110001;
    rom[6074] = 25'b1111101111001101101001000;
    rom[6075] = 25'b1111101111001011111101011;
    rom[6076] = 25'b1111101111001010010011101;
    rom[6077] = 25'b1111101111001000101011101;
    rom[6078] = 25'b1111101111000111000101010;
    rom[6079] = 25'b1111101111000101100000110;
    rom[6080] = 25'b1111101111000011111101111;
    rom[6081] = 25'b1111101111000010011100111;
    rom[6082] = 25'b1111101111000000111101101;
    rom[6083] = 25'b1111101110111111100000001;
    rom[6084] = 25'b1111101110111110000100011;
    rom[6085] = 25'b1111101110111100101010100;
    rom[6086] = 25'b1111101110111011010010100;
    rom[6087] = 25'b1111101110111001111100001;
    rom[6088] = 25'b1111101110111000100111101;
    rom[6089] = 25'b1111101110110111010100111;
    rom[6090] = 25'b1111101110110110000100001;
    rom[6091] = 25'b1111101110110100110101001;
    rom[6092] = 25'b1111101110110011100111111;
    rom[6093] = 25'b1111101110110010011100100;
    rom[6094] = 25'b1111101110110001010011001;
    rom[6095] = 25'b1111101110110000001011100;
    rom[6096] = 25'b1111101110101111000101110;
    rom[6097] = 25'b1111101110101110000010000;
    rom[6098] = 25'b1111101110101101000000000;
    rom[6099] = 25'b1111101110101011111111111;
    rom[6100] = 25'b1111101110101011000001110;
    rom[6101] = 25'b1111101110101010000101011;
    rom[6102] = 25'b1111101110101001001011000;
    rom[6103] = 25'b1111101110101000010010100;
    rom[6104] = 25'b1111101110100111011100000;
    rom[6105] = 25'b1111101110100110100111011;
    rom[6106] = 25'b1111101110100101110100110;
    rom[6107] = 25'b1111101110100101000100000;
    rom[6108] = 25'b1111101110100100010101010;
    rom[6109] = 25'b1111101110100011101000100;
    rom[6110] = 25'b1111101110100010111101100;
    rom[6111] = 25'b1111101110100010010100110;
    rom[6112] = 25'b1111101110100001101101101;
    rom[6113] = 25'b1111101110100001001000110;
    rom[6114] = 25'b1111101110100000100101110;
    rom[6115] = 25'b1111101110100000000100111;
    rom[6116] = 25'b1111101110011111100101110;
    rom[6117] = 25'b1111101110011111001000111;
    rom[6118] = 25'b1111101110011110101101111;
    rom[6119] = 25'b1111101110011110010101000;
    rom[6120] = 25'b1111101110011101111110000;
    rom[6121] = 25'b1111101110011101101001001;
    rom[6122] = 25'b1111101110011101010110010;
    rom[6123] = 25'b1111101110011101000101011;
    rom[6124] = 25'b1111101110011100110110101;
    rom[6125] = 25'b1111101110011100101001111;
    rom[6126] = 25'b1111101110011100011111010;
    rom[6127] = 25'b1111101110011100010110100;
    rom[6128] = 25'b1111101110011100010000000;
    rom[6129] = 25'b1111101110011100001011100;
    rom[6130] = 25'b1111101110011100001001001;
    rom[6131] = 25'b1111101110011100001000110;
    rom[6132] = 25'b1111101110011100001010100;
    rom[6133] = 25'b1111101110011100001110010;
    rom[6134] = 25'b1111101110011100010100010;
    rom[6135] = 25'b1111101110011100011100011;
    rom[6136] = 25'b1111101110011100100110100;
    rom[6137] = 25'b1111101110011100110010101;
    rom[6138] = 25'b1111101110011101000001001;
    rom[6139] = 25'b1111101110011101010001101;
    rom[6140] = 25'b1111101110011101100100010;
    rom[6141] = 25'b1111101110011101111001000;
    rom[6142] = 25'b1111101110011110001111111;
    rom[6143] = 25'b1111101110011110101000111;
    rom[6144] = 25'b1111101110011111000100001;
    rom[6145] = 25'b1111101110011111100001100;
    rom[6146] = 25'b1111101110100000000000111;
    rom[6147] = 25'b1111101110100000100010100;
    rom[6148] = 25'b1111101110100001000110011;
    rom[6149] = 25'b1111101110100001101100010;
    rom[6150] = 25'b1111101110100010010100100;
    rom[6151] = 25'b1111101110100010111110110;
    rom[6152] = 25'b1111101110100011101011011;
    rom[6153] = 25'b1111101110100100011010000;
    rom[6154] = 25'b1111101110100101001010111;
    rom[6155] = 25'b1111101110100101111110000;
    rom[6156] = 25'b1111101110100110110011010;
    rom[6157] = 25'b1111101110100111101010110;
    rom[6158] = 25'b1111101110101000100100011;
    rom[6159] = 25'b1111101110101001100000010;
    rom[6160] = 25'b1111101110101010011110011;
    rom[6161] = 25'b1111101110101011011110101;
    rom[6162] = 25'b1111101110101100100001010;
    rom[6163] = 25'b1111101110101101100110000;
    rom[6164] = 25'b1111101110101110101101000;
    rom[6165] = 25'b1111101110101111110110001;
    rom[6166] = 25'b1111101110110001000001101;
    rom[6167] = 25'b1111101110110010001111011;
    rom[6168] = 25'b1111101110110011011111011;
    rom[6169] = 25'b1111101110110100110001100;
    rom[6170] = 25'b1111101110110110000101111;
    rom[6171] = 25'b1111101110110111011100100;
    rom[6172] = 25'b1111101110111000110101100;
    rom[6173] = 25'b1111101110111010010000101;
    rom[6174] = 25'b1111101110111011101110001;
    rom[6175] = 25'b1111101110111101001101111;
    rom[6176] = 25'b1111101110111110101111110;
    rom[6177] = 25'b1111101111000000010100000;
    rom[6178] = 25'b1111101111000001111010101;
    rom[6179] = 25'b1111101111000011100011011;
    rom[6180] = 25'b1111101111000101001110100;
    rom[6181] = 25'b1111101111000110111011110;
    rom[6182] = 25'b1111101111001000101011100;
    rom[6183] = 25'b1111101111001010011101011;
    rom[6184] = 25'b1111101111001100010001101;
    rom[6185] = 25'b1111101111001110001000000;
    rom[6186] = 25'b1111101111010000000000110;
    rom[6187] = 25'b1111101111010001111011111;
    rom[6188] = 25'b1111101111010011111001010;
    rom[6189] = 25'b1111101111010101111001000;
    rom[6190] = 25'b1111101111010111111011000;
    rom[6191] = 25'b1111101111011001111111010;
    rom[6192] = 25'b1111101111011100000101110;
    rom[6193] = 25'b1111101111011110001110101;
    rom[6194] = 25'b1111101111100000011001111;
    rom[6195] = 25'b1111101111100010100111011;
    rom[6196] = 25'b1111101111100100110111001;
    rom[6197] = 25'b1111101111100111001001010;
    rom[6198] = 25'b1111101111101001011101110;
    rom[6199] = 25'b1111101111101011110100100;
    rom[6200] = 25'b1111101111101110001101101;
    rom[6201] = 25'b1111101111110000101000111;
    rom[6202] = 25'b1111101111110011000110101;
    rom[6203] = 25'b1111101111110101100110101;
    rom[6204] = 25'b1111101111111000001001000;
    rom[6205] = 25'b1111101111111010101101101;
    rom[6206] = 25'b1111101111111101010100101;
    rom[6207] = 25'b1111101111111111111101111;
    rom[6208] = 25'b1111110000000010101001101;
    rom[6209] = 25'b1111110000000101010111100;
    rom[6210] = 25'b1111110000001000000111111;
    rom[6211] = 25'b1111110000001010111010100;
    rom[6212] = 25'b1111110000001101101111100;
    rom[6213] = 25'b1111110000010000100110110;
    rom[6214] = 25'b1111110000010011100000010;
    rom[6215] = 25'b1111110000010110011100010;
    rom[6216] = 25'b1111110000011001011010100;
    rom[6217] = 25'b1111110000011100011011001;
    rom[6218] = 25'b1111110000011111011110000;
    rom[6219] = 25'b1111110000100010100011011;
    rom[6220] = 25'b1111110000100101101010111;
    rom[6221] = 25'b1111110000101000110100110;
    rom[6222] = 25'b1111110000101100000001000;
    rom[6223] = 25'b1111110000101111001111110;
    rom[6224] = 25'b1111110000110010100000101;
    rom[6225] = 25'b1111110000110101110011111;
    rom[6226] = 25'b1111110000111001001001011;
    rom[6227] = 25'b1111110000111100100001010;
    rom[6228] = 25'b1111110000111111111011100;
    rom[6229] = 25'b1111110001000011011000001;
    rom[6230] = 25'b1111110001000110110110111;
    rom[6231] = 25'b1111110001001010011000010;
    rom[6232] = 25'b1111110001001101111011110;
    rom[6233] = 25'b1111110001010001100001100;
    rom[6234] = 25'b1111110001010101001001110;
    rom[6235] = 25'b1111110001011000110100010;
    rom[6236] = 25'b1111110001011100100001000;
    rom[6237] = 25'b1111110001100000010000010;
    rom[6238] = 25'b1111110001100100000001101;
    rom[6239] = 25'b1111110001100111110101011;
    rom[6240] = 25'b1111110001101011101011100;
    rom[6241] = 25'b1111110001101111100100000;
    rom[6242] = 25'b1111110001110011011110110;
    rom[6243] = 25'b1111110001110111011011110;
    rom[6244] = 25'b1111110001111011011011001;
    rom[6245] = 25'b1111110001111111011100111;
    rom[6246] = 25'b1111110010000011100000110;
    rom[6247] = 25'b1111110010000111100111001;
    rom[6248] = 25'b1111110010001011101111110;
    rom[6249] = 25'b1111110010001111111010100;
    rom[6250] = 25'b1111110010010100000111110;
    rom[6251] = 25'b1111110010011000010111010;
    rom[6252] = 25'b1111110010011100101001000;
    rom[6253] = 25'b1111110010100000111101001;
    rom[6254] = 25'b1111110010100101010011100;
    rom[6255] = 25'b1111110010101001101100001;
    rom[6256] = 25'b1111110010101110000111001;
    rom[6257] = 25'b1111110010110010100100010;
    rom[6258] = 25'b1111110010110111000011110;
    rom[6259] = 25'b1111110010111011100101101;
    rom[6260] = 25'b1111110011000000001001101;
    rom[6261] = 25'b1111110011000100110000000;
    rom[6262] = 25'b1111110011001001011000101;
    rom[6263] = 25'b1111110011001110000011100;
    rom[6264] = 25'b1111110011010010110000101;
    rom[6265] = 25'b1111110011010111100000000;
    rom[6266] = 25'b1111110011011100010001110;
    rom[6267] = 25'b1111110011100001000101101;
    rom[6268] = 25'b1111110011100101111011110;
    rom[6269] = 25'b1111110011101010110100001;
    rom[6270] = 25'b1111110011101111101110111;
    rom[6271] = 25'b1111110011110100101011101;
    rom[6272] = 25'b1111110011111001101010110;
    rom[6273] = 25'b1111110011111110101100001;
    rom[6274] = 25'b1111110100000011101111110;
    rom[6275] = 25'b1111110100001000110101100;
    rom[6276] = 25'b1111110100001101111101101;
    rom[6277] = 25'b1111110100010011000111111;
    rom[6278] = 25'b1111110100011000010100011;
    rom[6279] = 25'b1111110100011101100011000;
    rom[6280] = 25'b1111110100100010110011111;
    rom[6281] = 25'b1111110100101000000111000;
    rom[6282] = 25'b1111110100101101011100010;
    rom[6283] = 25'b1111110100110010110011110;
    rom[6284] = 25'b1111110100111000001101011;
    rom[6285] = 25'b1111110100111101101001010;
    rom[6286] = 25'b1111110101000011000111001;
    rom[6287] = 25'b1111110101001000100111011;
    rom[6288] = 25'b1111110101001110001001110;
    rom[6289] = 25'b1111110101010011101110010;
    rom[6290] = 25'b1111110101011001010100111;
    rom[6291] = 25'b1111110101011110111101110;
    rom[6292] = 25'b1111110101100100101000101;
    rom[6293] = 25'b1111110101101010010101111;
    rom[6294] = 25'b1111110101110000000101000;
    rom[6295] = 25'b1111110101110101110110100;
    rom[6296] = 25'b1111110101111011101010000;
    rom[6297] = 25'b1111110110000001011111101;
    rom[6298] = 25'b1111110110000111010111011;
    rom[6299] = 25'b1111110110001101010001001;
    rom[6300] = 25'b1111110110010011001101001;
    rom[6301] = 25'b1111110110011001001011010;
    rom[6302] = 25'b1111110110011111001011011;
    rom[6303] = 25'b1111110110100101001101100;
    rom[6304] = 25'b1111110110101011010001111;
    rom[6305] = 25'b1111110110110001011000010;
    rom[6306] = 25'b1111110110110111100000110;
    rom[6307] = 25'b1111110110111101101011011;
    rom[6308] = 25'b1111110111000011110111111;
    rom[6309] = 25'b1111110111001010000110011;
    rom[6310] = 25'b1111110111010000010111001;
    rom[6311] = 25'b1111110111010110101001111;
    rom[6312] = 25'b1111110111011100111110101;
    rom[6313] = 25'b1111110111100011010101011;
    rom[6314] = 25'b1111110111101001101110001;
    rom[6315] = 25'b1111110111110000001000111;
    rom[6316] = 25'b1111110111110110100101101;
    rom[6317] = 25'b1111110111111101000100011;
    rom[6318] = 25'b1111111000000011100101001;
    rom[6319] = 25'b1111111000001010000111111;
    rom[6320] = 25'b1111111000010000101100101;
    rom[6321] = 25'b1111111000010111010011010;
    rom[6322] = 25'b1111111000011101111011111;
    rom[6323] = 25'b1111111000100100100110011;
    rom[6324] = 25'b1111111000101011010011000;
    rom[6325] = 25'b1111111000110010000001011;
    rom[6326] = 25'b1111111000111000110001110;
    rom[6327] = 25'b1111111000111111100100001;
    rom[6328] = 25'b1111111001000110011000010;
    rom[6329] = 25'b1111111001001101001110100;
    rom[6330] = 25'b1111111001010100000110011;
    rom[6331] = 25'b1111111001011011000000011;
    rom[6332] = 25'b1111111001100001111100001;
    rom[6333] = 25'b1111111001101000111001110;
    rom[6334] = 25'b1111111001101111111001011;
    rom[6335] = 25'b1111111001110110111010110;
    rom[6336] = 25'b1111111001111101111101111;
    rom[6337] = 25'b1111111010000101000011000;
    rom[6338] = 25'b1111111010001100001001111;
    rom[6339] = 25'b1111111010010011010010100;
    rom[6340] = 25'b1111111010011010011101001;
    rom[6341] = 25'b1111111010100001101001011;
    rom[6342] = 25'b1111111010101000110111100;
    rom[6343] = 25'b1111111010110000000111011;
    rom[6344] = 25'b1111111010110111011001000;
    rom[6345] = 25'b1111111010111110101100100;
    rom[6346] = 25'b1111111011000110000001110;
    rom[6347] = 25'b1111111011001101011000110;
    rom[6348] = 25'b1111111011010100110001011;
    rom[6349] = 25'b1111111011011100001011110;
    rom[6350] = 25'b1111111011100011100111111;
    rom[6351] = 25'b1111111011101011000101110;
    rom[6352] = 25'b1111111011110010100101010;
    rom[6353] = 25'b1111111011111010000110100;
    rom[6354] = 25'b1111111100000001101001011;
    rom[6355] = 25'b1111111100001001001110000;
    rom[6356] = 25'b1111111100010000110100010;
    rom[6357] = 25'b1111111100011000011100001;
    rom[6358] = 25'b1111111100100000000101101;
    rom[6359] = 25'b1111111100100111110000111;
    rom[6360] = 25'b1111111100101111011101110;
    rom[6361] = 25'b1111111100110111001100000;
    rom[6362] = 25'b1111111100111110111100001;
    rom[6363] = 25'b1111111101000110101101101;
    rom[6364] = 25'b1111111101001110100000110;
    rom[6365] = 25'b1111111101010110010101101;
    rom[6366] = 25'b1111111101011110001011111;
    rom[6367] = 25'b1111111101100110000011110;
    rom[6368] = 25'b1111111101101101111101001;
    rom[6369] = 25'b1111111101110101111000000;
    rom[6370] = 25'b1111111101111101110100100;
    rom[6371] = 25'b1111111110000101110010011;
    rom[6372] = 25'b1111111110001101110001110;
    rom[6373] = 25'b1111111110010101110010101;
    rom[6374] = 25'b1111111110011101110101001;
    rom[6375] = 25'b1111111110100101111000111;
    rom[6376] = 25'b1111111110101101111110001;
    rom[6377] = 25'b1111111110110110000100111;
    rom[6378] = 25'b1111111110111110001101000;
    rom[6379] = 25'b1111111111000110010110101;
    rom[6380] = 25'b1111111111001110100001100;
    rom[6381] = 25'b1111111111010110101101111;
    rom[6382] = 25'b1111111111011110111011101;
    rom[6383] = 25'b1111111111100111001010101;
    rom[6384] = 25'b1111111111101111011011000;
    rom[6385] = 25'b1111111111110111101100111;
    rom[6386] = 25'b0000000000000000000000000;
    rom[6387] = 25'b0000000000001000010100011;
    rom[6388] = 25'b0000000000010000101010000;
    rom[6389] = 25'b0000000000011001000001001;
    rom[6390] = 25'b0000000000100001011001011;
    rom[6391] = 25'b0000000000101001110011000;
    rom[6392] = 25'b0000000000110010001101110;
    rom[6393] = 25'b0000000000111010101001111;
    rom[6394] = 25'b0000000001000011000111001;
    rom[6395] = 25'b0000000001001011100101110;
    rom[6396] = 25'b0000000001010100000101100;
    rom[6397] = 25'b0000000001011100100110011;
    rom[6398] = 25'b0000000001100101001000100;
    rom[6399] = 25'b0000000001101101101011110;
    rom[6400] = 25'b0000000001110110010000010;
    rom[6401] = 25'b0000000001111110110101111;
    rom[6402] = 25'b0000000010000111011100100;
    rom[6403] = 25'b0000000010010000000100010;
    rom[6404] = 25'b0000000010011000101101010;
    rom[6405] = 25'b0000000010100001010111010;
    rom[6406] = 25'b0000000010101010000010010;
    rom[6407] = 25'b0000000010110010101110100;
    rom[6408] = 25'b0000000010111011011011101;
    rom[6409] = 25'b0000000011000100001001111;
    rom[6410] = 25'b0000000011001100111001001;
    rom[6411] = 25'b0000000011010101101001011;
    rom[6412] = 25'b0000000011011110011010101;
    rom[6413] = 25'b0000000011100111001100111;
    rom[6414] = 25'b0000000011110000000000000;
    rom[6415] = 25'b0000000011111000110100010;
    rom[6416] = 25'b0000000100000001101001010;
    rom[6417] = 25'b0000000100001010011111010;
    rom[6418] = 25'b0000000100010011010110010;
    rom[6419] = 25'b0000000100011100001110001;
    rom[6420] = 25'b0000000100100101000110110;
    rom[6421] = 25'b0000000100101110000000010;
    rom[6422] = 25'b0000000100110110111010110;
    rom[6423] = 25'b0000000100111111110110000;
    rom[6424] = 25'b0000000101001000110010000;
    rom[6425] = 25'b0000000101010001101110111;
    rom[6426] = 25'b0000000101011010101100101;
    rom[6427] = 25'b0000000101100011101011001;
    rom[6428] = 25'b0000000101101100101010011;
    rom[6429] = 25'b0000000101110101101010011;
    rom[6430] = 25'b0000000101111110101011000;
    rom[6431] = 25'b0000000110000111101100100;
    rom[6432] = 25'b0000000110010000101110101;
    rom[6433] = 25'b0000000110011001110001100;
    rom[6434] = 25'b0000000110100010110101000;
    rom[6435] = 25'b0000000110101011111001001;
    rom[6436] = 25'b0000000110110100111101111;
    rom[6437] = 25'b0000000110111110000011100;
    rom[6438] = 25'b0000000111000111001001100;
    rom[6439] = 25'b0000000111010000010000001;
    rom[6440] = 25'b0000000111011001010111011;
    rom[6441] = 25'b0000000111100010011111001;
    rom[6442] = 25'b0000000111101011100111101;
    rom[6443] = 25'b0000000111110100110000100;
    rom[6444] = 25'b0000000111111101111001111;
    rom[6445] = 25'b0000001000000111000011111;
    rom[6446] = 25'b0000001000010000001110010;
    rom[6447] = 25'b0000001000011001011001010;
    rom[6448] = 25'b0000001000100010100100101;
    rom[6449] = 25'b0000001000101011110000011;
    rom[6450] = 25'b0000001000110100111100101;
    rom[6451] = 25'b0000001000111110001001010;
    rom[6452] = 25'b0000001001000111010110011;
    rom[6453] = 25'b0000001001010000100011110;
    rom[6454] = 25'b0000001001011001110001101;
    rom[6455] = 25'b0000001001100010111111110;
    rom[6456] = 25'b0000001001101100001110001;
    rom[6457] = 25'b0000001001110101011101000;
    rom[6458] = 25'b0000001001111110101100000;
    rom[6459] = 25'b0000001010000111111011100;
    rom[6460] = 25'b0000001010010001001011001;
    rom[6461] = 25'b0000001010011010011010111;
    rom[6462] = 25'b0000001010100011101011001;
    rom[6463] = 25'b0000001010101100111011011;
    rom[6464] = 25'b0000001010110110001100000;
    rom[6465] = 25'b0000001010111111011100101;
    rom[6466] = 25'b0000001011001000101101100;
    rom[6467] = 25'b0000001011010001111110100;
    rom[6468] = 25'b0000001011011011001111110;
    rom[6469] = 25'b0000001011100100100001000;
    rom[6470] = 25'b0000001011101101110010011;
    rom[6471] = 25'b0000001011110111000011111;
    rom[6472] = 25'b0000001100000000010101011;
    rom[6473] = 25'b0000001100001001100111000;
    rom[6474] = 25'b0000001100010010111000110;
    rom[6475] = 25'b0000001100011100001010010;
    rom[6476] = 25'b0000001100100101011011111;
    rom[6477] = 25'b0000001100101110101101100;
    rom[6478] = 25'b0000001100110111111111001;
    rom[6479] = 25'b0000001101000001010000101;
    rom[6480] = 25'b0000001101001010100010000;
    rom[6481] = 25'b0000001101010011110011100;
    rom[6482] = 25'b0000001101011101000100110;
    rom[6483] = 25'b0000001101100110010101111;
    rom[6484] = 25'b0000001101101111100110111;
    rom[6485] = 25'b0000001101111000110111101;
    rom[6486] = 25'b0000001110000010001000011;
    rom[6487] = 25'b0000001110001011011000110;
    rom[6488] = 25'b0000001110010100101001001;
    rom[6489] = 25'b0000001110011101111001001;
    rom[6490] = 25'b0000001110100111001000111;
    rom[6491] = 25'b0000001110110000011000011;
    rom[6492] = 25'b0000001110111001100111101;
    rom[6493] = 25'b0000001111000010110110101;
    rom[6494] = 25'b0000001111001100000101010;
    rom[6495] = 25'b0000001111010101010011100;
    rom[6496] = 25'b0000001111011110100001011;
    rom[6497] = 25'b0000001111100111101111000;
    rom[6498] = 25'b0000001111110000111100010;
    rom[6499] = 25'b0000001111111010001001000;
    rom[6500] = 25'b0000010000000011010101011;
    rom[6501] = 25'b0000010000001100100001010;
    rom[6502] = 25'b0000010000010101101100101;
    rom[6503] = 25'b0000010000011110110111101;
    rom[6504] = 25'b0000010000101000000010001;
    rom[6505] = 25'b0000010000110001001100001;
    rom[6506] = 25'b0000010000111010010101100;
    rom[6507] = 25'b0000010001000011011110011;
    rom[6508] = 25'b0000010001001100100110110;
    rom[6509] = 25'b0000010001010101101110100;
    rom[6510] = 25'b0000010001011110110101101;
    rom[6511] = 25'b0000010001100111111100001;
    rom[6512] = 25'b0000010001110001000001111;
    rom[6513] = 25'b0000010001111010000111001;
    rom[6514] = 25'b0000010010000011001011101;
    rom[6515] = 25'b0000010010001100001111100;
    rom[6516] = 25'b0000010010010101010010100;
    rom[6517] = 25'b0000010010011110010101000;
    rom[6518] = 25'b0000010010100111010110100;
    rom[6519] = 25'b0000010010110000010111011;
    rom[6520] = 25'b0000010010111001010111011;
    rom[6521] = 25'b0000010011000010010110101;
    rom[6522] = 25'b0000010011001011010101001;
    rom[6523] = 25'b0000010011010100010010110;
    rom[6524] = 25'b0000010011011101001111011;
    rom[6525] = 25'b0000010011100110001011001;
    rom[6526] = 25'b0000010011101111000110001;
    rom[6527] = 25'b0000010011111000000000001;
    rom[6528] = 25'b0000010100000000111001010;
    rom[6529] = 25'b0000010100001001110001011;
    rom[6530] = 25'b0000010100010010101000100;
    rom[6531] = 25'b0000010100011011011110101;
    rom[6532] = 25'b0000010100100100010011110;
    rom[6533] = 25'b0000010100101101000111111;
    rom[6534] = 25'b0000010100110101111010111;
    rom[6535] = 25'b0000010100111110101100111;
    rom[6536] = 25'b0000010101000111011101110;
    rom[6537] = 25'b0000010101010000001101100;
    rom[6538] = 25'b0000010101011000111100010;
    rom[6539] = 25'b0000010101100001101001110;
    rom[6540] = 25'b0000010101101010010110001;
    rom[6541] = 25'b0000010101110011000001010;
    rom[6542] = 25'b0000010101111011101011001;
    rom[6543] = 25'b0000010110000100010100000;
    rom[6544] = 25'b0000010110001100111011100;
    rom[6545] = 25'b0000010110010101100001110;
    rom[6546] = 25'b0000010110011110000110110;
    rom[6547] = 25'b0000010110100110101010011;
    rom[6548] = 25'b0000010110101111001100110;
    rom[6549] = 25'b0000010110110111101101110;
    rom[6550] = 25'b0000010111000000001101011;
    rom[6551] = 25'b0000010111001000101011110;
    rom[6552] = 25'b0000010111010001001000101;
    rom[6553] = 25'b0000010111011001100100001;
    rom[6554] = 25'b0000010111100001111110010;
    rom[6555] = 25'b0000010111101010010110111;
    rom[6556] = 25'b0000010111110010101110000;
    rom[6557] = 25'b0000010111111011000011110;
    rom[6558] = 25'b0000011000000011010111111;
    rom[6559] = 25'b0000011000001011101010100;
    rom[6560] = 25'b0000011000010011111011101;
    rom[6561] = 25'b0000011000011100001011001;
    rom[6562] = 25'b0000011000100100011001001;
    rom[6563] = 25'b0000011000101100100101100;
    rom[6564] = 25'b0000011000110100110000010;
    rom[6565] = 25'b0000011000111100111001011;
    rom[6566] = 25'b0000011001000101000000111;
    rom[6567] = 25'b0000011001001101000110101;
    rom[6568] = 25'b0000011001010101001010101;
    rom[6569] = 25'b0000011001011101001101001;
    rom[6570] = 25'b0000011001100101001101110;
    rom[6571] = 25'b0000011001101101001100100;
    rom[6572] = 25'b0000011001110101001001110;
    rom[6573] = 25'b0000011001111101000101000;
    rom[6574] = 25'b0000011010000100111110100;
    rom[6575] = 25'b0000011010001100110110010;
    rom[6576] = 25'b0000011010010100101100000;
    rom[6577] = 25'b0000011010011100100000000;
    rom[6578] = 25'b0000011010100100010010001;
    rom[6579] = 25'b0000011010101100000010011;
    rom[6580] = 25'b0000011010110011110000101;
    rom[6581] = 25'b0000011010111011011100111;
    rom[6582] = 25'b0000011011000011000111010;
    rom[6583] = 25'b0000011011001010101111101;
    rom[6584] = 25'b0000011011010010010110000;
    rom[6585] = 25'b0000011011011001111010100;
    rom[6586] = 25'b0000011011100001011100111;
    rom[6587] = 25'b0000011011101000111101000;
    rom[6588] = 25'b0000011011110000011011010;
    rom[6589] = 25'b0000011011110111110111011;
    rom[6590] = 25'b0000011011111111010001100;
    rom[6591] = 25'b0000011100000110101001010;
    rom[6592] = 25'b0000011100001101111111000;
    rom[6593] = 25'b0000011100010101010010101;
    rom[6594] = 25'b0000011100011100100100000;
    rom[6595] = 25'b0000011100100011110011001;
    rom[6596] = 25'b0000011100101011000000001;
    rom[6597] = 25'b0000011100110010001010111;
    rom[6598] = 25'b0000011100111001010011010;
    rom[6599] = 25'b0000011101000000011001011;
    rom[6600] = 25'b0000011101000111011101011;
    rom[6601] = 25'b0000011101001110011110111;
    rom[6602] = 25'b0000011101010101011110001;
    rom[6603] = 25'b0000011101011100011010111;
    rom[6604] = 25'b0000011101100011010101100;
    rom[6605] = 25'b0000011101101010001101100;
    rom[6606] = 25'b0000011101110001000011010;
    rom[6607] = 25'b0000011101110111110110100;
    rom[6608] = 25'b0000011101111110100111011;
    rom[6609] = 25'b0000011110000101010101110;
    rom[6610] = 25'b0000011110001100000001101;
    rom[6611] = 25'b0000011110010010101011000;
    rom[6612] = 25'b0000011110011001010001111;
    rom[6613] = 25'b0000011110011111110110001;
    rom[6614] = 25'b0000011110100110010111111;
    rom[6615] = 25'b0000011110101100110111001;
    rom[6616] = 25'b0000011110110011010011101;
    rom[6617] = 25'b0000011110111001101101110;
    rom[6618] = 25'b0000011111000000000101000;
    rom[6619] = 25'b0000011111000110011001110;
    rom[6620] = 25'b0000011111001100101011110;
    rom[6621] = 25'b0000011111010010111011001;
    rom[6622] = 25'b0000011111011001000111110;
    rom[6623] = 25'b0000011111011111010001110;
    rom[6624] = 25'b0000011111100101011001000;
    rom[6625] = 25'b0000011111101011011101100;
    rom[6626] = 25'b0000011111110001011111000;
    rom[6627] = 25'b0000011111110111011110000;
    rom[6628] = 25'b0000011111111101011010000;
    rom[6629] = 25'b0000100000000011010011010;
    rom[6630] = 25'b0000100000001001001001101;
    rom[6631] = 25'b0000100000001110111101010;
    rom[6632] = 25'b0000100000010100101101111;
    rom[6633] = 25'b0000100000011010011011101;
    rom[6634] = 25'b0000100000100000000110100;
    rom[6635] = 25'b0000100000100101101110100;
    rom[6636] = 25'b0000100000101011010011100;
    rom[6637] = 25'b0000100000110000110101100;
    rom[6638] = 25'b0000100000110110010100011;
    rom[6639] = 25'b0000100000111011110000100;
    rom[6640] = 25'b0000100001000001001001100;
    rom[6641] = 25'b0000100001000110011111100;
    rom[6642] = 25'b0000100001001011110010010;
    rom[6643] = 25'b0000100001010001000010001;
    rom[6644] = 25'b0000100001010110001110111;
    rom[6645] = 25'b0000100001011011011000101;
    rom[6646] = 25'b0000100001100000011111000;
    rom[6647] = 25'b0000100001100101100010100;
    rom[6648] = 25'b0000100001101010100010101;
    rom[6649] = 25'b0000100001101111011111101;
    rom[6650] = 25'b0000100001110100011001101;
    rom[6651] = 25'b0000100001111001010000010;
    rom[6652] = 25'b0000100001111110000011101;
    rom[6653] = 25'b0000100010000010110011111;
    rom[6654] = 25'b0000100010000111100000110;
    rom[6655] = 25'b0000100010001100001010011;
    rom[6656] = 25'b0000100010010000110000110;
    rom[6657] = 25'b0000100010010101010011111;
    rom[6658] = 25'b0000100010011001110011101;
    rom[6659] = 25'b0000100010011110010000000;
    rom[6660] = 25'b0000100010100010101001000;
    rom[6661] = 25'b0000100010100110111110110;
    rom[6662] = 25'b0000100010101011010001000;
    rom[6663] = 25'b0000100010101111011111111;
    rom[6664] = 25'b0000100010110011101011010;
    rom[6665] = 25'b0000100010110111110011011;
    rom[6666] = 25'b0000100010111011110111111;
    rom[6667] = 25'b0000100010111111111001000;
    rom[6668] = 25'b0000100011000011110110101;
    rom[6669] = 25'b0000100011000111110000110;
    rom[6670] = 25'b0000100011001011100111011;
    rom[6671] = 25'b0000100011001111011010011;
    rom[6672] = 25'b0000100011010011001001111;
    rom[6673] = 25'b0000100011010110110101110;
    rom[6674] = 25'b0000100011011010011110010;
    rom[6675] = 25'b0000100011011110000011000;
    rom[6676] = 25'b0000100011100001100100001;
    rom[6677] = 25'b0000100011100101000001110;
    rom[6678] = 25'b0000100011101000011011100;
    rom[6679] = 25'b0000100011101011110001111;
    rom[6680] = 25'b0000100011101111000100011;
    rom[6681] = 25'b0000100011110010010011011;
    rom[6682] = 25'b0000100011110101011110100;
    rom[6683] = 25'b0000100011111000100110000;
    rom[6684] = 25'b0000100011111011101001101;
    rom[6685] = 25'b0000100011111110101001101;
    rom[6686] = 25'b0000100100000001100110000;
    rom[6687] = 25'b0000100100000100011110011;
    rom[6688] = 25'b0000100100000111010011001;
    rom[6689] = 25'b0000100100001010000011111;
    rom[6690] = 25'b0000100100001100110001000;
    rom[6691] = 25'b0000100100001111011010010;
    rom[6692] = 25'b0000100100010001111111101;
    rom[6693] = 25'b0000100100010100100001001;
    rom[6694] = 25'b0000100100010110111110111;
    rom[6695] = 25'b0000100100011001011000100;
    rom[6696] = 25'b0000100100011011101110011;
    rom[6697] = 25'b0000100100011110000000011;
    rom[6698] = 25'b0000100100100000001110011;
    rom[6699] = 25'b0000100100100010011000100;
    rom[6700] = 25'b0000100100100100011110100;
    rom[6701] = 25'b0000100100100110100000101;
    rom[6702] = 25'b0000100100101000011110111;
    rom[6703] = 25'b0000100100101010011001000;
    rom[6704] = 25'b0000100100101100001111001;
    rom[6705] = 25'b0000100100101110000001001;
    rom[6706] = 25'b0000100100101111101111010;
    rom[6707] = 25'b0000100100110001011001010;
    rom[6708] = 25'b0000100100110010111111010;
    rom[6709] = 25'b0000100100110100100001001;
    rom[6710] = 25'b0000100100110101111111000;
    rom[6711] = 25'b0000100100110111011000101;
    rom[6712] = 25'b0000100100111000101110010;
    rom[6713] = 25'b0000100100111001111111101;
    rom[6714] = 25'b0000100100111011001101000;
    rom[6715] = 25'b0000100100111100010110001;
    rom[6716] = 25'b0000100100111101011011001;
    rom[6717] = 25'b0000100100111110011100000;
    rom[6718] = 25'b0000100100111111011000100;
    rom[6719] = 25'b0000100101000000010001000;
    rom[6720] = 25'b0000100101000001000101010;
    rom[6721] = 25'b0000100101000001110101001;
    rom[6722] = 25'b0000100101000010100001000;
    rom[6723] = 25'b0000100101000011001000011;
    rom[6724] = 25'b0000100101000011101011110;
    rom[6725] = 25'b0000100101000100001010101;
    rom[6726] = 25'b0000100101000100100101011;
    rom[6727] = 25'b0000100101000100111011101;
    rom[6728] = 25'b0000100101000101001101111;
    rom[6729] = 25'b0000100101000101011011100;
    rom[6730] = 25'b0000100101000101100101000;
    rom[6731] = 25'b0000100101000101101010001;
    rom[6732] = 25'b0000100101000101101010111;
    rom[6733] = 25'b0000100101000101100111010;
    rom[6734] = 25'b0000100101000101011111010;
    rom[6735] = 25'b0000100101000101010010111;
    rom[6736] = 25'b0000100101000101000010001;
    rom[6737] = 25'b0000100101000100101101000;
    rom[6738] = 25'b0000100101000100010011100;
    rom[6739] = 25'b0000100101000011110101011;
    rom[6740] = 25'b0000100101000011010011000;
    rom[6741] = 25'b0000100101000010101100001;
    rom[6742] = 25'b0000100101000010000000111;
    rom[6743] = 25'b0000100101000001010001000;
    rom[6744] = 25'b0000100101000000011100110;
    rom[6745] = 25'b0000100100111111100100000;
    rom[6746] = 25'b0000100100111110100110110;
    rom[6747] = 25'b0000100100111101100101001;
    rom[6748] = 25'b0000100100111100011110111;
    rom[6749] = 25'b0000100100111011010100001;
    rom[6750] = 25'b0000100100111010000100110;
    rom[6751] = 25'b0000100100111000110001000;
    rom[6752] = 25'b0000100100110111011000100;
    rom[6753] = 25'b0000100100110101111011101;
    rom[6754] = 25'b0000100100110100011010001;
    rom[6755] = 25'b0000100100110010110100001;
    rom[6756] = 25'b0000100100110001001001100;
    rom[6757] = 25'b0000100100101111011010010;
    rom[6758] = 25'b0000100100101101100110100;
    rom[6759] = 25'b0000100100101011101110000;
    rom[6760] = 25'b0000100100101001110001000;
    rom[6761] = 25'b0000100100100111101111010;
    rom[6762] = 25'b0000100100100101101001000;
    rom[6763] = 25'b0000100100100011011110001;
    rom[6764] = 25'b0000100100100001001110101;
    rom[6765] = 25'b0000100100011110111010011;
    rom[6766] = 25'b0000100100011100100001100;
    rom[6767] = 25'b0000100100011010000011111;
    rom[6768] = 25'b0000100100010111100001110;
    rom[6769] = 25'b0000100100010100111010110;
    rom[6770] = 25'b0000100100010010001111010;
    rom[6771] = 25'b0000100100001111011111000;
    rom[6772] = 25'b0000100100001100101010000;
    rom[6773] = 25'b0000100100001001110000011;
    rom[6774] = 25'b0000100100000110110010000;
    rom[6775] = 25'b0000100100000011101110111;
    rom[6776] = 25'b0000100100000000100111000;
    rom[6777] = 25'b0000100011111101011010100;
    rom[6778] = 25'b0000100011111010001001010;
    rom[6779] = 25'b0000100011110110110011001;
    rom[6780] = 25'b0000100011110011011000011;
    rom[6781] = 25'b0000100011101111111000111;
    rom[6782] = 25'b0000100011101100010100100;
    rom[6783] = 25'b0000100011101000101011100;
    rom[6784] = 25'b0000100011100100111101101;
    rom[6785] = 25'b0000100011100001001011000;
    rom[6786] = 25'b0000100011011101010011101;
    rom[6787] = 25'b0000100011011001010111100;
    rom[6788] = 25'b0000100011010101010110100;
    rom[6789] = 25'b0000100011010001010000110;
    rom[6790] = 25'b0000100011001101000110010;
    rom[6791] = 25'b0000100011001000110111000;
    rom[6792] = 25'b0000100011000100100010110;
    rom[6793] = 25'b0000100011000000001001110;
    rom[6794] = 25'b0000100010111011101100000;
    rom[6795] = 25'b0000100010110111001001100;
    rom[6796] = 25'b0000100010110010100010000;
    rom[6797] = 25'b0000100010101101110101110;
    rom[6798] = 25'b0000100010101001000100101;
    rom[6799] = 25'b0000100010100100001110110;
    rom[6800] = 25'b0000100010011111010100001;
    rom[6801] = 25'b0000100010011010010100100;
    rom[6802] = 25'b0000100010010101010000000;
    rom[6803] = 25'b0000100010010000000110110;
    rom[6804] = 25'b0000100010001010111000101;
    rom[6805] = 25'b0000100010000101100101110;
    rom[6806] = 25'b0000100010000000001101111;
    rom[6807] = 25'b0000100001111010110001010;
    rom[6808] = 25'b0000100001110101001111110;
    rom[6809] = 25'b0000100001101111101001011;
    rom[6810] = 25'b0000100001101001111110001;
    rom[6811] = 25'b0000100001100100001110000;
    rom[6812] = 25'b0000100001011110011001001;
    rom[6813] = 25'b0000100001011000011111010;
    rom[6814] = 25'b0000100001010010100000100;
    rom[6815] = 25'b0000100001001100011100111;
    rom[6816] = 25'b0000100001000110010100100;
    rom[6817] = 25'b0000100001000000000111010;
    rom[6818] = 25'b0000100000111001110101000;
    rom[6819] = 25'b0000100000110011011110000;
    rom[6820] = 25'b0000100000101101000010001;
    rom[6821] = 25'b0000100000100110100001010;
    rom[6822] = 25'b0000100000011111111011101;
    rom[6823] = 25'b0000100000011001010001001;
    rom[6824] = 25'b0000100000010010100001110;
    rom[6825] = 25'b0000100000001011101101011;
    rom[6826] = 25'b0000100000000100110100010;
    rom[6827] = 25'b0000011111111101110110010;
    rom[6828] = 25'b0000011111110110110011011;
    rom[6829] = 25'b0000011111101111101011100;
    rom[6830] = 25'b0000011111101000011111000;
    rom[6831] = 25'b0000011111100001001101011;
    rom[6832] = 25'b0000011111011001110111000;
    rom[6833] = 25'b0000011111010010011011110;
    rom[6834] = 25'b0000011111001010111011101;
    rom[6835] = 25'b0000011111000011010110101;
    rom[6836] = 25'b0000011110111011101100111;
    rom[6837] = 25'b0000011110110011111110001;
    rom[6838] = 25'b0000011110101100001010100;
    rom[6839] = 25'b0000011110100100010010001;
    rom[6840] = 25'b0000011110011100010100111;
    rom[6841] = 25'b0000011110010100010010110;
    rom[6842] = 25'b0000011110001100001011110;
    rom[6843] = 25'b0000011110000011111111111;
    rom[6844] = 25'b0000011101111011101111010;
    rom[6845] = 25'b0000011101110011011001110;
    rom[6846] = 25'b0000011101101010111111011;
    rom[6847] = 25'b0000011101100010100000010;
    rom[6848] = 25'b0000011101011001111100001;
    rom[6849] = 25'b0000011101010001010011011;
    rom[6850] = 25'b0000011101001000100101101;
    rom[6851] = 25'b0000011100111111110011001;
    rom[6852] = 25'b0000011100110110111011111;
    rom[6853] = 25'b0000011100101101111111110;
    rom[6854] = 25'b0000011100100100111110110;
    rom[6855] = 25'b0000011100011011111001000;
    rom[6856] = 25'b0000011100010010101110100;
    rom[6857] = 25'b0000011100001001011111001;
    rom[6858] = 25'b0000011100000000001011000;
    rom[6859] = 25'b0000011011110110110010001;
    rom[6860] = 25'b0000011011101101010100011;
    rom[6861] = 25'b0000011011100011110001111;
    rom[6862] = 25'b0000011011011010001010101;
    rom[6863] = 25'b0000011011010000011110101;
    rom[6864] = 25'b0000011011000110101101111;
    rom[6865] = 25'b0000011010111100111000010;
    rom[6866] = 25'b0000011010110010111110000;
    rom[6867] = 25'b0000011010101000111111000;
    rom[6868] = 25'b0000011010011110111011001;
    rom[6869] = 25'b0000011010010100110010110;
    rom[6870] = 25'b0000011010001010100101011;
    rom[6871] = 25'b0000011010000000010011100;
    rom[6872] = 25'b0000011001110101111100111;
    rom[6873] = 25'b0000011001101011100001100;
    rom[6874] = 25'b0000011001100001000001100;
    rom[6875] = 25'b0000011001010110011100110;
    rom[6876] = 25'b0000011001001011110011010;
    rom[6877] = 25'b0000011001000001000101010;
    rom[6878] = 25'b0000011000110110010010011;
    rom[6879] = 25'b0000011000101011011011000;
    rom[6880] = 25'b0000011000100000011111000;
    rom[6881] = 25'b0000011000010101011110010;
    rom[6882] = 25'b0000011000001010011000111;
    rom[6883] = 25'b0000010111111111001110111;
    rom[6884] = 25'b0000010111110100000000010;
    rom[6885] = 25'b0000010111101000101101001;
    rom[6886] = 25'b0000010111011101010101010;
    rom[6887] = 25'b0000010111010001111000111;
    rom[6888] = 25'b0000010111000110010111111;
    rom[6889] = 25'b0000010110111010110010010;
    rom[6890] = 25'b0000010110101111001000010;
    rom[6891] = 25'b0000010110100011011001100;
    rom[6892] = 25'b0000010110010111100110010;
    rom[6893] = 25'b0000010110001011101110100;
    rom[6894] = 25'b0000010101111111110010010;
    rom[6895] = 25'b0000010101110011110001100;
    rom[6896] = 25'b0000010101100111101100001;
    rom[6897] = 25'b0000010101011011100010011;
    rom[6898] = 25'b0000010101001111010100001;
    rom[6899] = 25'b0000010101000011000001010;
    rom[6900] = 25'b0000010100110110101010001;
    rom[6901] = 25'b0000010100101010001110100;
    rom[6902] = 25'b0000010100011101101110011;
    rom[6903] = 25'b0000010100010001001001110;
    rom[6904] = 25'b0000010100000100100000111;
    rom[6905] = 25'b0000010011110111110011100;
    rom[6906] = 25'b0000010011101011000001110;
    rom[6907] = 25'b0000010011011110001011101;
    rom[6908] = 25'b0000010011010001010001001;
    rom[6909] = 25'b0000010011000100010010010;
    rom[6910] = 25'b0000010010110111001111001;
    rom[6911] = 25'b0000010010101010000111101;
    rom[6912] = 25'b0000010010011100111011110;
    rom[6913] = 25'b0000010010001111101011101;
    rom[6914] = 25'b0000010010000010010111001;
    rom[6915] = 25'b0000010001110100111110011;
    rom[6916] = 25'b0000010001100111100001011;
    rom[6917] = 25'b0000010001011010000000001;
    rom[6918] = 25'b0000010001001100011010110;
    rom[6919] = 25'b0000010000111110110000111;
    rom[6920] = 25'b0000010000110001000011000;
    rom[6921] = 25'b0000010000100011010000111;
    rom[6922] = 25'b0000010000010101011010101;
    rom[6923] = 25'b0000010000000111100000001;
    rom[6924] = 25'b0000001111111001100001100;
    rom[6925] = 25'b0000001111101011011110110;
    rom[6926] = 25'b0000001111011101010111111;
    rom[6927] = 25'b0000001111001111001100111;
    rom[6928] = 25'b0000001111000000111101110;
    rom[6929] = 25'b0000001110110010101010100;
    rom[6930] = 25'b0000001110100100010011010;
    rom[6931] = 25'b0000001110010101111000000;
    rom[6932] = 25'b0000001110000111011000110;
    rom[6933] = 25'b0000001101111000110101010;
    rom[6934] = 25'b0000001101101010001110000;
    rom[6935] = 25'b0000001101011011100010101;
    rom[6936] = 25'b0000001101001100110011011;
    rom[6937] = 25'b0000001100111110000000001;
    rom[6938] = 25'b0000001100101111001000111;
    rom[6939] = 25'b0000001100100000001101110;
    rom[6940] = 25'b0000001100010001001110110;
    rom[6941] = 25'b0000001100000010001011111;
    rom[6942] = 25'b0000001011110011000101001;
    rom[6943] = 25'b0000001011100011111010100;
    rom[6944] = 25'b0000001011010100101100000;
    rom[6945] = 25'b0000001011000101011001110;
    rom[6946] = 25'b0000001010110110000011101;
    rom[6947] = 25'b0000001010100110101001110;
    rom[6948] = 25'b0000001010010111001100010;
    rom[6949] = 25'b0000001010000111101010111;
    rom[6950] = 25'b0000001001111000000101110;
    rom[6951] = 25'b0000001001101000011101000;
    rom[6952] = 25'b0000001001011000110000100;
    rom[6953] = 25'b0000001001001001000000011;
    rom[6954] = 25'b0000001000111001001100101;
    rom[6955] = 25'b0000001000101001010101001;
    rom[6956] = 25'b0000001000011001011010001;
    rom[6957] = 25'b0000001000001001011011100;
    rom[6958] = 25'b0000000111111001011001010;
    rom[6959] = 25'b0000000111101001010011100;
    rom[6960] = 25'b0000000111011001001010001;
    rom[6961] = 25'b0000000111001000111101011;
    rom[6962] = 25'b0000000110111000101101000;
    rom[6963] = 25'b0000000110101000011001010;
    rom[6964] = 25'b0000000110011000000010000;
    rom[6965] = 25'b0000000110000111100111011;
    rom[6966] = 25'b0000000101110111001001010;
    rom[6967] = 25'b0000000101100110100111110;
    rom[6968] = 25'b0000000101010110000010111;
    rom[6969] = 25'b0000000101000101011010110;
    rom[6970] = 25'b0000000100110100101111010;
    rom[6971] = 25'b0000000100100100000000100;
    rom[6972] = 25'b0000000100010011001110010;
    rom[6973] = 25'b0000000100000010011000111;
    rom[6974] = 25'b0000000011110001100000011;
    rom[6975] = 25'b0000000011100000100100100;
    rom[6976] = 25'b0000000011001111100101100;
    rom[6977] = 25'b0000000010111110100011010;
    rom[6978] = 25'b0000000010101101011101111;
    rom[6979] = 25'b0000000010011100010101011;
    rom[6980] = 25'b0000000010001011001001111;
    rom[6981] = 25'b0000000001111001111011001;
    rom[6982] = 25'b0000000001101000101001011;
    rom[6983] = 25'b0000000001010111010100100;
    rom[6984] = 25'b0000000001000101111100110;
    rom[6985] = 25'b0000000000110100100010000;
    rom[6986] = 25'b0000000000100011000100010;
    rom[6987] = 25'b0000000000010001100011100;
    rom[6988] = 25'b0000000000000000000000000;
    rom[6989] = 25'b1111111111101110011001100;
    rom[6990] = 25'b1111111111011100110000001;
    rom[6991] = 25'b1111111111001011000011110;
    rom[6992] = 25'b1111111110111001010100110;
    rom[6993] = 25'b1111111110100111100010111;
    rom[6994] = 25'b1111111110010101101110001;
    rom[6995] = 25'b1111111110000011110110110;
    rom[6996] = 25'b1111111101110001111100101;
    rom[6997] = 25'b1111111101011111111111111;
    rom[6998] = 25'b1111111101001110000000011;
    rom[6999] = 25'b1111111100111011111110010;
    rom[7000] = 25'b1111111100101001111001100;
    rom[7001] = 25'b1111111100010111110010000;
    rom[7002] = 25'b1111111100000101101000001;
    rom[7003] = 25'b1111111011110011011011101;
    rom[7004] = 25'b1111111011100001001100101;
    rom[7005] = 25'b1111111011001110111011000;
    rom[7006] = 25'b1111111010111100100111001;
    rom[7007] = 25'b1111111010101010010000101;
    rom[7008] = 25'b1111111010010111110111110;
    rom[7009] = 25'b1111111010000101011100100;
    rom[7010] = 25'b1111111001110010111111000;
    rom[7011] = 25'b1111111001100000011111000;
    rom[7012] = 25'b1111111001001101111100110;
    rom[7013] = 25'b1111111000111011011000010;
    rom[7014] = 25'b1111111000101000110001100;
    rom[7015] = 25'b1111111000010110001000100;
    rom[7016] = 25'b1111111000000011011101010;
    rom[7017] = 25'b1111110111110000101111111;
    rom[7018] = 25'b1111110111011110000000011;
    rom[7019] = 25'b1111110111001011001110110;
    rom[7020] = 25'b1111110110111000011011000;
    rom[7021] = 25'b1111110110100101100101001;
    rom[7022] = 25'b1111110110010010101101011;
    rom[7023] = 25'b1111110101111111110011100;
    rom[7024] = 25'b1111110101101100110111101;
    rom[7025] = 25'b1111110101011001111001111;
    rom[7026] = 25'b1111110101000110111010010;
    rom[7027] = 25'b1111110100110011111000110;
    rom[7028] = 25'b1111110100100000110101010;
    rom[7029] = 25'b1111110100001101110000000;
    rom[7030] = 25'b1111110011111010101000111;
    rom[7031] = 25'b1111110011100111100000000;
    rom[7032] = 25'b1111110011010100010101100;
    rom[7033] = 25'b1111110011000001001001010;
    rom[7034] = 25'b1111110010101101111011010;
    rom[7035] = 25'b1111110010011010101011101;
    rom[7036] = 25'b1111110010000111011010011;
    rom[7037] = 25'b1111110001110100000111100;
    rom[7038] = 25'b1111110001100000110011010;
    rom[7039] = 25'b1111110001001101011101010;
    rom[7040] = 25'b1111110000111010000101110;
    rom[7041] = 25'b1111110000100110101100111;
    rom[7042] = 25'b1111110000010011010010100;
    rom[7043] = 25'b1111101111111111110110110;
    rom[7044] = 25'b1111101111101100011001101;
    rom[7045] = 25'b1111101111011000111011001;
    rom[7046] = 25'b1111101111000101011011010;
    rom[7047] = 25'b1111101110110001111010010;
    rom[7048] = 25'b1111101110011110010111111;
    rom[7049] = 25'b1111101110001010110100010;
    rom[7050] = 25'b1111101101110111001111100;
    rom[7051] = 25'b1111101101100011101001101;
    rom[7052] = 25'b1111101101010000000010100;
    rom[7053] = 25'b1111101100111100011010011;
    rom[7054] = 25'b1111101100101000110001001;
    rom[7055] = 25'b1111101100010101000110111;
    rom[7056] = 25'b1111101100000001011011110;
    rom[7057] = 25'b1111101011101101101111100;
    rom[7058] = 25'b1111101011011010000010010;
    rom[7059] = 25'b1111101011000110010100010;
    rom[7060] = 25'b1111101010110010100101011;
    rom[7061] = 25'b1111101010011110110101100;
    rom[7062] = 25'b1111101010001011000101001;
    rom[7063] = 25'b1111101001110111010011110;
    rom[7064] = 25'b1111101001100011100001101;
    rom[7065] = 25'b1111101001001111101110111;
    rom[7066] = 25'b1111101000111011111011011;
    rom[7067] = 25'b1111101000101000000111010;
    rom[7068] = 25'b1111101000010100010010101;
    rom[7069] = 25'b1111101000000000011101011;
    rom[7070] = 25'b1111100111101100100111101;
    rom[7071] = 25'b1111100111011000110001010;
    rom[7072] = 25'b1111100111000100111010100;
    rom[7073] = 25'b1111100110110001000011010;
    rom[7074] = 25'b1111100110011101001011101;
    rom[7075] = 25'b1111100110001001010011110;
    rom[7076] = 25'b1111100101110101011011011;
    rom[7077] = 25'b1111100101100001100010111;
    rom[7078] = 25'b1111100101001101101010000;
    rom[7079] = 25'b1111100100111001110000111;
    rom[7080] = 25'b1111100100100101110111101;
    rom[7081] = 25'b1111100100010001111110000;
    rom[7082] = 25'b1111100011111110000100100;
    rom[7083] = 25'b1111100011101010001010111;
    rom[7084] = 25'b1111100011010110010001001;
    rom[7085] = 25'b1111100011000010010111011;
    rom[7086] = 25'b1111100010101110011101101;
    rom[7087] = 25'b1111100010011010100011111;
    rom[7088] = 25'b1111100010000110101010011;
    rom[7089] = 25'b1111100001110010110000111;
    rom[7090] = 25'b1111100001011110110111101;
    rom[7091] = 25'b1111100001001010111110100;
    rom[7092] = 25'b1111100000110111000101101;
    rom[7093] = 25'b1111100000100011001101000;
    rom[7094] = 25'b1111100000001111010100101;
    rom[7095] = 25'b1111011111111011011100101;
    rom[7096] = 25'b1111011111100111100101000;
    rom[7097] = 25'b1111011111010011101101110;
    rom[7098] = 25'b1111011110111111110111000;
    rom[7099] = 25'b1111011110101100000000110;
    rom[7100] = 25'b1111011110011000001010111;
    rom[7101] = 25'b1111011110000100010101101;
    rom[7102] = 25'b1111011101110000100001000;
    rom[7103] = 25'b1111011101011100101101000;
    rom[7104] = 25'b1111011101001000111001110;
    rom[7105] = 25'b1111011100110101000111001;
    rom[7106] = 25'b1111011100100001010101010;
    rom[7107] = 25'b1111011100001101100100000;
    rom[7108] = 25'b1111011011111001110011110;
    rom[7109] = 25'b1111011011100110000100010;
    rom[7110] = 25'b1111011011010010010101101;
    rom[7111] = 25'b1111011010111110101000000;
    rom[7112] = 25'b1111011010101010111011010;
    rom[7113] = 25'b1111011010010111001111101;
    rom[7114] = 25'b1111011010000011100101000;
    rom[7115] = 25'b1111011001101111111011010;
    rom[7116] = 25'b1111011001011100010010111;
    rom[7117] = 25'b1111011001001000101011100;
    rom[7118] = 25'b1111011000110101000101010;
    rom[7119] = 25'b1111011000100001100000011;
    rom[7120] = 25'b1111011000001101111100110;
    rom[7121] = 25'b1111010111111010011010011;
    rom[7122] = 25'b1111010111100110111001010;
    rom[7123] = 25'b1111010111010011011001101;
    rom[7124] = 25'b1111010110111111111011011;
    rom[7125] = 25'b1111010110101100011110101;
    rom[7126] = 25'b1111010110011001000011010;
    rom[7127] = 25'b1111010110000101101001100;
    rom[7128] = 25'b1111010101110010010001010;
    rom[7129] = 25'b1111010101011110111010101;
    rom[7130] = 25'b1111010101001011100101101;
    rom[7131] = 25'b1111010100111000010010011;
    rom[7132] = 25'b1111010100100101000000110;
    rom[7133] = 25'b1111010100010001110000111;
    rom[7134] = 25'b1111010011111110100010111;
    rom[7135] = 25'b1111010011101011010110101;
    rom[7136] = 25'b1111010011011000001100011;
    rom[7137] = 25'b1111010011000101000011111;
    rom[7138] = 25'b1111010010110001111101100;
    rom[7139] = 25'b1111010010011110111001000;
    rom[7140] = 25'b1111010010001011110110100;
    rom[7141] = 25'b1111010001111000110110010;
    rom[7142] = 25'b1111010001100101110111111;
    rom[7143] = 25'b1111010001010010111011111;
    rom[7144] = 25'b1111010001000000000001111;
    rom[7145] = 25'b1111010000101101001010001;
    rom[7146] = 25'b1111010000011010010100110;
    rom[7147] = 25'b1111010000000111100001101;
    rom[7148] = 25'b1111001111110100110000101;
    rom[7149] = 25'b1111001111100010000010011;
    rom[7150] = 25'b1111001111001111010110011;
    rom[7151] = 25'b1111001110111100101100110;
    rom[7152] = 25'b1111001110101010000101110;
    rom[7153] = 25'b1111001110010111100001001;
    rom[7154] = 25'b1111001110000100111111010;
    rom[7155] = 25'b1111001101110010011111111;
    rom[7156] = 25'b1111001101100000000011010;
    rom[7157] = 25'b1111001101001101101001011;
    rom[7158] = 25'b1111001100111011010010001;
    rom[7159] = 25'b1111001100101000111101101;
    rom[7160] = 25'b1111001100010110101100000;
    rom[7161] = 25'b1111001100000100011101010;
    rom[7162] = 25'b1111001011110010010001011;
    rom[7163] = 25'b1111001011100000001000011;
    rom[7164] = 25'b1111001011001110000010011;
    rom[7165] = 25'b1111001010111011111111100;
    rom[7166] = 25'b1111001010101001111111100;
    rom[7167] = 25'b1111001010011000000010101;
    rom[7168] = 25'b1111001010000110001001000;
    rom[7169] = 25'b1111001001110100010010100;
    rom[7170] = 25'b1111001001100010011111010;
    rom[7171] = 25'b1111001001010000101111010;
    rom[7172] = 25'b1111001000111111000010100;
    rom[7173] = 25'b1111001000101101011001000;
    rom[7174] = 25'b1111001000011011110010111;
    rom[7175] = 25'b1111001000001010010000011;
    rom[7176] = 25'b1111000111111000110001001;
    rom[7177] = 25'b1111000111100111010101100;
    rom[7178] = 25'b1111000111010101111101011;
    rom[7179] = 25'b1111000111000100101000110;
    rom[7180] = 25'b1111000110110011010111111;
    rom[7181] = 25'b1111000110100010001010100;
    rom[7182] = 25'b1111000110010001000000111;
    rom[7183] = 25'b1111000101111111111011000;
    rom[7184] = 25'b1111000101101110111000111;
    rom[7185] = 25'b1111000101011101111010101;
    rom[7186] = 25'b1111000101001101000000010;
    rom[7187] = 25'b1111000100111100001001101;
    rom[7188] = 25'b1111000100101011010111001;
    rom[7189] = 25'b1111000100011010101000011;
    rom[7190] = 25'b1111000100001001111101110;
    rom[7191] = 25'b1111000011111001010111010;
    rom[7192] = 25'b1111000011101000110100111;
    rom[7193] = 25'b1111000011011000010110100;
    rom[7194] = 25'b1111000011000111111100010;
    rom[7195] = 25'b1111000010110111100110011;
    rom[7196] = 25'b1111000010100111010100110;
    rom[7197] = 25'b1111000010010111000111011;
    rom[7198] = 25'b1111000010000110111110010;
    rom[7199] = 25'b1111000001110110111001101;
    rom[7200] = 25'b1111000001100110111001011;
    rom[7201] = 25'b1111000001010110111101101;
    rom[7202] = 25'b1111000001000111000110010;
    rom[7203] = 25'b1111000000110111010011100;
    rom[7204] = 25'b1111000000100111100101011;
    rom[7205] = 25'b1111000000010111111011110;
    rom[7206] = 25'b1111000000001000010110111;
    rom[7207] = 25'b1110111111111000110110101;
    rom[7208] = 25'b1110111111101001011011001;
    rom[7209] = 25'b1110111111011010000100100;
    rom[7210] = 25'b1110111111001010110010101;
    rom[7211] = 25'b1110111110111011100101100;
    rom[7212] = 25'b1110111110101100011101100;
    rom[7213] = 25'b1110111110011101011010010;
    rom[7214] = 25'b1110111110001110011100001;
    rom[7215] = 25'b1110111101111111100010111;
    rom[7216] = 25'b1110111101110000101110101;
    rom[7217] = 25'b1110111101100001111111110;
    rom[7218] = 25'b1110111101010011010101110;
    rom[7219] = 25'b1110111101000100110001000;
    rom[7220] = 25'b1110111100110110010001100;
    rom[7221] = 25'b1110111100100111110111010;
    rom[7222] = 25'b1110111100011001100010011;
    rom[7223] = 25'b1110111100001011010010110;
    rom[7224] = 25'b1110111011111101001000011;
    rom[7225] = 25'b1110111011101111000011101;
    rom[7226] = 25'b1110111011100001000100010;
    rom[7227] = 25'b1110111011010011001010011;
    rom[7228] = 25'b1110111011000101010110000;
    rom[7229] = 25'b1110111010110111100111010;
    rom[7230] = 25'b1110111010101001111110000;
    rom[7231] = 25'b1110111010011100011010100;
    rom[7232] = 25'b1110111010001110111100110;
    rom[7233] = 25'b1110111010000001100100101;
    rom[7234] = 25'b1110111001110100010010010;
    rom[7235] = 25'b1110111001100111000101110;
    rom[7236] = 25'b1110111001011001111111001;
    rom[7237] = 25'b1110111001001100111110011;
    rom[7238] = 25'b1110111001000000000011011;
    rom[7239] = 25'b1110111000110011001110100;
    rom[7240] = 25'b1110111000100110011111101;
    rom[7241] = 25'b1110111000011001110110110;
    rom[7242] = 25'b1110111000001101010100000;
    rom[7243] = 25'b1110111000000000110111011;
    rom[7244] = 25'b1110110111110100100000111;
    rom[7245] = 25'b1110110111101000010000101;
    rom[7246] = 25'b1110110111011100000110101;
    rom[7247] = 25'b1110110111010000000010110;
    rom[7248] = 25'b1110110111000100000101011;
    rom[7249] = 25'b1110110110111000001110010;
    rom[7250] = 25'b1110110110101100011101101;
    rom[7251] = 25'b1110110110100000110011010;
    rom[7252] = 25'b1110110110010101001111100;
    rom[7253] = 25'b1110110110001001110010001;
    rom[7254] = 25'b1110110101111110011011011;
    rom[7255] = 25'b1110110101110011001011001;
    rom[7256] = 25'b1110110101101000000001101;
    rom[7257] = 25'b1110110101011100111110110;
    rom[7258] = 25'b1110110101010010000010101;
    rom[7259] = 25'b1110110101000111001101001;
    rom[7260] = 25'b1110110100111100011110011;
    rom[7261] = 25'b1110110100110001110110101;
    rom[7262] = 25'b1110110100100111010101100;
    rom[7263] = 25'b1110110100011100111011011;
    rom[7264] = 25'b1110110100010010101000001;
    rom[7265] = 25'b1110110100001000011011111;
    rom[7266] = 25'b1110110011111110010110101;
    rom[7267] = 25'b1110110011110100011000011;
    rom[7268] = 25'b1110110011101010100001010;
    rom[7269] = 25'b1110110011100000110001010;
    rom[7270] = 25'b1110110011010111001000011;
    rom[7271] = 25'b1110110011001101100110101;
    rom[7272] = 25'b1110110011000100001100001;
    rom[7273] = 25'b1110110010111010111000111;
    rom[7274] = 25'b1110110010110001101101000;
    rom[7275] = 25'b1110110010101000101000011;
    rom[7276] = 25'b1110110010011111101011010;
    rom[7277] = 25'b1110110010010110110101011;
    rom[7278] = 25'b1110110010001110000111000;
    rom[7279] = 25'b1110110010000101100000001;
    rom[7280] = 25'b1110110001111101000000101;
    rom[7281] = 25'b1110110001110100101000111;
    rom[7282] = 25'b1110110001101100011000110;
    rom[7283] = 25'b1110110001100100010000000;
    rom[7284] = 25'b1110110001011100001111000;
    rom[7285] = 25'b1110110001010100010101111;
    rom[7286] = 25'b1110110001001100100100010;
    rom[7287] = 25'b1110110001000100111010100;
    rom[7288] = 25'b1110110000111101011000101;
    rom[7289] = 25'b1110110000110101111110011;
    rom[7290] = 25'b1110110000101110101100001;
    rom[7291] = 25'b1110110000100111100001111;
    rom[7292] = 25'b1110110000100000011111011;
    rom[7293] = 25'b1110110000011001100101000;
    rom[7294] = 25'b1110110000010010110010101;
    rom[7295] = 25'b1110110000001100001000010;
    rom[7296] = 25'b1110110000000101100110000;
    rom[7297] = 25'b1110101111111111001011111;
    rom[7298] = 25'b1110101111111000111001111;
    rom[7299] = 25'b1110101111110010110000000;
    rom[7300] = 25'b1110101111101100101110011;
    rom[7301] = 25'b1110101111100110110101001;
    rom[7302] = 25'b1110101111100001000100001;
    rom[7303] = 25'b1110101111011011011011011;
    rom[7304] = 25'b1110101111010101111010111;
    rom[7305] = 25'b1110101111010000100011000;
    rom[7306] = 25'b1110101111001011010011100;
    rom[7307] = 25'b1110101111000110001100011;
    rom[7308] = 25'b1110101111000001001101110;
    rom[7309] = 25'b1110101110111100010111110;
    rom[7310] = 25'b1110101110110111101010001;
    rom[7311] = 25'b1110101110110011000101010;
    rom[7312] = 25'b1110101110101110101001000;
    rom[7313] = 25'b1110101110101010010101011;
    rom[7314] = 25'b1110101110100110001010100;
    rom[7315] = 25'b1110101110100010001000010;
    rom[7316] = 25'b1110101110011110001110110;
    rom[7317] = 25'b1110101110011010011110001;
    rom[7318] = 25'b1110101110010110110110010;
    rom[7319] = 25'b1110101110010011010111010;
    rom[7320] = 25'b1110101110010000000001001;
    rom[7321] = 25'b1110101110001100110011111;
    rom[7322] = 25'b1110101110001001101111101;
    rom[7323] = 25'b1110101110000110110100100;
    rom[7324] = 25'b1110101110000100000010001;
    rom[7325] = 25'b1110101110000001011001000;
    rom[7326] = 25'b1110101101111110111000111;
    rom[7327] = 25'b1110101101111100100001111;
    rom[7328] = 25'b1110101101111010010011111;
    rom[7329] = 25'b1110101101111000001111010;
    rom[7330] = 25'b1110101101110110010011110;
    rom[7331] = 25'b1110101101110100100001011;
    rom[7332] = 25'b1110101101110010111000011;
    rom[7333] = 25'b1110101101110001011000110;
    rom[7334] = 25'b1110101101110000000010010;
    rom[7335] = 25'b1110101101101110110101010;
    rom[7336] = 25'b1110101101101101110001100;
    rom[7337] = 25'b1110101101101100110111010;
    rom[7338] = 25'b1110101101101100000110011;
    rom[7339] = 25'b1110101101101011011111000;
    rom[7340] = 25'b1110101101101011000001001;
    rom[7341] = 25'b1110101101101010101100110;
    rom[7342] = 25'b1110101101101010100010000;
    rom[7343] = 25'b1110101101101010100000110;
    rom[7344] = 25'b1110101101101010101001001;
    rom[7345] = 25'b1110101101101010111011010;
    rom[7346] = 25'b1110101101101011010111000;
    rom[7347] = 25'b1110101101101011111100011;
    rom[7348] = 25'b1110101101101100101011101;
    rom[7349] = 25'b1110101101101101100100100;
    rom[7350] = 25'b1110101101101110100111010;
    rom[7351] = 25'b1110101101101111110011110;
    rom[7352] = 25'b1110101101110001001010000;
    rom[7353] = 25'b1110101101110010101010010;
    rom[7354] = 25'b1110101101110100010100011;
    rom[7355] = 25'b1110101101110110001000011;
    rom[7356] = 25'b1110101101111000000110011;
    rom[7357] = 25'b1110101101111010001110011;
    rom[7358] = 25'b1110101101111100100000010;
    rom[7359] = 25'b1110101101111110111100010;
    rom[7360] = 25'b1110101110000001100010010;
    rom[7361] = 25'b1110101110000100010010011;
    rom[7362] = 25'b1110101110000111001100101;
    rom[7363] = 25'b1110101110001010010000111;
    rom[7364] = 25'b1110101110001101011111100;
    rom[7365] = 25'b1110101110010000111000001;
    rom[7366] = 25'b1110101110010100011011000;
    rom[7367] = 25'b1110101110011000001000010;
    rom[7368] = 25'b1110101110011011111111100;
    rom[7369] = 25'b1110101110100000000001010;
    rom[7370] = 25'b1110101110100100001101010;
    rom[7371] = 25'b1110101110101000100011100;
    rom[7372] = 25'b1110101110101101000100001;
    rom[7373] = 25'b1110101110110001101111010;
    rom[7374] = 25'b1110101110110110100100101;
    rom[7375] = 25'b1110101110111011100100100;
    rom[7376] = 25'b1110101111000000101110110;
    rom[7377] = 25'b1110101111000110000011101;
    rom[7378] = 25'b1110101111001011100010111;
    rom[7379] = 25'b1110101111010001001100101;
    rom[7380] = 25'b1110101111010111000001001;
    rom[7381] = 25'b1110101111011101000000000;
    rom[7382] = 25'b1110101111100011001001100;
    rom[7383] = 25'b1110101111101001011101101;
    rom[7384] = 25'b1110101111101111111100011;
    rom[7385] = 25'b1110101111110110100101110;
    rom[7386] = 25'b1110101111111101011001111;
    rom[7387] = 25'b1110110000000100011000101;
    rom[7388] = 25'b1110110000001011100010001;
    rom[7389] = 25'b1110110000010010110110011;
    rom[7390] = 25'b1110110000011010010101011;
    rom[7391] = 25'b1110110000100001111111001;
    rom[7392] = 25'b1110110000101001110011110;
    rom[7393] = 25'b1110110000110001110011001;
    rom[7394] = 25'b1110110000111001111101011;
    rom[7395] = 25'b1110110001000010010010100;
    rom[7396] = 25'b1110110001001010110010100;
    rom[7397] = 25'b1110110001010011011101100;
    rom[7398] = 25'b1110110001011100010011010;
    rom[7399] = 25'b1110110001100101010100000;
    rom[7400] = 25'b1110110001101110011111111;
    rom[7401] = 25'b1110110001110111110110100;
    rom[7402] = 25'b1110110010000001011000001;
    rom[7403] = 25'b1110110010001011000100111;
    rom[7404] = 25'b1110110010010100111100110;
    rom[7405] = 25'b1110110010011110111111100;
    rom[7406] = 25'b1110110010101001001101011;
    rom[7407] = 25'b1110110010110011100110011;
    rom[7408] = 25'b1110110010111110001010100;
    rom[7409] = 25'b1110110011001000111001101;
    rom[7410] = 25'b1110110011010011110100000;
    rom[7411] = 25'b1110110011011110111001100;
    rom[7412] = 25'b1110110011101010001010010;
    rom[7413] = 25'b1110110011110101100110001;
    rom[7414] = 25'b1110110100000001001101010;
    rom[7415] = 25'b1110110100001100111111100;
    rom[7416] = 25'b1110110100011000111101000;
    rom[7417] = 25'b1110110100100101000101111;
    rom[7418] = 25'b1110110100110001011010000;
    rom[7419] = 25'b1110110100111101111001011;
    rom[7420] = 25'b1110110101001010100100000;
    rom[7421] = 25'b1110110101010111011010000;
    rom[7422] = 25'b1110110101100100011011010;
    rom[7423] = 25'b1110110101110001100111111;
    rom[7424] = 25'b1110110101111110111111111;
    rom[7425] = 25'b1110110110001100100011011;
    rom[7426] = 25'b1110110110011010010010001;
    rom[7427] = 25'b1110110110101000001100010;
    rom[7428] = 25'b1110110110110110010001111;
    rom[7429] = 25'b1110110111000100100010111;
    rom[7430] = 25'b1110110111010010111111011;
    rom[7431] = 25'b1110110111100001100111010;
    rom[7432] = 25'b1110110111110000011010110;
    rom[7433] = 25'b1110110111111111011001100;
    rom[7434] = 25'b1110111000001110100011111;
    rom[7435] = 25'b1110111000011101111001110;
    rom[7436] = 25'b1110111000101101011011001;
    rom[7437] = 25'b1110111000111101001000000;
    rom[7438] = 25'b1110111001001101000000100;
    rom[7439] = 25'b1110111001011101000100011;
    rom[7440] = 25'b1110111001101101010011111;
    rom[7441] = 25'b1110111001111101101111000;
    rom[7442] = 25'b1110111010001110010101110;
    rom[7443] = 25'b1110111010011111001000000;
    rom[7444] = 25'b1110111010110000000101111;
    rom[7445] = 25'b1110111011000001001111011;
    rom[7446] = 25'b1110111011010010100100100;
    rom[7447] = 25'b1110111011100100000101010;
    rom[7448] = 25'b1110111011110101110001100;
    rom[7449] = 25'b1110111100000111101001101;
    rom[7450] = 25'b1110111100011001101101010;
    rom[7451] = 25'b1110111100101011111100101;
    rom[7452] = 25'b1110111100111110010111101;
    rom[7453] = 25'b1110111101010000111110011;
    rom[7454] = 25'b1110111101100011110000110;
    rom[7455] = 25'b1110111101110110101110101;
    rom[7456] = 25'b1110111110001001111000100;
    rom[7457] = 25'b1110111110011101001110000;
    rom[7458] = 25'b1110111110110000101111001;
    rom[7459] = 25'b1110111111000100011100001;
    rom[7460] = 25'b1110111111011000010100110;
    rom[7461] = 25'b1110111111101100011001001;
    rom[7462] = 25'b1111000000000000101001001;
    rom[7463] = 25'b1111000000010101000101000;
    rom[7464] = 25'b1111000000101001101100101;
    rom[7465] = 25'b1111000000111110100000000;
    rom[7466] = 25'b1111000001010011011111001;
    rom[7467] = 25'b1111000001101000101010000;
    rom[7468] = 25'b1111000001111110000000101;
    rom[7469] = 25'b1111000010010011100011001;
    rom[7470] = 25'b1111000010101001010001011;
    rom[7471] = 25'b1111000010111111001011010;
    rom[7472] = 25'b1111000011010101010001001;
    rom[7473] = 25'b1111000011101011100010101;
    rom[7474] = 25'b1111000100000010000000000;
    rom[7475] = 25'b1111000100011000101001001;
    rom[7476] = 25'b1111000100101111011110001;
    rom[7477] = 25'b1111000101000110011110111;
    rom[7478] = 25'b1111000101011101101011011;
    rom[7479] = 25'b1111000101110101000011110;
    rom[7480] = 25'b1111000110001100100111111;
    rom[7481] = 25'b1111000110100100010111111;
    rom[7482] = 25'b1111000110111100010011101;
    rom[7483] = 25'b1111000111010100011011010;
    rom[7484] = 25'b1111000111101100101110101;
    rom[7485] = 25'b1111001000000101001101111;
    rom[7486] = 25'b1111001000011101111000111;
    rom[7487] = 25'b1111001000110110101111101;
    rom[7488] = 25'b1111001001001111110010010;
    rom[7489] = 25'b1111001001101001000000110;
    rom[7490] = 25'b1111001010000010011010111;
    rom[7491] = 25'b1111001010011100000001000;
    rom[7492] = 25'b1111001010110101110010111;
    rom[7493] = 25'b1111001011001111110000100;
    rom[7494] = 25'b1111001011101001111010000;
    rom[7495] = 25'b1111001100000100001111010;
    rom[7496] = 25'b1111001100011110110000010;
    rom[7497] = 25'b1111001100111001011101001;
    rom[7498] = 25'b1111001101010100010101110;
    rom[7499] = 25'b1111001101101111011010010;
    rom[7500] = 25'b1111001110001010101010011;
    rom[7501] = 25'b1111001110100110000110100;
    rom[7502] = 25'b1111001111000001101110010;
    rom[7503] = 25'b1111001111011101100001110;
    rom[7504] = 25'b1111001111111001100001001;
    rom[7505] = 25'b1111010000010101101100010;
    rom[7506] = 25'b1111010000110010000011001;
    rom[7507] = 25'b1111010001001110100101110;
    rom[7508] = 25'b1111010001101011010100001;
    rom[7509] = 25'b1111010010001000001110001;
    rom[7510] = 25'b1111010010100101010100001;
    rom[7511] = 25'b1111010011000010100101101;
    rom[7512] = 25'b1111010011100000000011000;
    rom[7513] = 25'b1111010011111101101100000;
    rom[7514] = 25'b1111010100011011100000110;
    rom[7515] = 25'b1111010100111001100001001;
    rom[7516] = 25'b1111010101010111101101011;
    rom[7517] = 25'b1111010101110110000101010;
    rom[7518] = 25'b1111010110010100101000110;
    rom[7519] = 25'b1111010110110011011000000;
    rom[7520] = 25'b1111010111010010010010111;
    rom[7521] = 25'b1111010111110001011001100;
    rom[7522] = 25'b1111011000010000101011101;
    rom[7523] = 25'b1111011000110000001001100;
    rom[7524] = 25'b1111011001001111110011000;
    rom[7525] = 25'b1111011001101111101000001;
    rom[7526] = 25'b1111011010001111101000111;
    rom[7527] = 25'b1111011010101111110101010;
    rom[7528] = 25'b1111011011010000001101001;
    rom[7529] = 25'b1111011011110000110000101;
    rom[7530] = 25'b1111011100010001011111110;
    rom[7531] = 25'b1111011100110010011010100;
    rom[7532] = 25'b1111011101010011100000101;
    rom[7533] = 25'b1111011101110100110010011;
    rom[7534] = 25'b1111011110010110001111110;
    rom[7535] = 25'b1111011110110111111000011;
    rom[7536] = 25'b1111011111011001101100110;
    rom[7537] = 25'b1111011111111011101100101;
    rom[7538] = 25'b1111100000011101110111111;
    rom[7539] = 25'b1111100001000000001110101;
    rom[7540] = 25'b1111100001100010110000111;
    rom[7541] = 25'b1111100010000101011110100;
    rom[7542] = 25'b1111100010101000010111101;
    rom[7543] = 25'b1111100011001011011100000;
    rom[7544] = 25'b1111100011101110101011111;
    rom[7545] = 25'b1111100100010010000111010;
    rom[7546] = 25'b1111100100110101101101110;
    rom[7547] = 25'b1111100101011001011111111;
    rom[7548] = 25'b1111100101111101011101010;
    rom[7549] = 25'b1111100110100001100101111;
    rom[7550] = 25'b1111100111000101111001110;
    rom[7551] = 25'b1111100111101010011001000;
    rom[7552] = 25'b1111101000001111000011101;
    rom[7553] = 25'b1111101000110011111001100;
    rom[7554] = 25'b1111101001011000111010011;
    rom[7555] = 25'b1111101001111110000110110;
    rom[7556] = 25'b1111101010100011011110010;
    rom[7557] = 25'b1111101011001001000000111;
    rom[7558] = 25'b1111101011101110101110110;
    rom[7559] = 25'b1111101100010100100111111;
    rom[7560] = 25'b1111101100111010101100000;
    rom[7561] = 25'b1111101101100000111011010;
    rom[7562] = 25'b1111101110000111010101101;
    rom[7563] = 25'b1111101110101101111011001;
    rom[7564] = 25'b1111101111010100101011100;
    rom[7565] = 25'b1111101111111011100111001;
    rom[7566] = 25'b1111110000100010101101110;
    rom[7567] = 25'b1111110001001001111111011;
    rom[7568] = 25'b1111110001110001011011111;
    rom[7569] = 25'b1111110010011001000011100;
    rom[7570] = 25'b1111110011000000110110000;
    rom[7571] = 25'b1111110011101000110011011;
    rom[7572] = 25'b1111110100010000111011110;
    rom[7573] = 25'b1111110100111001001111000;
    rom[7574] = 25'b1111110101100001101100111;
    rom[7575] = 25'b1111110110001010010101111;
    rom[7576] = 25'b1111110110110011001001100;
    rom[7577] = 25'b1111110111011100001000000;
    rom[7578] = 25'b1111111000000101010001010;
    rom[7579] = 25'b1111111000101110100101011;
    rom[7580] = 25'b1111111001011000000100001;
    rom[7581] = 25'b1111111010000001101101100;
    rom[7582] = 25'b1111111010101011100001101;
    rom[7583] = 25'b1111111011010101100000011;
    rom[7584] = 25'b1111111011111111101001111;
    rom[7585] = 25'b1111111100101001111101111;
    rom[7586] = 25'b1111111101010100011100011;
    rom[7587] = 25'b1111111101111111000101100;
    rom[7588] = 25'b1111111110101001111001001;
    rom[7589] = 25'b1111111111010100110111011;
    rom[7590] = 25'b0000000000000000000000000;
    rom[7591] = 25'b0000000000101011010011000;
    rom[7592] = 25'b0000000001010110110000100;
    rom[7593] = 25'b0000000010000010011000100;
    rom[7594] = 25'b0000000010101110001010110;
    rom[7595] = 25'b0000000011011010000111011;
    rom[7596] = 25'b0000000100000110001110011;
    rom[7597] = 25'b0000000100110010011111101;
    rom[7598] = 25'b0000000101011110111011001;
    rom[7599] = 25'b0000000110001011100001000;
    rom[7600] = 25'b0000000110111000010001000;
    rom[7601] = 25'b0000000111100101001011001;
    rom[7602] = 25'b0000001000010010001111100;
    rom[7603] = 25'b0000001000111111011101110;
    rom[7604] = 25'b0000001001101100110110011;
    rom[7605] = 25'b0000001010011010011001000;
    rom[7606] = 25'b0000001011001000000101100;
    rom[7607] = 25'b0000001011110101111100010;
    rom[7608] = 25'b0000001100100011111100111;
    rom[7609] = 25'b0000001101010010000111100;
    rom[7610] = 25'b0000001110000000011011111;
    rom[7611] = 25'b0000001110101110111010010;
    rom[7612] = 25'b0000001111011101100010100;
    rom[7613] = 25'b0000010000001100010100100;
    rom[7614] = 25'b0000010000111011010000011;
    rom[7615] = 25'b0000010001101010010110000;
    rom[7616] = 25'b0000010010011001100101011;
    rom[7617] = 25'b0000010011001000111110011;
    rom[7618] = 25'b0000010011111000100001000;
    rom[7619] = 25'b0000010100101000001101010;
    rom[7620] = 25'b0000010101011000000011011;
    rom[7621] = 25'b0000010110001000000010110;
    rom[7622] = 25'b0000010110111000001011111;
    rom[7623] = 25'b0000010111101000011110011;
    rom[7624] = 25'b0000011000011000111010010;
    rom[7625] = 25'b0000011001001001011111110;
    rom[7626] = 25'b0000011001111010001110100;
    rom[7627] = 25'b0000011010101011000110110;
    rom[7628] = 25'b0000011011011100001000010;
    rom[7629] = 25'b0000011100001101010011000;
    rom[7630] = 25'b0000011100111110100111000;
    rom[7631] = 25'b0000011101110000000100011;
    rom[7632] = 25'b0000011110100001101010111;
    rom[7633] = 25'b0000011111010011011010100;
    rom[7634] = 25'b0000100000000101010011001;
    rom[7635] = 25'b0000100000110111010101000;
    rom[7636] = 25'b0000100001101001011111111;
    rom[7637] = 25'b0000100010011011110011101;
    rom[7638] = 25'b0000100011001110010000101;
    rom[7639] = 25'b0000100100000000110110011;
    rom[7640] = 25'b0000100100110011100101000;
    rom[7641] = 25'b0000100101100110011100100;
    rom[7642] = 25'b0000100110011001011100111;
    rom[7643] = 25'b0000100111001100100110000;
    rom[7644] = 25'b0000100111111111110111111;
    rom[7645] = 25'b0000101000110011010010100;
    rom[7646] = 25'b0000101001100110110101101;
    rom[7647] = 25'b0000101010011010100001101;
    rom[7648] = 25'b0000101011001110010110000;
    rom[7649] = 25'b0000101100000010010011000;
    rom[7650] = 25'b0000101100110110011000100;
    rom[7651] = 25'b0000101101101010100110101;
    rom[7652] = 25'b0000101110011110111100111;
    rom[7653] = 25'b0000101111010011011011110;
    rom[7654] = 25'b0000110000001000000011000;
    rom[7655] = 25'b0000110000111100110010011;
    rom[7656] = 25'b0000110001110001101010001;
    rom[7657] = 25'b0000110010100110101010001;
    rom[7658] = 25'b0000110011011011110010010;
    rom[7659] = 25'b0000110100010001000010100;
    rom[7660] = 25'b0000110101000110011010111;
    rom[7661] = 25'b0000110101111011111011011;
    rom[7662] = 25'b0000110110110001100011110;
    rom[7663] = 25'b0000110111100111010100010;
    rom[7664] = 25'b0000111000011101001100101;
    rom[7665] = 25'b0000111001010011001101000;
    rom[7666] = 25'b0000111010001001010101000;
    rom[7667] = 25'b0000111010111111100101000;
    rom[7668] = 25'b0000111011110101111100101;
    rom[7669] = 25'b0000111100101100011100000;
    rom[7670] = 25'b0000111101100011000011001;
    rom[7671] = 25'b0000111110011001110001111;
    rom[7672] = 25'b0000111111010000101000001;
    rom[7673] = 25'b0001000000000111100101111;
    rom[7674] = 25'b0001000000111110101011011;
    rom[7675] = 25'b0001000001110101111000001;
    rom[7676] = 25'b0001000010101101001100010;
    rom[7677] = 25'b0001000011100100100111111;
    rom[7678] = 25'b0001000100011100001010110;
    rom[7679] = 25'b0001000101010011110100110;
    rom[7680] = 25'b0001000110001011100110010;
    rom[7681] = 25'b0001000111000011011110101;
    rom[7682] = 25'b0001000111111011011110011;
    rom[7683] = 25'b0001001000110011100101001;
    rom[7684] = 25'b0001001001101011110011000;
    rom[7685] = 25'b0001001010100100000111110;
    rom[7686] = 25'b0001001011011100100011100;
    rom[7687] = 25'b0001001100010101000110001;
    rom[7688] = 25'b0001001101001101101111101;
    rom[7689] = 25'b0001001110000110100000000;
    rom[7690] = 25'b0001001110111111010110111;
    rom[7691] = 25'b0001001111111000010100101;
    rom[7692] = 25'b0001010000110001011001001;
    rom[7693] = 25'b0001010001101010100100010;
    rom[7694] = 25'b0001010010100011110101110;
    rom[7695] = 25'b0001010011011101001101111;
    rom[7696] = 25'b0001010100010110101100011;
    rom[7697] = 25'b0001010101010000010001011;
    rom[7698] = 25'b0001010110001001111100110;
    rom[7699] = 25'b0001010111000011101110011;
    rom[7700] = 25'b0001010111111101100110011;
    rom[7701] = 25'b0001011000110111100100100;
    rom[7702] = 25'b0001011001110001101000111;
    rom[7703] = 25'b0001011010101011110011010;
    rom[7704] = 25'b0001011011100110000011111;
    rom[7705] = 25'b0001011100100000011010011;
    rom[7706] = 25'b0001011101011010110110111;
    rom[7707] = 25'b0001011110010101011001011;
    rom[7708] = 25'b0001011111010000000001101;
    rom[7709] = 25'b0001100000001010101111101;
    rom[7710] = 25'b0001100001000101100011100;
    rom[7711] = 25'b0001100010000000011101001;
    rom[7712] = 25'b0001100010111011011100011;
    rom[7713] = 25'b0001100011110110100001010;
    rom[7714] = 25'b0001100100110001101011101;
    rom[7715] = 25'b0001100101101100111011101;
    rom[7716] = 25'b0001100110101000010000111;
    rom[7717] = 25'b0001100111100011101011110;
    rom[7718] = 25'b0001101000011111001011111;
    rom[7719] = 25'b0001101001011010110001001;
    rom[7720] = 25'b0001101010010110011011110;
    rom[7721] = 25'b0001101011010010001011101;
    rom[7722] = 25'b0001101100001110000000101;
    rom[7723] = 25'b0001101101001001111010101;
    rom[7724] = 25'b0001101110000101111001110;
    rom[7725] = 25'b0001101111000001111101110;
    rom[7726] = 25'b0001101111111110000110110;
    rom[7727] = 25'b0001110000111010010100100;
    rom[7728] = 25'b0001110001110110100111010;
    rom[7729] = 25'b0001110010110010111110101;
    rom[7730] = 25'b0001110011101111011010110;
    rom[7731] = 25'b0001110100101011111011100;
    rom[7732] = 25'b0001110101101000100000110;
    rom[7733] = 25'b0001110110100101001010101;
    rom[7734] = 25'b0001110111100001111001000;
    rom[7735] = 25'b0001111000011110101011110;
    rom[7736] = 25'b0001111001011011100011000;
    rom[7737] = 25'b0001111010011000011110011;
    rom[7738] = 25'b0001111011010101011110010;
    rom[7739] = 25'b0001111100010010100010001;
    rom[7740] = 25'b0001111101001111101010010;
    rom[7741] = 25'b0001111110001100110110011;
    rom[7742] = 25'b0001111111001010000110101;
    rom[7743] = 25'b0010000000000111011010110;
    rom[7744] = 25'b0010000001000100110010111;
    rom[7745] = 25'b0010000010000010001110111;
    rom[7746] = 25'b0010000010111111101110101;
    rom[7747] = 25'b0010000011111101010010001;
    rom[7748] = 25'b0010000100111010111001011;
    rom[7749] = 25'b0010000101111000100100010;
    rom[7750] = 25'b0010000110110110010010110;
    rom[7751] = 25'b0010000111110100000100110;
    rom[7752] = 25'b0010001000110001111010001;
    rom[7753] = 25'b0010001001101111110011000;
    rom[7754] = 25'b0010001010101101101111010;
    rom[7755] = 25'b0010001011101011101110110;
    rom[7756] = 25'b0010001100101001110001011;
    rom[7757] = 25'b0010001101100111110111011;
    rom[7758] = 25'b0010001110100110000000011;
    rom[7759] = 25'b0010001111100100001100011;
    rom[7760] = 25'b0010010000100010011011100;
    rom[7761] = 25'b0010010001100000101101100;
    rom[7762] = 25'b0010010010011111000010011;
    rom[7763] = 25'b0010010011011101011010001;
    rom[7764] = 25'b0010010100011011110100101;
    rom[7765] = 25'b0010010101011010010001111;
    rom[7766] = 25'b0010010110011000110001101;
    rom[7767] = 25'b0010010111010111010100001;
    rom[7768] = 25'b0010011000010101111001000;
    rom[7769] = 25'b0010011001010100100000011;
    rom[7770] = 25'b0010011010010011001010010;
    rom[7771] = 25'b0010011011010001110110011;
    rom[7772] = 25'b0010011100010000100100111;
    rom[7773] = 25'b0010011101001111010101100;
    rom[7774] = 25'b0010011110001110001000011;
    rom[7775] = 25'b0010011111001100111101010;
    rom[7776] = 25'b0010100000001011110100010;
    rom[7777] = 25'b0010100001001010101101010;
    rom[7778] = 25'b0010100010001001101000001;
    rom[7779] = 25'b0010100011001000100101000;
    rom[7780] = 25'b0010100100000111100011101;
    rom[7781] = 25'b0010100101000110100011110;
    rom[7782] = 25'b0010100110000101100101110;
    rom[7783] = 25'b0010100111000100101001011;
    rom[7784] = 25'b0010101000000011101110101;
    rom[7785] = 25'b0010101001000010110101011;
    rom[7786] = 25'b0010101010000001111101011;
    rom[7787] = 25'b0010101011000001000110111;
    rom[7788] = 25'b0010101100000000010001110;
    rom[7789] = 25'b0010101100111111011101110;
    rom[7790] = 25'b0010101101111110101010111;
    rom[7791] = 25'b0010101110111101111001010;
    rom[7792] = 25'b0010101111111101001000110;
    rom[7793] = 25'b0010110000111100011001001;
    rom[7794] = 25'b0010110001111011101010100;
    rom[7795] = 25'b0010110010111010111100110;
    rom[7796] = 25'b0010110011111010001111111;
    rom[7797] = 25'b0010110100111001100011101;
    rom[7798] = 25'b0010110101111000111000001;
    rom[7799] = 25'b0010110110111000001101011;
    rom[7800] = 25'b0010110111110111100011000;
    rom[7801] = 25'b0010111000110110111001010;
    rom[7802] = 25'b0010111001110110001111111;
    rom[7803] = 25'b0010111010110101100111000;
    rom[7804] = 25'b0010111011110100111110011;
    rom[7805] = 25'b0010111100110100010110000;
    rom[7806] = 25'b0010111101110011101101110;
    rom[7807] = 25'b0010111110110011000101101;
    rom[7808] = 25'b0010111111110010011101110;
    rom[7809] = 25'b0011000000110001110101110;
    rom[7810] = 25'b0011000001110001001101101;
    rom[7811] = 25'b0011000010110000100101100;
    rom[7812] = 25'b0011000011101111111101000;
    rom[7813] = 25'b0011000100101111010100100;
    rom[7814] = 25'b0011000101101110101011100;
    rom[7815] = 25'b0011000110101110000010010;
    rom[7816] = 25'b0011000111101101011000100;
    rom[7817] = 25'b0011001000101100101110010;
    rom[7818] = 25'b0011001001101100000011011;
    rom[7819] = 25'b0011001010101011011000000;
    rom[7820] = 25'b0011001011101010101011111;
    rom[7821] = 25'b0011001100101001111110111;
    rom[7822] = 25'b0011001101101001010001001;
    rom[7823] = 25'b0011001110101000100010101;
    rom[7824] = 25'b0011001111100111110011000;
    rom[7825] = 25'b0011010000100111000010011;
    rom[7826] = 25'b0011010001100110010000110;
    rom[7827] = 25'b0011010010100101011101111;
    rom[7828] = 25'b0011010011100100101001111;
    rom[7829] = 25'b0011010100100011110100101;
    rom[7830] = 25'b0011010101100010111110000;
    rom[7831] = 25'b0011010110100010000110000;
    rom[7832] = 25'b0011010111100001001100100;
    rom[7833] = 25'b0011011000100000010001100;
    rom[7834] = 25'b0011011001011111010100111;
    rom[7835] = 25'b0011011010011110010110101;
    rom[7836] = 25'b0011011011011101010110101;
    rom[7837] = 25'b0011011100011100010101000;
    rom[7838] = 25'b0011011101011011010001011;
    rom[7839] = 25'b0011011110011010001011110;
    rom[7840] = 25'b0011011111011001000100010;
    rom[7841] = 25'b0011100000010111111010110;
    rom[7842] = 25'b0011100001010110101111001;
    rom[7843] = 25'b0011100010010101100001010;
    rom[7844] = 25'b0011100011010100010001010;
    rom[7845] = 25'b0011100100010010111110111;
    rom[7846] = 25'b0011100101010001101010010;
    rom[7847] = 25'b0011100110010000010011000;
    rom[7848] = 25'b0011100111001110111001011;
    rom[7849] = 25'b0011101000001101011101010;
    rom[7850] = 25'b0011101001001011111110011;
    rom[7851] = 25'b0011101010001010011100111;
    rom[7852] = 25'b0011101011001000111000101;
    rom[7853] = 25'b0011101100000111010001101;
    rom[7854] = 25'b0011101101000101100111101;
    rom[7855] = 25'b0011101110000011111010110;
    rom[7856] = 25'b0011101111000010001010111;
    rom[7857] = 25'b0011110000000000010111111;
    rom[7858] = 25'b0011110000111110100001110;
    rom[7859] = 25'b0011110001111100101000100;
    rom[7860] = 25'b0011110010111010101011111;
    rom[7861] = 25'b0011110011111000101100000;
    rom[7862] = 25'b0011110100110110101000110;
    rom[7863] = 25'b0011110101110100100010000;
    rom[7864] = 25'b0011110110110010010111101;
    rom[7865] = 25'b0011110111110000001001110;
    rom[7866] = 25'b0011111000101101111000010;
    rom[7867] = 25'b0011111001101011100011000;
    rom[7868] = 25'b0011111010101001001010000;
    rom[7869] = 25'b0011111011100110101101000;
    rom[7870] = 25'b0011111100100100001100010;
    rom[7871] = 25'b0011111101100001100111100;
    rom[7872] = 25'b0011111110011110111110101;
    rom[7873] = 25'b0011111111011100010001111;
    rom[7874] = 25'b0100000000011001100000110;
    rom[7875] = 25'b0100000001010110101011100;
    rom[7876] = 25'b0100000010010011110001111;
    rom[7877] = 25'b0100000011010000110011111;
    rom[7878] = 25'b0100000100001101110001100;
    rom[7879] = 25'b0100000101001010101010101;
    rom[7880] = 25'b0100000110000111011111010;
    rom[7881] = 25'b0100000111000100001111001;
    rom[7882] = 25'b0100001000000000111010011;
    rom[7883] = 25'b0100001000111101100000111;
    rom[7884] = 25'b0100001001111010000010101;
    rom[7885] = 25'b0100001010110110011111011;
    rom[7886] = 25'b0100001011110010110111011;
    rom[7887] = 25'b0100001100101111001010010;
    rom[7888] = 25'b0100001101101011011000001;
    rom[7889] = 25'b0100001110100111100000110;
    rom[7890] = 25'b0100001111100011100100010;
    rom[7891] = 25'b0100010000011111100010100;
    rom[7892] = 25'b0100010001011011011011100;
    rom[7893] = 25'b0100010010010111001111000;
    rom[7894] = 25'b0100010011010010111101001;
    rom[7895] = 25'b0100010100001110100101110;
    rom[7896] = 25'b0100010101001010001000110;
    rom[7897] = 25'b0100010110000101100110001;
    rom[7898] = 25'b0100010111000000111101110;
    rom[7899] = 25'b0100010111111100001111110;
    rom[7900] = 25'b0100011000110111011011111;
    rom[7901] = 25'b0100011001110010100010000;
    rom[7902] = 25'b0100011010101101100010010;
    rom[7903] = 25'b0100011011101000011100100;
    rom[7904] = 25'b0100011100100011010000110;
    rom[7905] = 25'b0100011101011101111110110;
    rom[7906] = 25'b0100011110011000100110100;
    rom[7907] = 25'b0100011111010011001000001;
    rom[7908] = 25'b0100100000001101100011011;
    rom[7909] = 25'b0100100001000111111000000;
    rom[7910] = 25'b0100100010000010000110100;
    rom[7911] = 25'b0100100010111100001110010;
    rom[7912] = 25'b0100100011110110001111100;
    rom[7913] = 25'b0100100100110000001010010;
    rom[7914] = 25'b0100100101101001111110001;
    rom[7915] = 25'b0100100110100011101011010;
    rom[7916] = 25'b0100100111011101010001101;
    rom[7917] = 25'b0100101000010110110001000;
    rom[7918] = 25'b0100101001010000001001101;
    rom[7919] = 25'b0100101010001001011011000;
    rom[7920] = 25'b0100101011000010100101100;
    rom[7921] = 25'b0100101011111011101000110;
    rom[7922] = 25'b0100101100110100100100110;
    rom[7923] = 25'b0100101101101101011001100;
    rom[7924] = 25'b0100101110100110000111000;
    rom[7925] = 25'b0100101111011110101101010;
    rom[7926] = 25'b0100110000010111001011110;
    rom[7927] = 25'b0100110001001111100011000;
    rom[7928] = 25'b0100110010000111110010100;
    rom[7929] = 25'b0100110010111111111010100;
    rom[7930] = 25'b0100110011110111111010110;
    rom[7931] = 25'b0100110100101111110011010;
    rom[7932] = 25'b0100110101100111100100000;
    rom[7933] = 25'b0100110110011111001100111;
    rom[7934] = 25'b0100110111010110101101110;
    rom[7935] = 25'b0100111000001110000110110;
    rom[7936] = 25'b0100111001000101010111101;
    rom[7937] = 25'b0100111001111100100000011;
    rom[7938] = 25'b0100111010110011100001000;
    rom[7939] = 25'b0100111011101010011001010;
    rom[7940] = 25'b0100111100100001001001011;
    rom[7941] = 25'b0100111101010111110001001;
    rom[7942] = 25'b0100111110001110010000011;
    rom[7943] = 25'b0100111111000100100111010;
    rom[7944] = 25'b0100111111111010110101101;
    rom[7945] = 25'b0101000000110000111011011;
    rom[7946] = 25'b0101000001100110111000100;
    rom[7947] = 25'b0101000010011100101100110;
    rom[7948] = 25'b0101000011010010011000100;
    rom[7949] = 25'b0101000100000111111011010;
    rom[7950] = 25'b0101000100111101010101001;
    rom[7951] = 25'b0101000101110010100110001;
    rom[7952] = 25'b0101000110100111101110001;
    rom[7953] = 25'b0101000111011100101101000;
    rom[7954] = 25'b0101001000010001100010111;
    rom[7955] = 25'b0101001001000110001111100;
    rom[7956] = 25'b0101001001111010110011000;
    rom[7957] = 25'b0101001010101111001101000;
    rom[7958] = 25'b0101001011100011011101111;
    rom[7959] = 25'b0101001100010111100101010;
    rom[7960] = 25'b0101001101001011100011010;
    rom[7961] = 25'b0101001101111111010111101;
    rom[7962] = 25'b0101001110110011000010100;
    rom[7963] = 25'b0101001111100110100011110;
    rom[7964] = 25'b0101010000011001111011010;
    rom[7965] = 25'b0101010001001101001001000;
    rom[7966] = 25'b0101010010000000001101000;
    rom[7967] = 25'b0101010010110011000111010;
    rom[7968] = 25'b0101010011100101110111100;
    rom[7969] = 25'b0101010100011000011101110;
    rom[7970] = 25'b0101010101001010111001111;
    rom[7971] = 25'b0101010101111101001100001;
    rom[7972] = 25'b0101010110101111010100001;
    rom[7973] = 25'b0101010111100001010010000;
    rom[7974] = 25'b0101011000010011000101101;
    rom[7975] = 25'b0101011001000100101110111;
    rom[7976] = 25'b0101011001110110001101111;
    rom[7977] = 25'b0101011010100111100010011;
    rom[7978] = 25'b0101011011011000101100100;
    rom[7979] = 25'b0101011100001001101100001;
    rom[7980] = 25'b0101011100111010100001000;
    rom[7981] = 25'b0101011101101011001011100;
    rom[7982] = 25'b0101011110011011101011001;
    rom[7983] = 25'b0101011111001100000000000;
    rom[7984] = 25'b0101011111111100001010010;
    rom[7985] = 25'b0101100000101100001001100;
    rom[7986] = 25'b0101100001011011111110000;
    rom[7987] = 25'b0101100010001011100111100;
    rom[7988] = 25'b0101100010111011000110000;
    rom[7989] = 25'b0101100011101010011001100;
    rom[7990] = 25'b0101100100011001100001110;
    rom[7991] = 25'b0101100101001000011111000;
    rom[7992] = 25'b0101100101110111010001000;
    rom[7993] = 25'b0101100110100101110111101;
    rom[7994] = 25'b0101100111010100010011001;
    rom[7995] = 25'b0101101000000010100011001;
    rom[7996] = 25'b0101101000110000100111110;
    rom[7997] = 25'b0101101001011110100000111;
    rom[7998] = 25'b0101101010001100001110101;
    rom[7999] = 25'b0101101010111001110000101;
    rom[8000] = 25'b0101101011100111000111001;
    rom[8001] = 25'b0101101100010100010001111;
    rom[8002] = 25'b0101101101000001010001000;
    rom[8003] = 25'b0101101101101110000100010;
    rom[8004] = 25'b0101101110011010101011110;
    rom[8005] = 25'b0101101111000111000111011;
    rom[8006] = 25'b0101101111110011010111001;
    rom[8007] = 25'b0101110000011111011010111;
    rom[8008] = 25'b0101110001001011010010100;
    rom[8009] = 25'b0101110001110110111110001;
    rom[8010] = 25'b0101110010100010011101110;
    rom[8011] = 25'b0101110011001101110001000;
    rom[8012] = 25'b0101110011111000111000001;
    rom[8013] = 25'b0101110100100011110011001;
    rom[8014] = 25'b0101110101001110100001101;
    rom[8015] = 25'b0101110101111001000011111;
    rom[8016] = 25'b0101110110100011011001110;
    rom[8017] = 25'b0101110111001101100011001;
    rom[8018] = 25'b0101110111110111100000000;
    rom[8019] = 25'b0101111000100001010000010;
    rom[8020] = 25'b0101111001001010110100000;
    rom[8021] = 25'b0101111001110100001011010;
    rom[8022] = 25'b0101111010011101010101101;
    rom[8023] = 25'b0101111011000110010011010;
    rom[8024] = 25'b0101111011101111000100001;
    rom[8025] = 25'b0101111100010111101000010;
    rom[8026] = 25'b0101111100111111111111100;
    rom[8027] = 25'b0101111101101000001001110;
    rom[8028] = 25'b0101111110010000000111001;
    rom[8029] = 25'b0101111110110111110111011;
    rom[8030] = 25'b0101111111011111011010110;
    rom[8031] = 25'b0110000000000110110000111;
    rom[8032] = 25'b0110000000101101111010000;
    rom[8033] = 25'b0110000001010100110101111;
    rom[8034] = 25'b0110000001111011100100101;
    rom[8035] = 25'b0110000010100010000110000;
    rom[8036] = 25'b0110000011001000011010000;
    rom[8037] = 25'b0110000011101110100000110;
    rom[8038] = 25'b0110000100010100011010001;
    rom[8039] = 25'b0110000100111010000110000;
    rom[8040] = 25'b0110000101011111100100011;
    rom[8041] = 25'b0110000110000100110101010;
    rom[8042] = 25'b0110000110101001111000101;
    rom[8043] = 25'b0110000111001110101110010;
    rom[8044] = 25'b0110000111110011010110011;
    rom[8045] = 25'b0110001000010111110000110;
    rom[8046] = 25'b0110001000111011111101010;
    rom[8047] = 25'b0110001001011111111100001;
    rom[8048] = 25'b0110001010000011101101010;
    rom[8049] = 25'b0110001010100111010000011;
    rom[8050] = 25'b0110001011001010100101101;
    rom[8051] = 25'b0110001011101101101101001;
    rom[8052] = 25'b0110001100010000100110011;
    rom[8053] = 25'b0110001100110011010001110;
    rom[8054] = 25'b0110001101010101101111001;
    rom[8055] = 25'b0110001101110111111110010;
    rom[8056] = 25'b0110001110011001111111100;
    rom[8057] = 25'b0110001110111011110010011;
    rom[8058] = 25'b0110001111011101010111001;
    rom[8059] = 25'b0110001111111110101101101;
    rom[8060] = 25'b0110010000011111110101110;
    rom[8061] = 25'b0110010001000000101111101;
    rom[8062] = 25'b0110010001100001011011010;
    rom[8063] = 25'b0110010010000001111000011;
    rom[8064] = 25'b0110010010100010000111000;
    rom[8065] = 25'b0110010011000010000111010;
    rom[8066] = 25'b0110010011100001111001000;
    rom[8067] = 25'b0110010100000001011100001;
    rom[8068] = 25'b0110010100100000110000110;
    rom[8069] = 25'b0110010100111111110110110;
    rom[8070] = 25'b0110010101011110101110001;
    rom[8071] = 25'b0110010101111101010110110;
    rom[8072] = 25'b0110010110011011110000110;
    rom[8073] = 25'b0110010110111001111100000;
    rom[8074] = 25'b0110010111010111111000011;
    rom[8075] = 25'b0110010111110101100110000;
    rom[8076] = 25'b0110011000010011000100101;
    rom[8077] = 25'b0110011000110000010100100;
    rom[8078] = 25'b0110011001001101010101100;
    rom[8079] = 25'b0110011001101010000111100;
    rom[8080] = 25'b0110011010000110101010100;
    rom[8081] = 25'b0110011010100010111110100;
    rom[8082] = 25'b0110011010111111000011011;
    rom[8083] = 25'b0110011011011010111001010;
    rom[8084] = 25'b0110011011110110100000001;
    rom[8085] = 25'b0110011100010001110111110;
    rom[8086] = 25'b0110011100101101000000001;
    rom[8087] = 25'b0110011101000111111001010;
    rom[8088] = 25'b0110011101100010100011010;
    rom[8089] = 25'b0110011101111100111110001;
    rom[8090] = 25'b0110011110010111001001100;
    rom[8091] = 25'b0110011110110001000101100;
    rom[8092] = 25'b0110011111001010110010010;
    rom[8093] = 25'b0110011111100100001111101;
    rom[8094] = 25'b0110011111111101011101100;
    rom[8095] = 25'b0110100000010110011100000;
    rom[8096] = 25'b0110100000101111001011001;
    rom[8097] = 25'b0110100001000111101010101;
    rom[8098] = 25'b0110100001011111111010101;
    rom[8099] = 25'b0110100001110111111011001;
    rom[8100] = 25'b0110100010001111101011111;
    rom[8101] = 25'b0110100010100111001101001;
    rom[8102] = 25'b0110100010111110011110111;
    rom[8103] = 25'b0110100011010101100000110;
    rom[8104] = 25'b0110100011101100010011000;
    rom[8105] = 25'b0110100100000010110101101;
    rom[8106] = 25'b0110100100011001001000011;
    rom[8107] = 25'b0110100100101111001011100;
    rom[8108] = 25'b0110100101000100111110110;
    rom[8109] = 25'b0110100101011010100010001;
    rom[8110] = 25'b0110100101101111110101101;
    rom[8111] = 25'b0110100110000100111001011;
    rom[8112] = 25'b0110100110011001101101010;
    rom[8113] = 25'b0110100110101110010001010;
    rom[8114] = 25'b0110100111000010100101010;
    rom[8115] = 25'b0110100111010110101001010;
    rom[8116] = 25'b0110100111101010011101010;
    rom[8117] = 25'b0110100111111110000001010;
    rom[8118] = 25'b0110101000010001010101011;
    rom[8119] = 25'b0110101000100100011001010;
    rom[8120] = 25'b0110101000110111001101001;
    rom[8121] = 25'b0110101001001001110001000;
    rom[8122] = 25'b0110101001011100000100101;
    rom[8123] = 25'b0110101001101110001000001;
    rom[8124] = 25'b0110101001111111111011101;
    rom[8125] = 25'b0110101010010001011110110;
    rom[8126] = 25'b0110101010100010110001111;
    rom[8127] = 25'b0110101010110011110100101;
    rom[8128] = 25'b0110101011000100100111010;
    rom[8129] = 25'b0110101011010101001001100;
    rom[8130] = 25'b0110101011100101011011101;
    rom[8131] = 25'b0110101011110101011101011;
    rom[8132] = 25'b0110101100000101001110110;
    rom[8133] = 25'b0110101100010100101111111;
    rom[8134] = 25'b0110101100100100000000101;
    rom[8135] = 25'b0110101100110011000001000;
    rom[8136] = 25'b0110101101000001110001001;
    rom[8137] = 25'b0110101101010000010000110;
    rom[8138] = 25'b0110101101011110100000000;
    rom[8139] = 25'b0110101101101100011110110;
    rom[8140] = 25'b0110101101111010001101000;
    rom[8141] = 25'b0110101110000111101010111;
    rom[8142] = 25'b0110101110010100111000011;
    rom[8143] = 25'b0110101110100001110101010;
    rom[8144] = 25'b0110101110101110100001101;
    rom[8145] = 25'b0110101110111010111101100;
    rom[8146] = 25'b0110101111000111001000110;
    rom[8147] = 25'b0110101111010011000011101;
    rom[8148] = 25'b0110101111011110101101111;
    rom[8149] = 25'b0110101111101010000111100;
    rom[8150] = 25'b0110101111110101010000100;
    rom[8151] = 25'b0110110000000000001001000;
    rom[8152] = 25'b0110110000001010110000111;
    rom[8153] = 25'b0110110000010101001000000;
    rom[8154] = 25'b0110110000011111001110101;
    rom[8155] = 25'b0110110000101001000100100;
    rom[8156] = 25'b0110110000110010101001111;
    rom[8157] = 25'b0110110000111011111110011;
    rom[8158] = 25'b0110110001000101000010010;
    rom[8159] = 25'b0110110001001101110101100;
    rom[8160] = 25'b0110110001010110011000000;
    rom[8161] = 25'b0110110001011110101001111;
    rom[8162] = 25'b0110110001100110101010111;
    rom[8163] = 25'b0110110001101110011011001;
    rom[8164] = 25'b0110110001110101111010110;
    rom[8165] = 25'b0110110001111101001001101;
    rom[8166] = 25'b0110110010000100000111110;
    rom[8167] = 25'b0110110010001010110101000;
    rom[8168] = 25'b0110110010010001010001101;
    rom[8169] = 25'b0110110010010111011101010;
    rom[8170] = 25'b0110110010011101011000010;
    rom[8171] = 25'b0110110010100011000010100;
    rom[8172] = 25'b0110110010101000011011111;
    rom[8173] = 25'b0110110010101101100100011;
    rom[8174] = 25'b0110110010110010011100001;
    rom[8175] = 25'b0110110010110111000011000;
    rom[8176] = 25'b0110110010111011011001001;
    rom[8177] = 25'b0110110010111111011110100;
    rom[8178] = 25'b0110110011000011010010111;
    rom[8179] = 25'b0110110011000110110110100;
    rom[8180] = 25'b0110110011001010001001011;
    rom[8181] = 25'b0110110011001101001011010;
    rom[8182] = 25'b0110110011001111111100010;
    rom[8183] = 25'b0110110011010010011100100;
    rom[8184] = 25'b0110110011010100101011111;
    rom[8185] = 25'b0110110011010110101010010;
    rom[8186] = 25'b0110110011011000011000000;
    rom[8187] = 25'b0110110011011001110100110;
    rom[8188] = 25'b0110110011011011000000101;
    rom[8189] = 25'b0110110011011011111011101;
    rom[8190] = 25'b0110110011011100100101110;
    rom[8191] = 25'b0110110011011100111111001;
    rom[8192] = 25'b0110110011011101000111101;
    rom[8193] = 25'b0110110011011100111111001;
    rom[8194] = 25'b0110110011011100100101110;
    rom[8195] = 25'b0110110011011011111011101;
    rom[8196] = 25'b0110110011011011000000101;
    rom[8197] = 25'b0110110011011001110100110;
    rom[8198] = 25'b0110110011011000011000000;
    rom[8199] = 25'b0110110011010110101010010;
    rom[8200] = 25'b0110110011010100101011111;
    rom[8201] = 25'b0110110011010010011100100;
    rom[8202] = 25'b0110110011001111111100010;
    rom[8203] = 25'b0110110011001101001011010;
    rom[8204] = 25'b0110110011001010001001011;
    rom[8205] = 25'b0110110011000110110110100;
    rom[8206] = 25'b0110110011000011010010111;
    rom[8207] = 25'b0110110010111111011110100;
    rom[8208] = 25'b0110110010111011011001001;
    rom[8209] = 25'b0110110010110111000011000;
    rom[8210] = 25'b0110110010110010011100001;
    rom[8211] = 25'b0110110010101101100100011;
    rom[8212] = 25'b0110110010101000011011111;
    rom[8213] = 25'b0110110010100011000010100;
    rom[8214] = 25'b0110110010011101011000010;
    rom[8215] = 25'b0110110010010111011101010;
    rom[8216] = 25'b0110110010010001010001101;
    rom[8217] = 25'b0110110010001010110101000;
    rom[8218] = 25'b0110110010000100000111110;
    rom[8219] = 25'b0110110001111101001001101;
    rom[8220] = 25'b0110110001110101111010110;
    rom[8221] = 25'b0110110001101110011011001;
    rom[8222] = 25'b0110110001100110101010111;
    rom[8223] = 25'b0110110001011110101001111;
    rom[8224] = 25'b0110110001010110011000000;
    rom[8225] = 25'b0110110001001101110101100;
    rom[8226] = 25'b0110110001000101000010010;
    rom[8227] = 25'b0110110000111011111110011;
    rom[8228] = 25'b0110110000110010101001111;
    rom[8229] = 25'b0110110000101001000100100;
    rom[8230] = 25'b0110110000011111001110101;
    rom[8231] = 25'b0110110000010101001000000;
    rom[8232] = 25'b0110110000001010110000111;
    rom[8233] = 25'b0110110000000000001001000;
    rom[8234] = 25'b0110101111110101010000100;
    rom[8235] = 25'b0110101111101010000111100;
    rom[8236] = 25'b0110101111011110101101111;
    rom[8237] = 25'b0110101111010011000011101;
    rom[8238] = 25'b0110101111000111001000110;
    rom[8239] = 25'b0110101110111010111101100;
    rom[8240] = 25'b0110101110101110100001101;
    rom[8241] = 25'b0110101110100001110101010;
    rom[8242] = 25'b0110101110010100111000011;
    rom[8243] = 25'b0110101110000111101010111;
    rom[8244] = 25'b0110101101111010001101000;
    rom[8245] = 25'b0110101101101100011110110;
    rom[8246] = 25'b0110101101011110100000000;
    rom[8247] = 25'b0110101101010000010000110;
    rom[8248] = 25'b0110101101000001110001001;
    rom[8249] = 25'b0110101100110011000001000;
    rom[8250] = 25'b0110101100100100000000101;
    rom[8251] = 25'b0110101100010100101111111;
    rom[8252] = 25'b0110101100000101001110110;
    rom[8253] = 25'b0110101011110101011101011;
    rom[8254] = 25'b0110101011100101011011101;
    rom[8255] = 25'b0110101011010101001001100;
    rom[8256] = 25'b0110101011000100100111010;
    rom[8257] = 25'b0110101010110011110100101;
    rom[8258] = 25'b0110101010100010110001111;
    rom[8259] = 25'b0110101010010001011110110;
    rom[8260] = 25'b0110101001111111111011101;
    rom[8261] = 25'b0110101001101110001000001;
    rom[8262] = 25'b0110101001011100000100101;
    rom[8263] = 25'b0110101001001001110001000;
    rom[8264] = 25'b0110101000110111001101001;
    rom[8265] = 25'b0110101000100100011001010;
    rom[8266] = 25'b0110101000010001010101011;
    rom[8267] = 25'b0110100111111110000001010;
    rom[8268] = 25'b0110100111101010011101010;
    rom[8269] = 25'b0110100111010110101001010;
    rom[8270] = 25'b0110100111000010100101010;
    rom[8271] = 25'b0110100110101110010001010;
    rom[8272] = 25'b0110100110011001101101010;
    rom[8273] = 25'b0110100110000100111001011;
    rom[8274] = 25'b0110100101101111110101101;
    rom[8275] = 25'b0110100101011010100010001;
    rom[8276] = 25'b0110100101000100111110110;
    rom[8277] = 25'b0110100100101111001011100;
    rom[8278] = 25'b0110100100011001001000011;
    rom[8279] = 25'b0110100100000010110101101;
    rom[8280] = 25'b0110100011101100010011000;
    rom[8281] = 25'b0110100011010101100000110;
    rom[8282] = 25'b0110100010111110011110111;
    rom[8283] = 25'b0110100010100111001101001;
    rom[8284] = 25'b0110100010001111101011111;
    rom[8285] = 25'b0110100001110111111011001;
    rom[8286] = 25'b0110100001011111111010101;
    rom[8287] = 25'b0110100001000111101010101;
    rom[8288] = 25'b0110100000101111001011001;
    rom[8289] = 25'b0110100000010110011100000;
    rom[8290] = 25'b0110011111111101011101100;
    rom[8291] = 25'b0110011111100100001111101;
    rom[8292] = 25'b0110011111001010110010010;
    rom[8293] = 25'b0110011110110001000101100;
    rom[8294] = 25'b0110011110010111001001100;
    rom[8295] = 25'b0110011101111100111110001;
    rom[8296] = 25'b0110011101100010100011010;
    rom[8297] = 25'b0110011101000111111001010;
    rom[8298] = 25'b0110011100101101000000001;
    rom[8299] = 25'b0110011100010001110111110;
    rom[8300] = 25'b0110011011110110100000001;
    rom[8301] = 25'b0110011011011010111001010;
    rom[8302] = 25'b0110011010111111000011011;
    rom[8303] = 25'b0110011010100010111110100;
    rom[8304] = 25'b0110011010000110101010100;
    rom[8305] = 25'b0110011001101010000111100;
    rom[8306] = 25'b0110011001001101010101100;
    rom[8307] = 25'b0110011000110000010100100;
    rom[8308] = 25'b0110011000010011000100101;
    rom[8309] = 25'b0110010111110101100110000;
    rom[8310] = 25'b0110010111010111111000011;
    rom[8311] = 25'b0110010110111001111100000;
    rom[8312] = 25'b0110010110011011110000110;
    rom[8313] = 25'b0110010101111101010110110;
    rom[8314] = 25'b0110010101011110101110001;
    rom[8315] = 25'b0110010100111111110110110;
    rom[8316] = 25'b0110010100100000110000110;
    rom[8317] = 25'b0110010100000001011100001;
    rom[8318] = 25'b0110010011100001111001000;
    rom[8319] = 25'b0110010011000010000111010;
    rom[8320] = 25'b0110010010100010000111000;
    rom[8321] = 25'b0110010010000001111000011;
    rom[8322] = 25'b0110010001100001011011010;
    rom[8323] = 25'b0110010001000000101111101;
    rom[8324] = 25'b0110010000011111110101110;
    rom[8325] = 25'b0110001111111110101101101;
    rom[8326] = 25'b0110001111011101010111001;
    rom[8327] = 25'b0110001110111011110010011;
    rom[8328] = 25'b0110001110011001111111100;
    rom[8329] = 25'b0110001101110111111110010;
    rom[8330] = 25'b0110001101010101101111001;
    rom[8331] = 25'b0110001100110011010001110;
    rom[8332] = 25'b0110001100010000100110011;
    rom[8333] = 25'b0110001011101101101101001;
    rom[8334] = 25'b0110001011001010100101101;
    rom[8335] = 25'b0110001010100111010000011;
    rom[8336] = 25'b0110001010000011101101010;
    rom[8337] = 25'b0110001001011111111100001;
    rom[8338] = 25'b0110001000111011111101010;
    rom[8339] = 25'b0110001000010111110000110;
    rom[8340] = 25'b0110000111110011010110011;
    rom[8341] = 25'b0110000111001110101110010;
    rom[8342] = 25'b0110000110101001111000101;
    rom[8343] = 25'b0110000110000100110101010;
    rom[8344] = 25'b0110000101011111100100011;
    rom[8345] = 25'b0110000100111010000110000;
    rom[8346] = 25'b0110000100010100011010001;
    rom[8347] = 25'b0110000011101110100000110;
    rom[8348] = 25'b0110000011001000011010000;
    rom[8349] = 25'b0110000010100010000110000;
    rom[8350] = 25'b0110000001111011100100101;
    rom[8351] = 25'b0110000001010100110101111;
    rom[8352] = 25'b0110000000101101111010000;
    rom[8353] = 25'b0110000000000110110000111;
    rom[8354] = 25'b0101111111011111011010110;
    rom[8355] = 25'b0101111110110111110111011;
    rom[8356] = 25'b0101111110010000000111001;
    rom[8357] = 25'b0101111101101000001001110;
    rom[8358] = 25'b0101111100111111111111100;
    rom[8359] = 25'b0101111100010111101000010;
    rom[8360] = 25'b0101111011101111000100001;
    rom[8361] = 25'b0101111011000110010011010;
    rom[8362] = 25'b0101111010011101010101101;
    rom[8363] = 25'b0101111001110100001011010;
    rom[8364] = 25'b0101111001001010110100000;
    rom[8365] = 25'b0101111000100001010000010;
    rom[8366] = 25'b0101110111110111100000000;
    rom[8367] = 25'b0101110111001101100011001;
    rom[8368] = 25'b0101110110100011011001110;
    rom[8369] = 25'b0101110101111001000011111;
    rom[8370] = 25'b0101110101001110100001101;
    rom[8371] = 25'b0101110100100011110011001;
    rom[8372] = 25'b0101110011111000111000001;
    rom[8373] = 25'b0101110011001101110001000;
    rom[8374] = 25'b0101110010100010011101110;
    rom[8375] = 25'b0101110001110110111110001;
    rom[8376] = 25'b0101110001001011010010100;
    rom[8377] = 25'b0101110000011111011010111;
    rom[8378] = 25'b0101101111110011010111001;
    rom[8379] = 25'b0101101111000111000111011;
    rom[8380] = 25'b0101101110011010101011110;
    rom[8381] = 25'b0101101101101110000100010;
    rom[8382] = 25'b0101101101000001010001000;
    rom[8383] = 25'b0101101100010100010001111;
    rom[8384] = 25'b0101101011100111000111001;
    rom[8385] = 25'b0101101010111001110000101;
    rom[8386] = 25'b0101101010001100001110101;
    rom[8387] = 25'b0101101001011110100000111;
    rom[8388] = 25'b0101101000110000100111110;
    rom[8389] = 25'b0101101000000010100011001;
    rom[8390] = 25'b0101100111010100010011001;
    rom[8391] = 25'b0101100110100101110111101;
    rom[8392] = 25'b0101100101110111010001000;
    rom[8393] = 25'b0101100101001000011111000;
    rom[8394] = 25'b0101100100011001100001110;
    rom[8395] = 25'b0101100011101010011001100;
    rom[8396] = 25'b0101100010111011000110000;
    rom[8397] = 25'b0101100010001011100111100;
    rom[8398] = 25'b0101100001011011111110000;
    rom[8399] = 25'b0101100000101100001001100;
    rom[8400] = 25'b0101011111111100001010010;
    rom[8401] = 25'b0101011111001100000000000;
    rom[8402] = 25'b0101011110011011101011001;
    rom[8403] = 25'b0101011101101011001011100;
    rom[8404] = 25'b0101011100111010100001000;
    rom[8405] = 25'b0101011100001001101100001;
    rom[8406] = 25'b0101011011011000101100100;
    rom[8407] = 25'b0101011010100111100010011;
    rom[8408] = 25'b0101011001110110001101111;
    rom[8409] = 25'b0101011001000100101110111;
    rom[8410] = 25'b0101011000010011000101101;
    rom[8411] = 25'b0101010111100001010010000;
    rom[8412] = 25'b0101010110101111010100001;
    rom[8413] = 25'b0101010101111101001100001;
    rom[8414] = 25'b0101010101001010111001111;
    rom[8415] = 25'b0101010100011000011101110;
    rom[8416] = 25'b0101010011100101110111100;
    rom[8417] = 25'b0101010010110011000111010;
    rom[8418] = 25'b0101010010000000001101000;
    rom[8419] = 25'b0101010001001101001001000;
    rom[8420] = 25'b0101010000011001111011010;
    rom[8421] = 25'b0101001111100110100011110;
    rom[8422] = 25'b0101001110110011000010100;
    rom[8423] = 25'b0101001101111111010111101;
    rom[8424] = 25'b0101001101001011100011010;
    rom[8425] = 25'b0101001100010111100101010;
    rom[8426] = 25'b0101001011100011011101111;
    rom[8427] = 25'b0101001010101111001101000;
    rom[8428] = 25'b0101001001111010110011000;
    rom[8429] = 25'b0101001001000110001111100;
    rom[8430] = 25'b0101001000010001100010111;
    rom[8431] = 25'b0101000111011100101101000;
    rom[8432] = 25'b0101000110100111101110001;
    rom[8433] = 25'b0101000101110010100110001;
    rom[8434] = 25'b0101000100111101010101001;
    rom[8435] = 25'b0101000100000111111011010;
    rom[8436] = 25'b0101000011010010011000100;
    rom[8437] = 25'b0101000010011100101100110;
    rom[8438] = 25'b0101000001100110111000100;
    rom[8439] = 25'b0101000000110000111011011;
    rom[8440] = 25'b0100111111111010110101101;
    rom[8441] = 25'b0100111111000100100111010;
    rom[8442] = 25'b0100111110001110010000011;
    rom[8443] = 25'b0100111101010111110001001;
    rom[8444] = 25'b0100111100100001001001011;
    rom[8445] = 25'b0100111011101010011001010;
    rom[8446] = 25'b0100111010110011100001000;
    rom[8447] = 25'b0100111001111100100000011;
    rom[8448] = 25'b0100111001000101010111101;
    rom[8449] = 25'b0100111000001110000110110;
    rom[8450] = 25'b0100110111010110101101110;
    rom[8451] = 25'b0100110110011111001100111;
    rom[8452] = 25'b0100110101100111100100000;
    rom[8453] = 25'b0100110100101111110011010;
    rom[8454] = 25'b0100110011110111111010110;
    rom[8455] = 25'b0100110010111111111010100;
    rom[8456] = 25'b0100110010000111110010100;
    rom[8457] = 25'b0100110001001111100011000;
    rom[8458] = 25'b0100110000010111001011110;
    rom[8459] = 25'b0100101111011110101101010;
    rom[8460] = 25'b0100101110100110000111000;
    rom[8461] = 25'b0100101101101101011001100;
    rom[8462] = 25'b0100101100110100100100110;
    rom[8463] = 25'b0100101011111011101000110;
    rom[8464] = 25'b0100101011000010100101100;
    rom[8465] = 25'b0100101010001001011011000;
    rom[8466] = 25'b0100101001010000001001101;
    rom[8467] = 25'b0100101000010110110001000;
    rom[8468] = 25'b0100100111011101010001101;
    rom[8469] = 25'b0100100110100011101011010;
    rom[8470] = 25'b0100100101101001111110001;
    rom[8471] = 25'b0100100100110000001010010;
    rom[8472] = 25'b0100100011110110001111100;
    rom[8473] = 25'b0100100010111100001110010;
    rom[8474] = 25'b0100100010000010000110100;
    rom[8475] = 25'b0100100001000111111000000;
    rom[8476] = 25'b0100100000001101100011011;
    rom[8477] = 25'b0100011111010011001000001;
    rom[8478] = 25'b0100011110011000100110100;
    rom[8479] = 25'b0100011101011101111110110;
    rom[8480] = 25'b0100011100100011010000110;
    rom[8481] = 25'b0100011011101000011100100;
    rom[8482] = 25'b0100011010101101100010010;
    rom[8483] = 25'b0100011001110010100010000;
    rom[8484] = 25'b0100011000110111011011111;
    rom[8485] = 25'b0100010111111100001111110;
    rom[8486] = 25'b0100010111000000111101110;
    rom[8487] = 25'b0100010110000101100110001;
    rom[8488] = 25'b0100010101001010001000110;
    rom[8489] = 25'b0100010100001110100101110;
    rom[8490] = 25'b0100010011010010111101001;
    rom[8491] = 25'b0100010010010111001111000;
    rom[8492] = 25'b0100010001011011011011100;
    rom[8493] = 25'b0100010000011111100010100;
    rom[8494] = 25'b0100001111100011100100010;
    rom[8495] = 25'b0100001110100111100000110;
    rom[8496] = 25'b0100001101101011011000001;
    rom[8497] = 25'b0100001100101111001010010;
    rom[8498] = 25'b0100001011110010110111011;
    rom[8499] = 25'b0100001010110110011111011;
    rom[8500] = 25'b0100001001111010000010101;
    rom[8501] = 25'b0100001000111101100000111;
    rom[8502] = 25'b0100001000000000111010011;
    rom[8503] = 25'b0100000111000100001111001;
    rom[8504] = 25'b0100000110000111011111010;
    rom[8505] = 25'b0100000101001010101010101;
    rom[8506] = 25'b0100000100001101110001100;
    rom[8507] = 25'b0100000011010000110011111;
    rom[8508] = 25'b0100000010010011110001111;
    rom[8509] = 25'b0100000001010110101011100;
    rom[8510] = 25'b0100000000011001100000110;
    rom[8511] = 25'b0011111111011100010001111;
    rom[8512] = 25'b0011111110011110111110101;
    rom[8513] = 25'b0011111101100001100111100;
    rom[8514] = 25'b0011111100100100001100010;
    rom[8515] = 25'b0011111011100110101101000;
    rom[8516] = 25'b0011111010101001001010000;
    rom[8517] = 25'b0011111001101011100011000;
    rom[8518] = 25'b0011111000101101111000010;
    rom[8519] = 25'b0011110111110000001001110;
    rom[8520] = 25'b0011110110110010010111101;
    rom[8521] = 25'b0011110101110100100010000;
    rom[8522] = 25'b0011110100110110101000110;
    rom[8523] = 25'b0011110011111000101100000;
    rom[8524] = 25'b0011110010111010101011111;
    rom[8525] = 25'b0011110001111100101000100;
    rom[8526] = 25'b0011110000111110100001110;
    rom[8527] = 25'b0011110000000000010111111;
    rom[8528] = 25'b0011101111000010001010111;
    rom[8529] = 25'b0011101110000011111010110;
    rom[8530] = 25'b0011101101000101100111101;
    rom[8531] = 25'b0011101100000111010001101;
    rom[8532] = 25'b0011101011001000111000101;
    rom[8533] = 25'b0011101010001010011100111;
    rom[8534] = 25'b0011101001001011111110011;
    rom[8535] = 25'b0011101000001101011101010;
    rom[8536] = 25'b0011100111001110111001011;
    rom[8537] = 25'b0011100110010000010011000;
    rom[8538] = 25'b0011100101010001101010010;
    rom[8539] = 25'b0011100100010010111110111;
    rom[8540] = 25'b0011100011010100010001010;
    rom[8541] = 25'b0011100010010101100001010;
    rom[8542] = 25'b0011100001010110101111001;
    rom[8543] = 25'b0011100000010111111010110;
    rom[8544] = 25'b0011011111011001000100010;
    rom[8545] = 25'b0011011110011010001011110;
    rom[8546] = 25'b0011011101011011010001011;
    rom[8547] = 25'b0011011100011100010101000;
    rom[8548] = 25'b0011011011011101010110101;
    rom[8549] = 25'b0011011010011110010110101;
    rom[8550] = 25'b0011011001011111010100111;
    rom[8551] = 25'b0011011000100000010001100;
    rom[8552] = 25'b0011010111100001001100100;
    rom[8553] = 25'b0011010110100010000110000;
    rom[8554] = 25'b0011010101100010111110000;
    rom[8555] = 25'b0011010100100011110100101;
    rom[8556] = 25'b0011010011100100101001111;
    rom[8557] = 25'b0011010010100101011101111;
    rom[8558] = 25'b0011010001100110010000110;
    rom[8559] = 25'b0011010000100111000010011;
    rom[8560] = 25'b0011001111100111110011000;
    rom[8561] = 25'b0011001110101000100010101;
    rom[8562] = 25'b0011001101101001010001001;
    rom[8563] = 25'b0011001100101001111110111;
    rom[8564] = 25'b0011001011101010101011111;
    rom[8565] = 25'b0011001010101011011000000;
    rom[8566] = 25'b0011001001101100000011011;
    rom[8567] = 25'b0011001000101100101110010;
    rom[8568] = 25'b0011000111101101011000100;
    rom[8569] = 25'b0011000110101110000010010;
    rom[8570] = 25'b0011000101101110101011100;
    rom[8571] = 25'b0011000100101111010100100;
    rom[8572] = 25'b0011000011101111111101000;
    rom[8573] = 25'b0011000010110000100101100;
    rom[8574] = 25'b0011000001110001001101101;
    rom[8575] = 25'b0011000000110001110101110;
    rom[8576] = 25'b0010111111110010011101110;
    rom[8577] = 25'b0010111110110011000101101;
    rom[8578] = 25'b0010111101110011101101110;
    rom[8579] = 25'b0010111100110100010110000;
    rom[8580] = 25'b0010111011110100111110011;
    rom[8581] = 25'b0010111010110101100111000;
    rom[8582] = 25'b0010111001110110001111111;
    rom[8583] = 25'b0010111000110110111001010;
    rom[8584] = 25'b0010110111110111100011000;
    rom[8585] = 25'b0010110110111000001101011;
    rom[8586] = 25'b0010110101111000111000001;
    rom[8587] = 25'b0010110100111001100011101;
    rom[8588] = 25'b0010110011111010001111111;
    rom[8589] = 25'b0010110010111010111100110;
    rom[8590] = 25'b0010110001111011101010100;
    rom[8591] = 25'b0010110000111100011001001;
    rom[8592] = 25'b0010101111111101001000110;
    rom[8593] = 25'b0010101110111101111001010;
    rom[8594] = 25'b0010101101111110101010111;
    rom[8595] = 25'b0010101100111111011101110;
    rom[8596] = 25'b0010101100000000010001110;
    rom[8597] = 25'b0010101011000001000110111;
    rom[8598] = 25'b0010101010000001111101011;
    rom[8599] = 25'b0010101001000010110101011;
    rom[8600] = 25'b0010101000000011101110101;
    rom[8601] = 25'b0010100111000100101001011;
    rom[8602] = 25'b0010100110000101100101110;
    rom[8603] = 25'b0010100101000110100011110;
    rom[8604] = 25'b0010100100000111100011101;
    rom[8605] = 25'b0010100011001000100101000;
    rom[8606] = 25'b0010100010001001101000001;
    rom[8607] = 25'b0010100001001010101101010;
    rom[8608] = 25'b0010100000001011110100010;
    rom[8609] = 25'b0010011111001100111101010;
    rom[8610] = 25'b0010011110001110001000011;
    rom[8611] = 25'b0010011101001111010101100;
    rom[8612] = 25'b0010011100010000100100111;
    rom[8613] = 25'b0010011011010001110110011;
    rom[8614] = 25'b0010011010010011001010010;
    rom[8615] = 25'b0010011001010100100000011;
    rom[8616] = 25'b0010011000010101111001000;
    rom[8617] = 25'b0010010111010111010100001;
    rom[8618] = 25'b0010010110011000110001101;
    rom[8619] = 25'b0010010101011010010001111;
    rom[8620] = 25'b0010010100011011110100101;
    rom[8621] = 25'b0010010011011101011010001;
    rom[8622] = 25'b0010010010011111000010011;
    rom[8623] = 25'b0010010001100000101101100;
    rom[8624] = 25'b0010010000100010011011100;
    rom[8625] = 25'b0010001111100100001100011;
    rom[8626] = 25'b0010001110100110000000011;
    rom[8627] = 25'b0010001101100111110111011;
    rom[8628] = 25'b0010001100101001110001011;
    rom[8629] = 25'b0010001011101011101110110;
    rom[8630] = 25'b0010001010101101101111010;
    rom[8631] = 25'b0010001001101111110011000;
    rom[8632] = 25'b0010001000110001111010001;
    rom[8633] = 25'b0010000111110100000100110;
    rom[8634] = 25'b0010000110110110010010110;
    rom[8635] = 25'b0010000101111000100100010;
    rom[8636] = 25'b0010000100111010111001011;
    rom[8637] = 25'b0010000011111101010010001;
    rom[8638] = 25'b0010000010111111101110101;
    rom[8639] = 25'b0010000010000010001110111;
    rom[8640] = 25'b0010000001000100110010111;
    rom[8641] = 25'b0010000000000111011010110;
    rom[8642] = 25'b0001111111001010000110101;
    rom[8643] = 25'b0001111110001100110110011;
    rom[8644] = 25'b0001111101001111101010010;
    rom[8645] = 25'b0001111100010010100010001;
    rom[8646] = 25'b0001111011010101011110010;
    rom[8647] = 25'b0001111010011000011110011;
    rom[8648] = 25'b0001111001011011100011000;
    rom[8649] = 25'b0001111000011110101011110;
    rom[8650] = 25'b0001110111100001111001000;
    rom[8651] = 25'b0001110110100101001010101;
    rom[8652] = 25'b0001110101101000100000110;
    rom[8653] = 25'b0001110100101011111011100;
    rom[8654] = 25'b0001110011101111011010110;
    rom[8655] = 25'b0001110010110010111110101;
    rom[8656] = 25'b0001110001110110100111010;
    rom[8657] = 25'b0001110000111010010100100;
    rom[8658] = 25'b0001101111111110000110110;
    rom[8659] = 25'b0001101111000001111101110;
    rom[8660] = 25'b0001101110000101111001110;
    rom[8661] = 25'b0001101101001001111010101;
    rom[8662] = 25'b0001101100001110000000101;
    rom[8663] = 25'b0001101011010010001011101;
    rom[8664] = 25'b0001101010010110011011110;
    rom[8665] = 25'b0001101001011010110001001;
    rom[8666] = 25'b0001101000011111001011111;
    rom[8667] = 25'b0001100111100011101011110;
    rom[8668] = 25'b0001100110101000010000111;
    rom[8669] = 25'b0001100101101100111011101;
    rom[8670] = 25'b0001100100110001101011101;
    rom[8671] = 25'b0001100011110110100001010;
    rom[8672] = 25'b0001100010111011011100011;
    rom[8673] = 25'b0001100010000000011101001;
    rom[8674] = 25'b0001100001000101100011100;
    rom[8675] = 25'b0001100000001010101111101;
    rom[8676] = 25'b0001011111010000000001101;
    rom[8677] = 25'b0001011110010101011001011;
    rom[8678] = 25'b0001011101011010110110111;
    rom[8679] = 25'b0001011100100000011010011;
    rom[8680] = 25'b0001011011100110000011111;
    rom[8681] = 25'b0001011010101011110011010;
    rom[8682] = 25'b0001011001110001101000111;
    rom[8683] = 25'b0001011000110111100100100;
    rom[8684] = 25'b0001010111111101100110011;
    rom[8685] = 25'b0001010111000011101110011;
    rom[8686] = 25'b0001010110001001111100110;
    rom[8687] = 25'b0001010101010000010001011;
    rom[8688] = 25'b0001010100010110101100011;
    rom[8689] = 25'b0001010011011101001101111;
    rom[8690] = 25'b0001010010100011110101110;
    rom[8691] = 25'b0001010001101010100100010;
    rom[8692] = 25'b0001010000110001011001001;
    rom[8693] = 25'b0001001111111000010100101;
    rom[8694] = 25'b0001001110111111010110111;
    rom[8695] = 25'b0001001110000110100000000;
    rom[8696] = 25'b0001001101001101101111101;
    rom[8697] = 25'b0001001100010101000110001;
    rom[8698] = 25'b0001001011011100100011100;
    rom[8699] = 25'b0001001010100100000111110;
    rom[8700] = 25'b0001001001101011110011000;
    rom[8701] = 25'b0001001000110011100101001;
    rom[8702] = 25'b0001000111111011011110011;
    rom[8703] = 25'b0001000111000011011110101;
    rom[8704] = 25'b0001000110001011100110010;
    rom[8705] = 25'b0001000101010011110100110;
    rom[8706] = 25'b0001000100011100001010110;
    rom[8707] = 25'b0001000011100100100111111;
    rom[8708] = 25'b0001000010101101001100010;
    rom[8709] = 25'b0001000001110101111000001;
    rom[8710] = 25'b0001000000111110101011011;
    rom[8711] = 25'b0001000000000111100101111;
    rom[8712] = 25'b0000111111010000101000001;
    rom[8713] = 25'b0000111110011001110001111;
    rom[8714] = 25'b0000111101100011000011001;
    rom[8715] = 25'b0000111100101100011100000;
    rom[8716] = 25'b0000111011110101111100101;
    rom[8717] = 25'b0000111010111111100101000;
    rom[8718] = 25'b0000111010001001010101000;
    rom[8719] = 25'b0000111001010011001101000;
    rom[8720] = 25'b0000111000011101001100101;
    rom[8721] = 25'b0000110111100111010100010;
    rom[8722] = 25'b0000110110110001100011110;
    rom[8723] = 25'b0000110101111011111011011;
    rom[8724] = 25'b0000110101000110011010111;
    rom[8725] = 25'b0000110100010001000010100;
    rom[8726] = 25'b0000110011011011110010010;
    rom[8727] = 25'b0000110010100110101010001;
    rom[8728] = 25'b0000110001110001101010001;
    rom[8729] = 25'b0000110000111100110010011;
    rom[8730] = 25'b0000110000001000000011000;
    rom[8731] = 25'b0000101111010011011011110;
    rom[8732] = 25'b0000101110011110111100111;
    rom[8733] = 25'b0000101101101010100110101;
    rom[8734] = 25'b0000101100110110011000100;
    rom[8735] = 25'b0000101100000010010011000;
    rom[8736] = 25'b0000101011001110010110000;
    rom[8737] = 25'b0000101010011010100001101;
    rom[8738] = 25'b0000101001100110110101101;
    rom[8739] = 25'b0000101000110011010010100;
    rom[8740] = 25'b0000100111111111110111111;
    rom[8741] = 25'b0000100111001100100110000;
    rom[8742] = 25'b0000100110011001011100111;
    rom[8743] = 25'b0000100101100110011100100;
    rom[8744] = 25'b0000100100110011100101000;
    rom[8745] = 25'b0000100100000000110110011;
    rom[8746] = 25'b0000100011001110010000101;
    rom[8747] = 25'b0000100010011011110011101;
    rom[8748] = 25'b0000100001101001011111111;
    rom[8749] = 25'b0000100000110111010101000;
    rom[8750] = 25'b0000100000000101010011001;
    rom[8751] = 25'b0000011111010011011010100;
    rom[8752] = 25'b0000011110100001101010111;
    rom[8753] = 25'b0000011101110000000100011;
    rom[8754] = 25'b0000011100111110100111000;
    rom[8755] = 25'b0000011100001101010011000;
    rom[8756] = 25'b0000011011011100001000010;
    rom[8757] = 25'b0000011010101011000110110;
    rom[8758] = 25'b0000011001111010001110100;
    rom[8759] = 25'b0000011001001001011111110;
    rom[8760] = 25'b0000011000011000111010010;
    rom[8761] = 25'b0000010111101000011110011;
    rom[8762] = 25'b0000010110111000001011111;
    rom[8763] = 25'b0000010110001000000010110;
    rom[8764] = 25'b0000010101011000000011011;
    rom[8765] = 25'b0000010100101000001101010;
    rom[8766] = 25'b0000010011111000100001000;
    rom[8767] = 25'b0000010011001000111110011;
    rom[8768] = 25'b0000010010011001100101011;
    rom[8769] = 25'b0000010001101010010110000;
    rom[8770] = 25'b0000010000111011010000011;
    rom[8771] = 25'b0000010000001100010100100;
    rom[8772] = 25'b0000001111011101100010100;
    rom[8773] = 25'b0000001110101110111010010;
    rom[8774] = 25'b0000001110000000011011111;
    rom[8775] = 25'b0000001101010010000111100;
    rom[8776] = 25'b0000001100100011111100111;
    rom[8777] = 25'b0000001011110101111100010;
    rom[8778] = 25'b0000001011001000000101100;
    rom[8779] = 25'b0000001010011010011001000;
    rom[8780] = 25'b0000001001101100110110011;
    rom[8781] = 25'b0000001000111111011101110;
    rom[8782] = 25'b0000001000010010001111100;
    rom[8783] = 25'b0000000111100101001011001;
    rom[8784] = 25'b0000000110111000010001000;
    rom[8785] = 25'b0000000110001011100001000;
    rom[8786] = 25'b0000000101011110111011001;
    rom[8787] = 25'b0000000100110010011111101;
    rom[8788] = 25'b0000000100000110001110011;
    rom[8789] = 25'b0000000011011010000111011;
    rom[8790] = 25'b0000000010101110001010110;
    rom[8791] = 25'b0000000010000010011000100;
    rom[8792] = 25'b0000000001010110110000100;
    rom[8793] = 25'b0000000000101011010011000;
    rom[8794] = 25'b0000000000000000000000000;
    rom[8795] = 25'b1111111111010100110111011;
    rom[8796] = 25'b1111111110101001111001001;
    rom[8797] = 25'b1111111101111111000101100;
    rom[8798] = 25'b1111111101010100011100011;
    rom[8799] = 25'b1111111100101001111101111;
    rom[8800] = 25'b1111111011111111101001111;
    rom[8801] = 25'b1111111011010101100000011;
    rom[8802] = 25'b1111111010101011100001101;
    rom[8803] = 25'b1111111010000001101101100;
    rom[8804] = 25'b1111111001011000000100001;
    rom[8805] = 25'b1111111000101110100101011;
    rom[8806] = 25'b1111111000000101010001010;
    rom[8807] = 25'b1111110111011100001000000;
    rom[8808] = 25'b1111110110110011001001100;
    rom[8809] = 25'b1111110110001010010101111;
    rom[8810] = 25'b1111110101100001101100111;
    rom[8811] = 25'b1111110100111001001111000;
    rom[8812] = 25'b1111110100010000111011110;
    rom[8813] = 25'b1111110011101000110011011;
    rom[8814] = 25'b1111110011000000110110000;
    rom[8815] = 25'b1111110010011001000011100;
    rom[8816] = 25'b1111110001110001011011111;
    rom[8817] = 25'b1111110001001001111111011;
    rom[8818] = 25'b1111110000100010101101110;
    rom[8819] = 25'b1111101111111011100111001;
    rom[8820] = 25'b1111101111010100101011100;
    rom[8821] = 25'b1111101110101101111011001;
    rom[8822] = 25'b1111101110000111010101101;
    rom[8823] = 25'b1111101101100000111011010;
    rom[8824] = 25'b1111101100111010101100000;
    rom[8825] = 25'b1111101100010100100111111;
    rom[8826] = 25'b1111101011101110101110110;
    rom[8827] = 25'b1111101011001001000000111;
    rom[8828] = 25'b1111101010100011011110010;
    rom[8829] = 25'b1111101001111110000110110;
    rom[8830] = 25'b1111101001011000111010011;
    rom[8831] = 25'b1111101000110011111001100;
    rom[8832] = 25'b1111101000001111000011101;
    rom[8833] = 25'b1111100111101010011001000;
    rom[8834] = 25'b1111100111000101111001110;
    rom[8835] = 25'b1111100110100001100101111;
    rom[8836] = 25'b1111100101111101011101010;
    rom[8837] = 25'b1111100101011001011111111;
    rom[8838] = 25'b1111100100110101101101110;
    rom[8839] = 25'b1111100100010010000111010;
    rom[8840] = 25'b1111100011101110101011111;
    rom[8841] = 25'b1111100011001011011100000;
    rom[8842] = 25'b1111100010101000010111101;
    rom[8843] = 25'b1111100010000101011110100;
    rom[8844] = 25'b1111100001100010110000111;
    rom[8845] = 25'b1111100001000000001110101;
    rom[8846] = 25'b1111100000011101110111111;
    rom[8847] = 25'b1111011111111011101100101;
    rom[8848] = 25'b1111011111011001101100110;
    rom[8849] = 25'b1111011110110111111000011;
    rom[8850] = 25'b1111011110010110001111110;
    rom[8851] = 25'b1111011101110100110010011;
    rom[8852] = 25'b1111011101010011100000101;
    rom[8853] = 25'b1111011100110010011010100;
    rom[8854] = 25'b1111011100010001011111110;
    rom[8855] = 25'b1111011011110000110000101;
    rom[8856] = 25'b1111011011010000001101001;
    rom[8857] = 25'b1111011010101111110101010;
    rom[8858] = 25'b1111011010001111101000111;
    rom[8859] = 25'b1111011001101111101000001;
    rom[8860] = 25'b1111011001001111110011000;
    rom[8861] = 25'b1111011000110000001001100;
    rom[8862] = 25'b1111011000010000101011101;
    rom[8863] = 25'b1111010111110001011001100;
    rom[8864] = 25'b1111010111010010010010111;
    rom[8865] = 25'b1111010110110011011000000;
    rom[8866] = 25'b1111010110010100101000110;
    rom[8867] = 25'b1111010101110110000101010;
    rom[8868] = 25'b1111010101010111101101011;
    rom[8869] = 25'b1111010100111001100001001;
    rom[8870] = 25'b1111010100011011100000110;
    rom[8871] = 25'b1111010011111101101100000;
    rom[8872] = 25'b1111010011100000000011000;
    rom[8873] = 25'b1111010011000010100101101;
    rom[8874] = 25'b1111010010100101010100001;
    rom[8875] = 25'b1111010010001000001110001;
    rom[8876] = 25'b1111010001101011010100001;
    rom[8877] = 25'b1111010001001110100101110;
    rom[8878] = 25'b1111010000110010000011001;
    rom[8879] = 25'b1111010000010101101100010;
    rom[8880] = 25'b1111001111111001100001001;
    rom[8881] = 25'b1111001111011101100001110;
    rom[8882] = 25'b1111001111000001101110010;
    rom[8883] = 25'b1111001110100110000110100;
    rom[8884] = 25'b1111001110001010101010011;
    rom[8885] = 25'b1111001101101111011010010;
    rom[8886] = 25'b1111001101010100010101110;
    rom[8887] = 25'b1111001100111001011101001;
    rom[8888] = 25'b1111001100011110110000010;
    rom[8889] = 25'b1111001100000100001111010;
    rom[8890] = 25'b1111001011101001111010000;
    rom[8891] = 25'b1111001011001111110000100;
    rom[8892] = 25'b1111001010110101110010111;
    rom[8893] = 25'b1111001010011100000001000;
    rom[8894] = 25'b1111001010000010011010111;
    rom[8895] = 25'b1111001001101001000000110;
    rom[8896] = 25'b1111001001001111110010010;
    rom[8897] = 25'b1111001000110110101111101;
    rom[8898] = 25'b1111001000011101111000111;
    rom[8899] = 25'b1111001000000101001101111;
    rom[8900] = 25'b1111000111101100101110101;
    rom[8901] = 25'b1111000111010100011011010;
    rom[8902] = 25'b1111000110111100010011101;
    rom[8903] = 25'b1111000110100100010111111;
    rom[8904] = 25'b1111000110001100100111111;
    rom[8905] = 25'b1111000101110101000011110;
    rom[8906] = 25'b1111000101011101101011011;
    rom[8907] = 25'b1111000101000110011110111;
    rom[8908] = 25'b1111000100101111011110001;
    rom[8909] = 25'b1111000100011000101001001;
    rom[8910] = 25'b1111000100000010000000000;
    rom[8911] = 25'b1111000011101011100010101;
    rom[8912] = 25'b1111000011010101010001001;
    rom[8913] = 25'b1111000010111111001011010;
    rom[8914] = 25'b1111000010101001010001011;
    rom[8915] = 25'b1111000010010011100011001;
    rom[8916] = 25'b1111000001111110000000101;
    rom[8917] = 25'b1111000001101000101010000;
    rom[8918] = 25'b1111000001010011011111001;
    rom[8919] = 25'b1111000000111110100000000;
    rom[8920] = 25'b1111000000101001101100101;
    rom[8921] = 25'b1111000000010101000101000;
    rom[8922] = 25'b1111000000000000101001001;
    rom[8923] = 25'b1110111111101100011001001;
    rom[8924] = 25'b1110111111011000010100110;
    rom[8925] = 25'b1110111111000100011100001;
    rom[8926] = 25'b1110111110110000101111001;
    rom[8927] = 25'b1110111110011101001110000;
    rom[8928] = 25'b1110111110001001111000100;
    rom[8929] = 25'b1110111101110110101110101;
    rom[8930] = 25'b1110111101100011110000110;
    rom[8931] = 25'b1110111101010000111110011;
    rom[8932] = 25'b1110111100111110010111101;
    rom[8933] = 25'b1110111100101011111100101;
    rom[8934] = 25'b1110111100011001101101010;
    rom[8935] = 25'b1110111100000111101001101;
    rom[8936] = 25'b1110111011110101110001100;
    rom[8937] = 25'b1110111011100100000101010;
    rom[8938] = 25'b1110111011010010100100100;
    rom[8939] = 25'b1110111011000001001111011;
    rom[8940] = 25'b1110111010110000000101111;
    rom[8941] = 25'b1110111010011111001000000;
    rom[8942] = 25'b1110111010001110010101110;
    rom[8943] = 25'b1110111001111101101111000;
    rom[8944] = 25'b1110111001101101010011111;
    rom[8945] = 25'b1110111001011101000100011;
    rom[8946] = 25'b1110111001001101000000100;
    rom[8947] = 25'b1110111000111101001000000;
    rom[8948] = 25'b1110111000101101011011001;
    rom[8949] = 25'b1110111000011101111001110;
    rom[8950] = 25'b1110111000001110100011111;
    rom[8951] = 25'b1110110111111111011001100;
    rom[8952] = 25'b1110110111110000011010110;
    rom[8953] = 25'b1110110111100001100111010;
    rom[8954] = 25'b1110110111010010111111011;
    rom[8955] = 25'b1110110111000100100010111;
    rom[8956] = 25'b1110110110110110010001111;
    rom[8957] = 25'b1110110110101000001100010;
    rom[8958] = 25'b1110110110011010010010001;
    rom[8959] = 25'b1110110110001100100011011;
    rom[8960] = 25'b1110110101111110111111111;
    rom[8961] = 25'b1110110101110001100111111;
    rom[8962] = 25'b1110110101100100011011010;
    rom[8963] = 25'b1110110101010111011010000;
    rom[8964] = 25'b1110110101001010100100000;
    rom[8965] = 25'b1110110100111101111001011;
    rom[8966] = 25'b1110110100110001011010000;
    rom[8967] = 25'b1110110100100101000101111;
    rom[8968] = 25'b1110110100011000111101000;
    rom[8969] = 25'b1110110100001100111111100;
    rom[8970] = 25'b1110110100000001001101010;
    rom[8971] = 25'b1110110011110101100110001;
    rom[8972] = 25'b1110110011101010001010010;
    rom[8973] = 25'b1110110011011110111001100;
    rom[8974] = 25'b1110110011010011110100000;
    rom[8975] = 25'b1110110011001000111001101;
    rom[8976] = 25'b1110110010111110001010100;
    rom[8977] = 25'b1110110010110011100110011;
    rom[8978] = 25'b1110110010101001001101011;
    rom[8979] = 25'b1110110010011110111111100;
    rom[8980] = 25'b1110110010010100111100110;
    rom[8981] = 25'b1110110010001011000100111;
    rom[8982] = 25'b1110110010000001011000001;
    rom[8983] = 25'b1110110001110111110110100;
    rom[8984] = 25'b1110110001101110011111111;
    rom[8985] = 25'b1110110001100101010100000;
    rom[8986] = 25'b1110110001011100010011010;
    rom[8987] = 25'b1110110001010011011101100;
    rom[8988] = 25'b1110110001001010110010100;
    rom[8989] = 25'b1110110001000010010010100;
    rom[8990] = 25'b1110110000111001111101011;
    rom[8991] = 25'b1110110000110001110011001;
    rom[8992] = 25'b1110110000101001110011110;
    rom[8993] = 25'b1110110000100001111111001;
    rom[8994] = 25'b1110110000011010010101011;
    rom[8995] = 25'b1110110000010010110110011;
    rom[8996] = 25'b1110110000001011100010001;
    rom[8997] = 25'b1110110000000100011000101;
    rom[8998] = 25'b1110101111111101011001111;
    rom[8999] = 25'b1110101111110110100101110;
    rom[9000] = 25'b1110101111101111111100011;
    rom[9001] = 25'b1110101111101001011101101;
    rom[9002] = 25'b1110101111100011001001100;
    rom[9003] = 25'b1110101111011101000000000;
    rom[9004] = 25'b1110101111010111000001001;
    rom[9005] = 25'b1110101111010001001100101;
    rom[9006] = 25'b1110101111001011100010111;
    rom[9007] = 25'b1110101111000110000011101;
    rom[9008] = 25'b1110101111000000101110110;
    rom[9009] = 25'b1110101110111011100100100;
    rom[9010] = 25'b1110101110110110100100101;
    rom[9011] = 25'b1110101110110001101111010;
    rom[9012] = 25'b1110101110101101000100001;
    rom[9013] = 25'b1110101110101000100011100;
    rom[9014] = 25'b1110101110100100001101010;
    rom[9015] = 25'b1110101110100000000001010;
    rom[9016] = 25'b1110101110011011111111100;
    rom[9017] = 25'b1110101110011000001000010;
    rom[9018] = 25'b1110101110010100011011000;
    rom[9019] = 25'b1110101110010000111000001;
    rom[9020] = 25'b1110101110001101011111100;
    rom[9021] = 25'b1110101110001010010000111;
    rom[9022] = 25'b1110101110000111001100101;
    rom[9023] = 25'b1110101110000100010010011;
    rom[9024] = 25'b1110101110000001100010010;
    rom[9025] = 25'b1110101101111110111100010;
    rom[9026] = 25'b1110101101111100100000010;
    rom[9027] = 25'b1110101101111010001110011;
    rom[9028] = 25'b1110101101111000000110011;
    rom[9029] = 25'b1110101101110110001000011;
    rom[9030] = 25'b1110101101110100010100011;
    rom[9031] = 25'b1110101101110010101010010;
    rom[9032] = 25'b1110101101110001001010000;
    rom[9033] = 25'b1110101101101111110011110;
    rom[9034] = 25'b1110101101101110100111010;
    rom[9035] = 25'b1110101101101101100100100;
    rom[9036] = 25'b1110101101101100101011101;
    rom[9037] = 25'b1110101101101011111100011;
    rom[9038] = 25'b1110101101101011010111000;
    rom[9039] = 25'b1110101101101010111011010;
    rom[9040] = 25'b1110101101101010101001001;
    rom[9041] = 25'b1110101101101010100000110;
    rom[9042] = 25'b1110101101101010100010000;
    rom[9043] = 25'b1110101101101010101100110;
    rom[9044] = 25'b1110101101101011000001001;
    rom[9045] = 25'b1110101101101011011111000;
    rom[9046] = 25'b1110101101101100000110011;
    rom[9047] = 25'b1110101101101100110111010;
    rom[9048] = 25'b1110101101101101110001100;
    rom[9049] = 25'b1110101101101110110101010;
    rom[9050] = 25'b1110101101110000000010010;
    rom[9051] = 25'b1110101101110001011000110;
    rom[9052] = 25'b1110101101110010111000011;
    rom[9053] = 25'b1110101101110100100001011;
    rom[9054] = 25'b1110101101110110010011110;
    rom[9055] = 25'b1110101101111000001111010;
    rom[9056] = 25'b1110101101111010010011111;
    rom[9057] = 25'b1110101101111100100001111;
    rom[9058] = 25'b1110101101111110111000111;
    rom[9059] = 25'b1110101110000001011001000;
    rom[9060] = 25'b1110101110000100000010001;
    rom[9061] = 25'b1110101110000110110100100;
    rom[9062] = 25'b1110101110001001101111101;
    rom[9063] = 25'b1110101110001100110011111;
    rom[9064] = 25'b1110101110010000000001001;
    rom[9065] = 25'b1110101110010011010111010;
    rom[9066] = 25'b1110101110010110110110010;
    rom[9067] = 25'b1110101110011010011110001;
    rom[9068] = 25'b1110101110011110001110110;
    rom[9069] = 25'b1110101110100010001000010;
    rom[9070] = 25'b1110101110100110001010100;
    rom[9071] = 25'b1110101110101010010101011;
    rom[9072] = 25'b1110101110101110101001000;
    rom[9073] = 25'b1110101110110011000101010;
    rom[9074] = 25'b1110101110110111101010001;
    rom[9075] = 25'b1110101110111100010111110;
    rom[9076] = 25'b1110101111000001001101110;
    rom[9077] = 25'b1110101111000110001100011;
    rom[9078] = 25'b1110101111001011010011100;
    rom[9079] = 25'b1110101111010000100011000;
    rom[9080] = 25'b1110101111010101111010111;
    rom[9081] = 25'b1110101111011011011011011;
    rom[9082] = 25'b1110101111100001000100001;
    rom[9083] = 25'b1110101111100110110101001;
    rom[9084] = 25'b1110101111101100101110011;
    rom[9085] = 25'b1110101111110010110000000;
    rom[9086] = 25'b1110101111111000111001111;
    rom[9087] = 25'b1110101111111111001011111;
    rom[9088] = 25'b1110110000000101100110000;
    rom[9089] = 25'b1110110000001100001000010;
    rom[9090] = 25'b1110110000010010110010101;
    rom[9091] = 25'b1110110000011001100101000;
    rom[9092] = 25'b1110110000100000011111011;
    rom[9093] = 25'b1110110000100111100001111;
    rom[9094] = 25'b1110110000101110101100001;
    rom[9095] = 25'b1110110000110101111110011;
    rom[9096] = 25'b1110110000111101011000101;
    rom[9097] = 25'b1110110001000100111010100;
    rom[9098] = 25'b1110110001001100100100010;
    rom[9099] = 25'b1110110001010100010101111;
    rom[9100] = 25'b1110110001011100001111000;
    rom[9101] = 25'b1110110001100100010000000;
    rom[9102] = 25'b1110110001101100011000110;
    rom[9103] = 25'b1110110001110100101000111;
    rom[9104] = 25'b1110110001111101000000101;
    rom[9105] = 25'b1110110010000101100000001;
    rom[9106] = 25'b1110110010001110000111000;
    rom[9107] = 25'b1110110010010110110101011;
    rom[9108] = 25'b1110110010011111101011010;
    rom[9109] = 25'b1110110010101000101000011;
    rom[9110] = 25'b1110110010110001101101000;
    rom[9111] = 25'b1110110010111010111000111;
    rom[9112] = 25'b1110110011000100001100001;
    rom[9113] = 25'b1110110011001101100110101;
    rom[9114] = 25'b1110110011010111001000011;
    rom[9115] = 25'b1110110011100000110001010;
    rom[9116] = 25'b1110110011101010100001010;
    rom[9117] = 25'b1110110011110100011000011;
    rom[9118] = 25'b1110110011111110010110101;
    rom[9119] = 25'b1110110100001000011011111;
    rom[9120] = 25'b1110110100010010101000001;
    rom[9121] = 25'b1110110100011100111011011;
    rom[9122] = 25'b1110110100100111010101100;
    rom[9123] = 25'b1110110100110001110110101;
    rom[9124] = 25'b1110110100111100011110011;
    rom[9125] = 25'b1110110101000111001101001;
    rom[9126] = 25'b1110110101010010000010101;
    rom[9127] = 25'b1110110101011100111110110;
    rom[9128] = 25'b1110110101101000000001101;
    rom[9129] = 25'b1110110101110011001011001;
    rom[9130] = 25'b1110110101111110011011011;
    rom[9131] = 25'b1110110110001001110010001;
    rom[9132] = 25'b1110110110010101001111100;
    rom[9133] = 25'b1110110110100000110011010;
    rom[9134] = 25'b1110110110101100011101101;
    rom[9135] = 25'b1110110110111000001110010;
    rom[9136] = 25'b1110110111000100000101011;
    rom[9137] = 25'b1110110111010000000010110;
    rom[9138] = 25'b1110110111011100000110101;
    rom[9139] = 25'b1110110111101000010000101;
    rom[9140] = 25'b1110110111110100100000111;
    rom[9141] = 25'b1110111000000000110111011;
    rom[9142] = 25'b1110111000001101010100000;
    rom[9143] = 25'b1110111000011001110110110;
    rom[9144] = 25'b1110111000100110011111101;
    rom[9145] = 25'b1110111000110011001110100;
    rom[9146] = 25'b1110111001000000000011011;
    rom[9147] = 25'b1110111001001100111110011;
    rom[9148] = 25'b1110111001011001111111001;
    rom[9149] = 25'b1110111001100111000101110;
    rom[9150] = 25'b1110111001110100010010010;
    rom[9151] = 25'b1110111010000001100100101;
    rom[9152] = 25'b1110111010001110111100110;
    rom[9153] = 25'b1110111010011100011010100;
    rom[9154] = 25'b1110111010101001111110000;
    rom[9155] = 25'b1110111010110111100111010;
    rom[9156] = 25'b1110111011000101010110000;
    rom[9157] = 25'b1110111011010011001010011;
    rom[9158] = 25'b1110111011100001000100010;
    rom[9159] = 25'b1110111011101111000011101;
    rom[9160] = 25'b1110111011111101001000011;
    rom[9161] = 25'b1110111100001011010010110;
    rom[9162] = 25'b1110111100011001100010011;
    rom[9163] = 25'b1110111100100111110111010;
    rom[9164] = 25'b1110111100110110010001100;
    rom[9165] = 25'b1110111101000100110001000;
    rom[9166] = 25'b1110111101010011010101110;
    rom[9167] = 25'b1110111101100001111111110;
    rom[9168] = 25'b1110111101110000101110101;
    rom[9169] = 25'b1110111101111111100010111;
    rom[9170] = 25'b1110111110001110011100001;
    rom[9171] = 25'b1110111110011101011010010;
    rom[9172] = 25'b1110111110101100011101100;
    rom[9173] = 25'b1110111110111011100101100;
    rom[9174] = 25'b1110111111001010110010101;
    rom[9175] = 25'b1110111111011010000100100;
    rom[9176] = 25'b1110111111101001011011001;
    rom[9177] = 25'b1110111111111000110110101;
    rom[9178] = 25'b1111000000001000010110111;
    rom[9179] = 25'b1111000000010111111011110;
    rom[9180] = 25'b1111000000100111100101011;
    rom[9181] = 25'b1111000000110111010011100;
    rom[9182] = 25'b1111000001000111000110010;
    rom[9183] = 25'b1111000001010110111101101;
    rom[9184] = 25'b1111000001100110111001011;
    rom[9185] = 25'b1111000001110110111001101;
    rom[9186] = 25'b1111000010000110111110010;
    rom[9187] = 25'b1111000010010111000111011;
    rom[9188] = 25'b1111000010100111010100110;
    rom[9189] = 25'b1111000010110111100110011;
    rom[9190] = 25'b1111000011000111111100010;
    rom[9191] = 25'b1111000011011000010110100;
    rom[9192] = 25'b1111000011101000110100111;
    rom[9193] = 25'b1111000011111001010111010;
    rom[9194] = 25'b1111000100001001111101110;
    rom[9195] = 25'b1111000100011010101000011;
    rom[9196] = 25'b1111000100101011010111001;
    rom[9197] = 25'b1111000100111100001001101;
    rom[9198] = 25'b1111000101001101000000010;
    rom[9199] = 25'b1111000101011101111010101;
    rom[9200] = 25'b1111000101101110111000111;
    rom[9201] = 25'b1111000101111111111011000;
    rom[9202] = 25'b1111000110010001000000111;
    rom[9203] = 25'b1111000110100010001010100;
    rom[9204] = 25'b1111000110110011010111111;
    rom[9205] = 25'b1111000111000100101000110;
    rom[9206] = 25'b1111000111010101111101011;
    rom[9207] = 25'b1111000111100111010101100;
    rom[9208] = 25'b1111000111111000110001001;
    rom[9209] = 25'b1111001000001010010000011;
    rom[9210] = 25'b1111001000011011110010111;
    rom[9211] = 25'b1111001000101101011001000;
    rom[9212] = 25'b1111001000111111000010100;
    rom[9213] = 25'b1111001001010000101111010;
    rom[9214] = 25'b1111001001100010011111010;
    rom[9215] = 25'b1111001001110100010010100;
    rom[9216] = 25'b1111001010000110001001000;
    rom[9217] = 25'b1111001010011000000010101;
    rom[9218] = 25'b1111001010101001111111100;
    rom[9219] = 25'b1111001010111011111111100;
    rom[9220] = 25'b1111001011001110000010011;
    rom[9221] = 25'b1111001011100000001000011;
    rom[9222] = 25'b1111001011110010010001011;
    rom[9223] = 25'b1111001100000100011101010;
    rom[9224] = 25'b1111001100010110101100000;
    rom[9225] = 25'b1111001100101000111101101;
    rom[9226] = 25'b1111001100111011010010001;
    rom[9227] = 25'b1111001101001101101001011;
    rom[9228] = 25'b1111001101100000000011010;
    rom[9229] = 25'b1111001101110010011111111;
    rom[9230] = 25'b1111001110000100111111010;
    rom[9231] = 25'b1111001110010111100001001;
    rom[9232] = 25'b1111001110101010000101110;
    rom[9233] = 25'b1111001110111100101100110;
    rom[9234] = 25'b1111001111001111010110011;
    rom[9235] = 25'b1111001111100010000010011;
    rom[9236] = 25'b1111001111110100110000101;
    rom[9237] = 25'b1111010000000111100001101;
    rom[9238] = 25'b1111010000011010010100110;
    rom[9239] = 25'b1111010000101101001010001;
    rom[9240] = 25'b1111010001000000000001111;
    rom[9241] = 25'b1111010001010010111011111;
    rom[9242] = 25'b1111010001100101110111111;
    rom[9243] = 25'b1111010001111000110110010;
    rom[9244] = 25'b1111010010001011110110100;
    rom[9245] = 25'b1111010010011110111001000;
    rom[9246] = 25'b1111010010110001111101100;
    rom[9247] = 25'b1111010011000101000011111;
    rom[9248] = 25'b1111010011011000001100011;
    rom[9249] = 25'b1111010011101011010110101;
    rom[9250] = 25'b1111010011111110100010111;
    rom[9251] = 25'b1111010100010001110000111;
    rom[9252] = 25'b1111010100100101000000110;
    rom[9253] = 25'b1111010100111000010010011;
    rom[9254] = 25'b1111010101001011100101101;
    rom[9255] = 25'b1111010101011110111010101;
    rom[9256] = 25'b1111010101110010010001010;
    rom[9257] = 25'b1111010110000101101001100;
    rom[9258] = 25'b1111010110011001000011010;
    rom[9259] = 25'b1111010110101100011110101;
    rom[9260] = 25'b1111010110111111111011011;
    rom[9261] = 25'b1111010111010011011001101;
    rom[9262] = 25'b1111010111100110111001010;
    rom[9263] = 25'b1111010111111010011010011;
    rom[9264] = 25'b1111011000001101111100110;
    rom[9265] = 25'b1111011000100001100000011;
    rom[9266] = 25'b1111011000110101000101010;
    rom[9267] = 25'b1111011001001000101011100;
    rom[9268] = 25'b1111011001011100010010111;
    rom[9269] = 25'b1111011001101111111011010;
    rom[9270] = 25'b1111011010000011100101000;
    rom[9271] = 25'b1111011010010111001111101;
    rom[9272] = 25'b1111011010101010111011010;
    rom[9273] = 25'b1111011010111110101000000;
    rom[9274] = 25'b1111011011010010010101101;
    rom[9275] = 25'b1111011011100110000100010;
    rom[9276] = 25'b1111011011111001110011110;
    rom[9277] = 25'b1111011100001101100100000;
    rom[9278] = 25'b1111011100100001010101010;
    rom[9279] = 25'b1111011100110101000111001;
    rom[9280] = 25'b1111011101001000111001110;
    rom[9281] = 25'b1111011101011100101101000;
    rom[9282] = 25'b1111011101110000100001000;
    rom[9283] = 25'b1111011110000100010101101;
    rom[9284] = 25'b1111011110011000001010111;
    rom[9285] = 25'b1111011110101100000000110;
    rom[9286] = 25'b1111011110111111110111000;
    rom[9287] = 25'b1111011111010011101101110;
    rom[9288] = 25'b1111011111100111100101000;
    rom[9289] = 25'b1111011111111011011100101;
    rom[9290] = 25'b1111100000001111010100101;
    rom[9291] = 25'b1111100000100011001101000;
    rom[9292] = 25'b1111100000110111000101101;
    rom[9293] = 25'b1111100001001010111110100;
    rom[9294] = 25'b1111100001011110110111101;
    rom[9295] = 25'b1111100001110010110000111;
    rom[9296] = 25'b1111100010000110101010011;
    rom[9297] = 25'b1111100010011010100011111;
    rom[9298] = 25'b1111100010101110011101101;
    rom[9299] = 25'b1111100011000010010111011;
    rom[9300] = 25'b1111100011010110010001001;
    rom[9301] = 25'b1111100011101010001010111;
    rom[9302] = 25'b1111100011111110000100100;
    rom[9303] = 25'b1111100100010001111110000;
    rom[9304] = 25'b1111100100100101110111101;
    rom[9305] = 25'b1111100100111001110000111;
    rom[9306] = 25'b1111100101001101101010000;
    rom[9307] = 25'b1111100101100001100010111;
    rom[9308] = 25'b1111100101110101011011011;
    rom[9309] = 25'b1111100110001001010011110;
    rom[9310] = 25'b1111100110011101001011101;
    rom[9311] = 25'b1111100110110001000011010;
    rom[9312] = 25'b1111100111000100111010100;
    rom[9313] = 25'b1111100111011000110001010;
    rom[9314] = 25'b1111100111101100100111101;
    rom[9315] = 25'b1111101000000000011101011;
    rom[9316] = 25'b1111101000010100010010101;
    rom[9317] = 25'b1111101000101000000111010;
    rom[9318] = 25'b1111101000111011111011011;
    rom[9319] = 25'b1111101001001111101110111;
    rom[9320] = 25'b1111101001100011100001101;
    rom[9321] = 25'b1111101001110111010011110;
    rom[9322] = 25'b1111101010001011000101001;
    rom[9323] = 25'b1111101010011110110101100;
    rom[9324] = 25'b1111101010110010100101011;
    rom[9325] = 25'b1111101011000110010100010;
    rom[9326] = 25'b1111101011011010000010010;
    rom[9327] = 25'b1111101011101101101111100;
    rom[9328] = 25'b1111101100000001011011110;
    rom[9329] = 25'b1111101100010101000110111;
    rom[9330] = 25'b1111101100101000110001001;
    rom[9331] = 25'b1111101100111100011010011;
    rom[9332] = 25'b1111101101010000000010100;
    rom[9333] = 25'b1111101101100011101001101;
    rom[9334] = 25'b1111101101110111001111100;
    rom[9335] = 25'b1111101110001010110100010;
    rom[9336] = 25'b1111101110011110010111111;
    rom[9337] = 25'b1111101110110001111010010;
    rom[9338] = 25'b1111101111000101011011010;
    rom[9339] = 25'b1111101111011000111011001;
    rom[9340] = 25'b1111101111101100011001101;
    rom[9341] = 25'b1111101111111111110110110;
    rom[9342] = 25'b1111110000010011010010100;
    rom[9343] = 25'b1111110000100110101100111;
    rom[9344] = 25'b1111110000111010000101110;
    rom[9345] = 25'b1111110001001101011101010;
    rom[9346] = 25'b1111110001100000110011010;
    rom[9347] = 25'b1111110001110100000111100;
    rom[9348] = 25'b1111110010000111011010011;
    rom[9349] = 25'b1111110010011010101011101;
    rom[9350] = 25'b1111110010101101111011010;
    rom[9351] = 25'b1111110011000001001001010;
    rom[9352] = 25'b1111110011010100010101100;
    rom[9353] = 25'b1111110011100111100000000;
    rom[9354] = 25'b1111110011111010101000111;
    rom[9355] = 25'b1111110100001101110000000;
    rom[9356] = 25'b1111110100100000110101010;
    rom[9357] = 25'b1111110100110011111000110;
    rom[9358] = 25'b1111110101000110111010010;
    rom[9359] = 25'b1111110101011001111001111;
    rom[9360] = 25'b1111110101101100110111101;
    rom[9361] = 25'b1111110101111111110011100;
    rom[9362] = 25'b1111110110010010101101011;
    rom[9363] = 25'b1111110110100101100101001;
    rom[9364] = 25'b1111110110111000011011000;
    rom[9365] = 25'b1111110111001011001110110;
    rom[9366] = 25'b1111110111011110000000011;
    rom[9367] = 25'b1111110111110000101111111;
    rom[9368] = 25'b1111111000000011011101010;
    rom[9369] = 25'b1111111000010110001000100;
    rom[9370] = 25'b1111111000101000110001100;
    rom[9371] = 25'b1111111000111011011000010;
    rom[9372] = 25'b1111111001001101111100110;
    rom[9373] = 25'b1111111001100000011111000;
    rom[9374] = 25'b1111111001110010111111000;
    rom[9375] = 25'b1111111010000101011100100;
    rom[9376] = 25'b1111111010010111110111110;
    rom[9377] = 25'b1111111010101010010000101;
    rom[9378] = 25'b1111111010111100100111001;
    rom[9379] = 25'b1111111011001110111011000;
    rom[9380] = 25'b1111111011100001001100101;
    rom[9381] = 25'b1111111011110011011011101;
    rom[9382] = 25'b1111111100000101101000001;
    rom[9383] = 25'b1111111100010111110010000;
    rom[9384] = 25'b1111111100101001111001100;
    rom[9385] = 25'b1111111100111011111110010;
    rom[9386] = 25'b1111111101001110000000011;
    rom[9387] = 25'b1111111101011111111111111;
    rom[9388] = 25'b1111111101110001111100101;
    rom[9389] = 25'b1111111110000011110110110;
    rom[9390] = 25'b1111111110010101101110001;
    rom[9391] = 25'b1111111110100111100010111;
    rom[9392] = 25'b1111111110111001010100110;
    rom[9393] = 25'b1111111111001011000011110;
    rom[9394] = 25'b1111111111011100110000001;
    rom[9395] = 25'b1111111111101110011001100;
    rom[9396] = 25'b0000000000000000000000000;
    rom[9397] = 25'b0000000000010001100011100;
    rom[9398] = 25'b0000000000100011000100010;
    rom[9399] = 25'b0000000000110100100010000;
    rom[9400] = 25'b0000000001000101111100110;
    rom[9401] = 25'b0000000001010111010100100;
    rom[9402] = 25'b0000000001101000101001011;
    rom[9403] = 25'b0000000001111001111011001;
    rom[9404] = 25'b0000000010001011001001111;
    rom[9405] = 25'b0000000010011100010101011;
    rom[9406] = 25'b0000000010101101011101111;
    rom[9407] = 25'b0000000010111110100011010;
    rom[9408] = 25'b0000000011001111100101100;
    rom[9409] = 25'b0000000011100000100100100;
    rom[9410] = 25'b0000000011110001100000011;
    rom[9411] = 25'b0000000100000010011000111;
    rom[9412] = 25'b0000000100010011001110010;
    rom[9413] = 25'b0000000100100100000000100;
    rom[9414] = 25'b0000000100110100101111010;
    rom[9415] = 25'b0000000101000101011010110;
    rom[9416] = 25'b0000000101010110000010111;
    rom[9417] = 25'b0000000101100110100111110;
    rom[9418] = 25'b0000000101110111001001010;
    rom[9419] = 25'b0000000110000111100111011;
    rom[9420] = 25'b0000000110011000000010000;
    rom[9421] = 25'b0000000110101000011001010;
    rom[9422] = 25'b0000000110111000101101000;
    rom[9423] = 25'b0000000111001000111101011;
    rom[9424] = 25'b0000000111011001001010001;
    rom[9425] = 25'b0000000111101001010011100;
    rom[9426] = 25'b0000000111111001011001010;
    rom[9427] = 25'b0000001000001001011011100;
    rom[9428] = 25'b0000001000011001011010001;
    rom[9429] = 25'b0000001000101001010101001;
    rom[9430] = 25'b0000001000111001001100101;
    rom[9431] = 25'b0000001001001001000000011;
    rom[9432] = 25'b0000001001011000110000100;
    rom[9433] = 25'b0000001001101000011101000;
    rom[9434] = 25'b0000001001111000000101110;
    rom[9435] = 25'b0000001010000111101010111;
    rom[9436] = 25'b0000001010010111001100010;
    rom[9437] = 25'b0000001010100110101001110;
    rom[9438] = 25'b0000001010110110000011101;
    rom[9439] = 25'b0000001011000101011001110;
    rom[9440] = 25'b0000001011010100101100000;
    rom[9441] = 25'b0000001011100011111010100;
    rom[9442] = 25'b0000001011110011000101001;
    rom[9443] = 25'b0000001100000010001011111;
    rom[9444] = 25'b0000001100010001001110110;
    rom[9445] = 25'b0000001100100000001101110;
    rom[9446] = 25'b0000001100101111001000111;
    rom[9447] = 25'b0000001100111110000000001;
    rom[9448] = 25'b0000001101001100110011011;
    rom[9449] = 25'b0000001101011011100010101;
    rom[9450] = 25'b0000001101101010001110000;
    rom[9451] = 25'b0000001101111000110101010;
    rom[9452] = 25'b0000001110000111011000110;
    rom[9453] = 25'b0000001110010101111000000;
    rom[9454] = 25'b0000001110100100010011010;
    rom[9455] = 25'b0000001110110010101010100;
    rom[9456] = 25'b0000001111000000111101110;
    rom[9457] = 25'b0000001111001111001100111;
    rom[9458] = 25'b0000001111011101010111111;
    rom[9459] = 25'b0000001111101011011110110;
    rom[9460] = 25'b0000001111111001100001100;
    rom[9461] = 25'b0000010000000111100000001;
    rom[9462] = 25'b0000010000010101011010101;
    rom[9463] = 25'b0000010000100011010000111;
    rom[9464] = 25'b0000010000110001000011000;
    rom[9465] = 25'b0000010000111110110000111;
    rom[9466] = 25'b0000010001001100011010110;
    rom[9467] = 25'b0000010001011010000000001;
    rom[9468] = 25'b0000010001100111100001011;
    rom[9469] = 25'b0000010001110100111110011;
    rom[9470] = 25'b0000010010000010010111001;
    rom[9471] = 25'b0000010010001111101011101;
    rom[9472] = 25'b0000010010011100111011110;
    rom[9473] = 25'b0000010010101010000111101;
    rom[9474] = 25'b0000010010110111001111001;
    rom[9475] = 25'b0000010011000100010010010;
    rom[9476] = 25'b0000010011010001010001001;
    rom[9477] = 25'b0000010011011110001011101;
    rom[9478] = 25'b0000010011101011000001110;
    rom[9479] = 25'b0000010011110111110011100;
    rom[9480] = 25'b0000010100000100100000111;
    rom[9481] = 25'b0000010100010001001001110;
    rom[9482] = 25'b0000010100011101101110011;
    rom[9483] = 25'b0000010100101010001110100;
    rom[9484] = 25'b0000010100110110101010001;
    rom[9485] = 25'b0000010101000011000001010;
    rom[9486] = 25'b0000010101001111010100001;
    rom[9487] = 25'b0000010101011011100010011;
    rom[9488] = 25'b0000010101100111101100001;
    rom[9489] = 25'b0000010101110011110001100;
    rom[9490] = 25'b0000010101111111110010010;
    rom[9491] = 25'b0000010110001011101110100;
    rom[9492] = 25'b0000010110010111100110010;
    rom[9493] = 25'b0000010110100011011001100;
    rom[9494] = 25'b0000010110101111001000010;
    rom[9495] = 25'b0000010110111010110010010;
    rom[9496] = 25'b0000010111000110010111111;
    rom[9497] = 25'b0000010111010001111000111;
    rom[9498] = 25'b0000010111011101010101010;
    rom[9499] = 25'b0000010111101000101101001;
    rom[9500] = 25'b0000010111110100000000010;
    rom[9501] = 25'b0000010111111111001110111;
    rom[9502] = 25'b0000011000001010011000111;
    rom[9503] = 25'b0000011000010101011110010;
    rom[9504] = 25'b0000011000100000011111000;
    rom[9505] = 25'b0000011000101011011011000;
    rom[9506] = 25'b0000011000110110010010011;
    rom[9507] = 25'b0000011001000001000101010;
    rom[9508] = 25'b0000011001001011110011010;
    rom[9509] = 25'b0000011001010110011100110;
    rom[9510] = 25'b0000011001100001000001100;
    rom[9511] = 25'b0000011001101011100001100;
    rom[9512] = 25'b0000011001110101111100111;
    rom[9513] = 25'b0000011010000000010011100;
    rom[9514] = 25'b0000011010001010100101011;
    rom[9515] = 25'b0000011010010100110010110;
    rom[9516] = 25'b0000011010011110111011001;
    rom[9517] = 25'b0000011010101000111111000;
    rom[9518] = 25'b0000011010110010111110000;
    rom[9519] = 25'b0000011010111100111000010;
    rom[9520] = 25'b0000011011000110101101111;
    rom[9521] = 25'b0000011011010000011110101;
    rom[9522] = 25'b0000011011011010001010101;
    rom[9523] = 25'b0000011011100011110001111;
    rom[9524] = 25'b0000011011101101010100011;
    rom[9525] = 25'b0000011011110110110010001;
    rom[9526] = 25'b0000011100000000001011000;
    rom[9527] = 25'b0000011100001001011111001;
    rom[9528] = 25'b0000011100010010101110100;
    rom[9529] = 25'b0000011100011011111001000;
    rom[9530] = 25'b0000011100100100111110110;
    rom[9531] = 25'b0000011100101101111111110;
    rom[9532] = 25'b0000011100110110111011111;
    rom[9533] = 25'b0000011100111111110011001;
    rom[9534] = 25'b0000011101001000100101101;
    rom[9535] = 25'b0000011101010001010011011;
    rom[9536] = 25'b0000011101011001111100001;
    rom[9537] = 25'b0000011101100010100000010;
    rom[9538] = 25'b0000011101101010111111011;
    rom[9539] = 25'b0000011101110011011001110;
    rom[9540] = 25'b0000011101111011101111010;
    rom[9541] = 25'b0000011110000011111111111;
    rom[9542] = 25'b0000011110001100001011110;
    rom[9543] = 25'b0000011110010100010010110;
    rom[9544] = 25'b0000011110011100010100111;
    rom[9545] = 25'b0000011110100100010010001;
    rom[9546] = 25'b0000011110101100001010100;
    rom[9547] = 25'b0000011110110011111110001;
    rom[9548] = 25'b0000011110111011101100111;
    rom[9549] = 25'b0000011111000011010110101;
    rom[9550] = 25'b0000011111001010111011101;
    rom[9551] = 25'b0000011111010010011011110;
    rom[9552] = 25'b0000011111011001110111000;
    rom[9553] = 25'b0000011111100001001101011;
    rom[9554] = 25'b0000011111101000011111000;
    rom[9555] = 25'b0000011111101111101011100;
    rom[9556] = 25'b0000011111110110110011011;
    rom[9557] = 25'b0000011111111101110110010;
    rom[9558] = 25'b0000100000000100110100010;
    rom[9559] = 25'b0000100000001011101101011;
    rom[9560] = 25'b0000100000010010100001110;
    rom[9561] = 25'b0000100000011001010001001;
    rom[9562] = 25'b0000100000011111111011101;
    rom[9563] = 25'b0000100000100110100001010;
    rom[9564] = 25'b0000100000101101000010001;
    rom[9565] = 25'b0000100000110011011110000;
    rom[9566] = 25'b0000100000111001110101000;
    rom[9567] = 25'b0000100001000000000111010;
    rom[9568] = 25'b0000100001000110010100100;
    rom[9569] = 25'b0000100001001100011100111;
    rom[9570] = 25'b0000100001010010100000100;
    rom[9571] = 25'b0000100001011000011111010;
    rom[9572] = 25'b0000100001011110011001001;
    rom[9573] = 25'b0000100001100100001110000;
    rom[9574] = 25'b0000100001101001111110001;
    rom[9575] = 25'b0000100001101111101001011;
    rom[9576] = 25'b0000100001110101001111110;
    rom[9577] = 25'b0000100001111010110001010;
    rom[9578] = 25'b0000100010000000001101111;
    rom[9579] = 25'b0000100010000101100101110;
    rom[9580] = 25'b0000100010001010111000101;
    rom[9581] = 25'b0000100010010000000110110;
    rom[9582] = 25'b0000100010010101010000000;
    rom[9583] = 25'b0000100010011010010100100;
    rom[9584] = 25'b0000100010011111010100001;
    rom[9585] = 25'b0000100010100100001110110;
    rom[9586] = 25'b0000100010101001000100101;
    rom[9587] = 25'b0000100010101101110101110;
    rom[9588] = 25'b0000100010110010100010000;
    rom[9589] = 25'b0000100010110111001001100;
    rom[9590] = 25'b0000100010111011101100000;
    rom[9591] = 25'b0000100011000000001001110;
    rom[9592] = 25'b0000100011000100100010110;
    rom[9593] = 25'b0000100011001000110111000;
    rom[9594] = 25'b0000100011001101000110010;
    rom[9595] = 25'b0000100011010001010000110;
    rom[9596] = 25'b0000100011010101010110100;
    rom[9597] = 25'b0000100011011001010111100;
    rom[9598] = 25'b0000100011011101010011101;
    rom[9599] = 25'b0000100011100001001011000;
    rom[9600] = 25'b0000100011100100111101101;
    rom[9601] = 25'b0000100011101000101011100;
    rom[9602] = 25'b0000100011101100010100100;
    rom[9603] = 25'b0000100011101111111000111;
    rom[9604] = 25'b0000100011110011011000011;
    rom[9605] = 25'b0000100011110110110011001;
    rom[9606] = 25'b0000100011111010001001010;
    rom[9607] = 25'b0000100011111101011010100;
    rom[9608] = 25'b0000100100000000100111000;
    rom[9609] = 25'b0000100100000011101110111;
    rom[9610] = 25'b0000100100000110110010000;
    rom[9611] = 25'b0000100100001001110000011;
    rom[9612] = 25'b0000100100001100101010000;
    rom[9613] = 25'b0000100100001111011111000;
    rom[9614] = 25'b0000100100010010001111010;
    rom[9615] = 25'b0000100100010100111010110;
    rom[9616] = 25'b0000100100010111100001110;
    rom[9617] = 25'b0000100100011010000011111;
    rom[9618] = 25'b0000100100011100100001100;
    rom[9619] = 25'b0000100100011110111010011;
    rom[9620] = 25'b0000100100100001001110101;
    rom[9621] = 25'b0000100100100011011110001;
    rom[9622] = 25'b0000100100100101101001000;
    rom[9623] = 25'b0000100100100111101111010;
    rom[9624] = 25'b0000100100101001110001000;
    rom[9625] = 25'b0000100100101011101110000;
    rom[9626] = 25'b0000100100101101100110100;
    rom[9627] = 25'b0000100100101111011010010;
    rom[9628] = 25'b0000100100110001001001100;
    rom[9629] = 25'b0000100100110010110100001;
    rom[9630] = 25'b0000100100110100011010001;
    rom[9631] = 25'b0000100100110101111011101;
    rom[9632] = 25'b0000100100110111011000100;
    rom[9633] = 25'b0000100100111000110001000;
    rom[9634] = 25'b0000100100111010000100110;
    rom[9635] = 25'b0000100100111011010100001;
    rom[9636] = 25'b0000100100111100011110111;
    rom[9637] = 25'b0000100100111101100101001;
    rom[9638] = 25'b0000100100111110100110110;
    rom[9639] = 25'b0000100100111111100100000;
    rom[9640] = 25'b0000100101000000011100110;
    rom[9641] = 25'b0000100101000001010001000;
    rom[9642] = 25'b0000100101000010000000111;
    rom[9643] = 25'b0000100101000010101100001;
    rom[9644] = 25'b0000100101000011010011000;
    rom[9645] = 25'b0000100101000011110101011;
    rom[9646] = 25'b0000100101000100010011100;
    rom[9647] = 25'b0000100101000100101101000;
    rom[9648] = 25'b0000100101000101000010001;
    rom[9649] = 25'b0000100101000101010010111;
    rom[9650] = 25'b0000100101000101011111010;
    rom[9651] = 25'b0000100101000101100111010;
    rom[9652] = 25'b0000100101000101101010111;
    rom[9653] = 25'b0000100101000101101010001;
    rom[9654] = 25'b0000100101000101100101000;
    rom[9655] = 25'b0000100101000101011011100;
    rom[9656] = 25'b0000100101000101001101111;
    rom[9657] = 25'b0000100101000100111011101;
    rom[9658] = 25'b0000100101000100100101011;
    rom[9659] = 25'b0000100101000100001010101;
    rom[9660] = 25'b0000100101000011101011110;
    rom[9661] = 25'b0000100101000011001000011;
    rom[9662] = 25'b0000100101000010100001000;
    rom[9663] = 25'b0000100101000001110101001;
    rom[9664] = 25'b0000100101000001000101010;
    rom[9665] = 25'b0000100101000000010001000;
    rom[9666] = 25'b0000100100111111011000100;
    rom[9667] = 25'b0000100100111110011100000;
    rom[9668] = 25'b0000100100111101011011001;
    rom[9669] = 25'b0000100100111100010110001;
    rom[9670] = 25'b0000100100111011001101000;
    rom[9671] = 25'b0000100100111001111111101;
    rom[9672] = 25'b0000100100111000101110010;
    rom[9673] = 25'b0000100100110111011000101;
    rom[9674] = 25'b0000100100110101111111000;
    rom[9675] = 25'b0000100100110100100001001;
    rom[9676] = 25'b0000100100110010111111010;
    rom[9677] = 25'b0000100100110001011001010;
    rom[9678] = 25'b0000100100101111101111010;
    rom[9679] = 25'b0000100100101110000001001;
    rom[9680] = 25'b0000100100101100001111001;
    rom[9681] = 25'b0000100100101010011001000;
    rom[9682] = 25'b0000100100101000011110111;
    rom[9683] = 25'b0000100100100110100000101;
    rom[9684] = 25'b0000100100100100011110100;
    rom[9685] = 25'b0000100100100010011000100;
    rom[9686] = 25'b0000100100100000001110011;
    rom[9687] = 25'b0000100100011110000000011;
    rom[9688] = 25'b0000100100011011101110011;
    rom[9689] = 25'b0000100100011001011000100;
    rom[9690] = 25'b0000100100010110111110111;
    rom[9691] = 25'b0000100100010100100001001;
    rom[9692] = 25'b0000100100010001111111101;
    rom[9693] = 25'b0000100100001111011010010;
    rom[9694] = 25'b0000100100001100110001000;
    rom[9695] = 25'b0000100100001010000011111;
    rom[9696] = 25'b0000100100000111010011001;
    rom[9697] = 25'b0000100100000100011110011;
    rom[9698] = 25'b0000100100000001100110000;
    rom[9699] = 25'b0000100011111110101001101;
    rom[9700] = 25'b0000100011111011101001101;
    rom[9701] = 25'b0000100011111000100110000;
    rom[9702] = 25'b0000100011110101011110100;
    rom[9703] = 25'b0000100011110010010011011;
    rom[9704] = 25'b0000100011101111000100011;
    rom[9705] = 25'b0000100011101011110001111;
    rom[9706] = 25'b0000100011101000011011100;
    rom[9707] = 25'b0000100011100101000001110;
    rom[9708] = 25'b0000100011100001100100001;
    rom[9709] = 25'b0000100011011110000011000;
    rom[9710] = 25'b0000100011011010011110010;
    rom[9711] = 25'b0000100011010110110101110;
    rom[9712] = 25'b0000100011010011001001111;
    rom[9713] = 25'b0000100011001111011010011;
    rom[9714] = 25'b0000100011001011100111011;
    rom[9715] = 25'b0000100011000111110000110;
    rom[9716] = 25'b0000100011000011110110101;
    rom[9717] = 25'b0000100010111111111001000;
    rom[9718] = 25'b0000100010111011110111111;
    rom[9719] = 25'b0000100010110111110011011;
    rom[9720] = 25'b0000100010110011101011010;
    rom[9721] = 25'b0000100010101111011111111;
    rom[9722] = 25'b0000100010101011010001000;
    rom[9723] = 25'b0000100010100110111110110;
    rom[9724] = 25'b0000100010100010101001000;
    rom[9725] = 25'b0000100010011110010000000;
    rom[9726] = 25'b0000100010011001110011101;
    rom[9727] = 25'b0000100010010101010011111;
    rom[9728] = 25'b0000100010010000110000110;
    rom[9729] = 25'b0000100010001100001010011;
    rom[9730] = 25'b0000100010000111100000110;
    rom[9731] = 25'b0000100010000010110011111;
    rom[9732] = 25'b0000100001111110000011101;
    rom[9733] = 25'b0000100001111001010000010;
    rom[9734] = 25'b0000100001110100011001101;
    rom[9735] = 25'b0000100001101111011111101;
    rom[9736] = 25'b0000100001101010100010101;
    rom[9737] = 25'b0000100001100101100010100;
    rom[9738] = 25'b0000100001100000011111000;
    rom[9739] = 25'b0000100001011011011000101;
    rom[9740] = 25'b0000100001010110001110111;
    rom[9741] = 25'b0000100001010001000010001;
    rom[9742] = 25'b0000100001001011110010010;
    rom[9743] = 25'b0000100001000110011111100;
    rom[9744] = 25'b0000100001000001001001100;
    rom[9745] = 25'b0000100000111011110000100;
    rom[9746] = 25'b0000100000110110010100011;
    rom[9747] = 25'b0000100000110000110101100;
    rom[9748] = 25'b0000100000101011010011100;
    rom[9749] = 25'b0000100000100101101110100;
    rom[9750] = 25'b0000100000100000000110100;
    rom[9751] = 25'b0000100000011010011011101;
    rom[9752] = 25'b0000100000010100101101111;
    rom[9753] = 25'b0000100000001110111101010;
    rom[9754] = 25'b0000100000001001001001101;
    rom[9755] = 25'b0000100000000011010011010;
    rom[9756] = 25'b0000011111111101011010000;
    rom[9757] = 25'b0000011111110111011110000;
    rom[9758] = 25'b0000011111110001011111000;
    rom[9759] = 25'b0000011111101011011101100;
    rom[9760] = 25'b0000011111100101011001000;
    rom[9761] = 25'b0000011111011111010001110;
    rom[9762] = 25'b0000011111011001000111110;
    rom[9763] = 25'b0000011111010010111011001;
    rom[9764] = 25'b0000011111001100101011110;
    rom[9765] = 25'b0000011111000110011001110;
    rom[9766] = 25'b0000011111000000000101000;
    rom[9767] = 25'b0000011110111001101101110;
    rom[9768] = 25'b0000011110110011010011101;
    rom[9769] = 25'b0000011110101100110111001;
    rom[9770] = 25'b0000011110100110010111111;
    rom[9771] = 25'b0000011110011111110110001;
    rom[9772] = 25'b0000011110011001010001111;
    rom[9773] = 25'b0000011110010010101011000;
    rom[9774] = 25'b0000011110001100000001101;
    rom[9775] = 25'b0000011110000101010101110;
    rom[9776] = 25'b0000011101111110100111011;
    rom[9777] = 25'b0000011101110111110110100;
    rom[9778] = 25'b0000011101110001000011010;
    rom[9779] = 25'b0000011101101010001101100;
    rom[9780] = 25'b0000011101100011010101100;
    rom[9781] = 25'b0000011101011100011010111;
    rom[9782] = 25'b0000011101010101011110001;
    rom[9783] = 25'b0000011101001110011110111;
    rom[9784] = 25'b0000011101000111011101011;
    rom[9785] = 25'b0000011101000000011001011;
    rom[9786] = 25'b0000011100111001010011010;
    rom[9787] = 25'b0000011100110010001010111;
    rom[9788] = 25'b0000011100101011000000001;
    rom[9789] = 25'b0000011100100011110011001;
    rom[9790] = 25'b0000011100011100100100000;
    rom[9791] = 25'b0000011100010101010010101;
    rom[9792] = 25'b0000011100001101111111000;
    rom[9793] = 25'b0000011100000110101001010;
    rom[9794] = 25'b0000011011111111010001100;
    rom[9795] = 25'b0000011011110111110111011;
    rom[9796] = 25'b0000011011110000011011010;
    rom[9797] = 25'b0000011011101000111101000;
    rom[9798] = 25'b0000011011100001011100111;
    rom[9799] = 25'b0000011011011001111010100;
    rom[9800] = 25'b0000011011010010010110000;
    rom[9801] = 25'b0000011011001010101111101;
    rom[9802] = 25'b0000011011000011000111010;
    rom[9803] = 25'b0000011010111011011100111;
    rom[9804] = 25'b0000011010110011110000101;
    rom[9805] = 25'b0000011010101100000010011;
    rom[9806] = 25'b0000011010100100010010001;
    rom[9807] = 25'b0000011010011100100000000;
    rom[9808] = 25'b0000011010010100101100000;
    rom[9809] = 25'b0000011010001100110110010;
    rom[9810] = 25'b0000011010000100111110100;
    rom[9811] = 25'b0000011001111101000101000;
    rom[9812] = 25'b0000011001110101001001110;
    rom[9813] = 25'b0000011001101101001100100;
    rom[9814] = 25'b0000011001100101001101110;
    rom[9815] = 25'b0000011001011101001101001;
    rom[9816] = 25'b0000011001010101001010101;
    rom[9817] = 25'b0000011001001101000110101;
    rom[9818] = 25'b0000011001000101000000111;
    rom[9819] = 25'b0000011000111100111001011;
    rom[9820] = 25'b0000011000110100110000010;
    rom[9821] = 25'b0000011000101100100101100;
    rom[9822] = 25'b0000011000100100011001001;
    rom[9823] = 25'b0000011000011100001011001;
    rom[9824] = 25'b0000011000010011111011101;
    rom[9825] = 25'b0000011000001011101010100;
    rom[9826] = 25'b0000011000000011010111111;
    rom[9827] = 25'b0000010111111011000011110;
    rom[9828] = 25'b0000010111110010101110000;
    rom[9829] = 25'b0000010111101010010110111;
    rom[9830] = 25'b0000010111100001111110010;
    rom[9831] = 25'b0000010111011001100100001;
    rom[9832] = 25'b0000010111010001001000101;
    rom[9833] = 25'b0000010111001000101011110;
    rom[9834] = 25'b0000010111000000001101011;
    rom[9835] = 25'b0000010110110111101101110;
    rom[9836] = 25'b0000010110101111001100110;
    rom[9837] = 25'b0000010110100110101010011;
    rom[9838] = 25'b0000010110011110000110110;
    rom[9839] = 25'b0000010110010101100001110;
    rom[9840] = 25'b0000010110001100111011100;
    rom[9841] = 25'b0000010110000100010100000;
    rom[9842] = 25'b0000010101111011101011001;
    rom[9843] = 25'b0000010101110011000001010;
    rom[9844] = 25'b0000010101101010010110001;
    rom[9845] = 25'b0000010101100001101001110;
    rom[9846] = 25'b0000010101011000111100010;
    rom[9847] = 25'b0000010101010000001101100;
    rom[9848] = 25'b0000010101000111011101110;
    rom[9849] = 25'b0000010100111110101100111;
    rom[9850] = 25'b0000010100110101111010111;
    rom[9851] = 25'b0000010100101101000111111;
    rom[9852] = 25'b0000010100100100010011110;
    rom[9853] = 25'b0000010100011011011110101;
    rom[9854] = 25'b0000010100010010101000100;
    rom[9855] = 25'b0000010100001001110001011;
    rom[9856] = 25'b0000010100000000111001010;
    rom[9857] = 25'b0000010011111000000000001;
    rom[9858] = 25'b0000010011101111000110001;
    rom[9859] = 25'b0000010011100110001011001;
    rom[9860] = 25'b0000010011011101001111011;
    rom[9861] = 25'b0000010011010100010010110;
    rom[9862] = 25'b0000010011001011010101001;
    rom[9863] = 25'b0000010011000010010110101;
    rom[9864] = 25'b0000010010111001010111011;
    rom[9865] = 25'b0000010010110000010111011;
    rom[9866] = 25'b0000010010100111010110100;
    rom[9867] = 25'b0000010010011110010101000;
    rom[9868] = 25'b0000010010010101010010100;
    rom[9869] = 25'b0000010010001100001111100;
    rom[9870] = 25'b0000010010000011001011101;
    rom[9871] = 25'b0000010001111010000111001;
    rom[9872] = 25'b0000010001110001000001111;
    rom[9873] = 25'b0000010001100111111100001;
    rom[9874] = 25'b0000010001011110110101101;
    rom[9875] = 25'b0000010001010101101110100;
    rom[9876] = 25'b0000010001001100100110110;
    rom[9877] = 25'b0000010001000011011110011;
    rom[9878] = 25'b0000010000111010010101100;
    rom[9879] = 25'b0000010000110001001100001;
    rom[9880] = 25'b0000010000101000000010001;
    rom[9881] = 25'b0000010000011110110111101;
    rom[9882] = 25'b0000010000010101101100101;
    rom[9883] = 25'b0000010000001100100001010;
    rom[9884] = 25'b0000010000000011010101011;
    rom[9885] = 25'b0000001111111010001001000;
    rom[9886] = 25'b0000001111110000111100010;
    rom[9887] = 25'b0000001111100111101111000;
    rom[9888] = 25'b0000001111011110100001011;
    rom[9889] = 25'b0000001111010101010011100;
    rom[9890] = 25'b0000001111001100000101010;
    rom[9891] = 25'b0000001111000010110110101;
    rom[9892] = 25'b0000001110111001100111101;
    rom[9893] = 25'b0000001110110000011000011;
    rom[9894] = 25'b0000001110100111001000111;
    rom[9895] = 25'b0000001110011101111001001;
    rom[9896] = 25'b0000001110010100101001001;
    rom[9897] = 25'b0000001110001011011000110;
    rom[9898] = 25'b0000001110000010001000011;
    rom[9899] = 25'b0000001101111000110111101;
    rom[9900] = 25'b0000001101101111100110111;
    rom[9901] = 25'b0000001101100110010101111;
    rom[9902] = 25'b0000001101011101000100110;
    rom[9903] = 25'b0000001101010011110011100;
    rom[9904] = 25'b0000001101001010100010000;
    rom[9905] = 25'b0000001101000001010000101;
    rom[9906] = 25'b0000001100110111111111001;
    rom[9907] = 25'b0000001100101110101101100;
    rom[9908] = 25'b0000001100100101011011111;
    rom[9909] = 25'b0000001100011100001010010;
    rom[9910] = 25'b0000001100010010111000110;
    rom[9911] = 25'b0000001100001001100111000;
    rom[9912] = 25'b0000001100000000010101011;
    rom[9913] = 25'b0000001011110111000011111;
    rom[9914] = 25'b0000001011101101110010011;
    rom[9915] = 25'b0000001011100100100001000;
    rom[9916] = 25'b0000001011011011001111110;
    rom[9917] = 25'b0000001011010001111110100;
    rom[9918] = 25'b0000001011001000101101100;
    rom[9919] = 25'b0000001010111111011100101;
    rom[9920] = 25'b0000001010110110001100000;
    rom[9921] = 25'b0000001010101100111011011;
    rom[9922] = 25'b0000001010100011101011001;
    rom[9923] = 25'b0000001010011010011010111;
    rom[9924] = 25'b0000001010010001001011001;
    rom[9925] = 25'b0000001010000111111011100;
    rom[9926] = 25'b0000001001111110101100000;
    rom[9927] = 25'b0000001001110101011101000;
    rom[9928] = 25'b0000001001101100001110001;
    rom[9929] = 25'b0000001001100010111111110;
    rom[9930] = 25'b0000001001011001110001101;
    rom[9931] = 25'b0000001001010000100011110;
    rom[9932] = 25'b0000001001000111010110011;
    rom[9933] = 25'b0000001000111110001001010;
    rom[9934] = 25'b0000001000110100111100101;
    rom[9935] = 25'b0000001000101011110000011;
    rom[9936] = 25'b0000001000100010100100101;
    rom[9937] = 25'b0000001000011001011001010;
    rom[9938] = 25'b0000001000010000001110010;
    rom[9939] = 25'b0000001000000111000011111;
    rom[9940] = 25'b0000000111111101111001111;
    rom[9941] = 25'b0000000111110100110000100;
    rom[9942] = 25'b0000000111101011100111101;
    rom[9943] = 25'b0000000111100010011111001;
    rom[9944] = 25'b0000000111011001010111011;
    rom[9945] = 25'b0000000111010000010000001;
    rom[9946] = 25'b0000000111000111001001100;
    rom[9947] = 25'b0000000110111110000011100;
    rom[9948] = 25'b0000000110110100111101111;
    rom[9949] = 25'b0000000110101011111001001;
    rom[9950] = 25'b0000000110100010110101000;
    rom[9951] = 25'b0000000110011001110001100;
    rom[9952] = 25'b0000000110010000101110101;
    rom[9953] = 25'b0000000110000111101100100;
    rom[9954] = 25'b0000000101111110101011000;
    rom[9955] = 25'b0000000101110101101010011;
    rom[9956] = 25'b0000000101101100101010011;
    rom[9957] = 25'b0000000101100011101011001;
    rom[9958] = 25'b0000000101011010101100101;
    rom[9959] = 25'b0000000101010001101110111;
    rom[9960] = 25'b0000000101001000110010000;
    rom[9961] = 25'b0000000100111111110110000;
    rom[9962] = 25'b0000000100110110111010110;
    rom[9963] = 25'b0000000100101110000000010;
    rom[9964] = 25'b0000000100100101000110110;
    rom[9965] = 25'b0000000100011100001110001;
    rom[9966] = 25'b0000000100010011010110010;
    rom[9967] = 25'b0000000100001010011111010;
    rom[9968] = 25'b0000000100000001101001010;
    rom[9969] = 25'b0000000011111000110100010;
    rom[9970] = 25'b0000000011110000000000000;
    rom[9971] = 25'b0000000011100111001100111;
    rom[9972] = 25'b0000000011011110011010101;
    rom[9973] = 25'b0000000011010101101001011;
    rom[9974] = 25'b0000000011001100111001001;
    rom[9975] = 25'b0000000011000100001001111;
    rom[9976] = 25'b0000000010111011011011101;
    rom[9977] = 25'b0000000010110010101110100;
    rom[9978] = 25'b0000000010101010000010010;
    rom[9979] = 25'b0000000010100001010111010;
    rom[9980] = 25'b0000000010011000101101010;
    rom[9981] = 25'b0000000010010000000100010;
    rom[9982] = 25'b0000000010000111011100100;
    rom[9983] = 25'b0000000001111110110101111;
    rom[9984] = 25'b0000000001110110010000010;
    rom[9985] = 25'b0000000001101101101011110;
    rom[9986] = 25'b0000000001100101001000100;
    rom[9987] = 25'b0000000001011100100110011;
    rom[9988] = 25'b0000000001010100000101100;
    rom[9989] = 25'b0000000001001011100101110;
    rom[9990] = 25'b0000000001000011000111001;
    rom[9991] = 25'b0000000000111010101001111;
    rom[9992] = 25'b0000000000110010001101110;
    rom[9993] = 25'b0000000000101001110011000;
    rom[9994] = 25'b0000000000100001011001011;
    rom[9995] = 25'b0000000000011001000001001;
    rom[9996] = 25'b0000000000010000101010000;
    rom[9997] = 25'b0000000000001000010100011;
    rom[9998] = 25'b0000000000000000000000000;
    rom[9999] = 25'b1111111111110111101100111;
    rom[10000] = 25'b1111111111101111011011000;
    rom[10001] = 25'b1111111111100111001010101;
    rom[10002] = 25'b1111111111011110111011101;
    rom[10003] = 25'b1111111111010110101101111;
    rom[10004] = 25'b1111111111001110100001100;
    rom[10005] = 25'b1111111111000110010110101;
    rom[10006] = 25'b1111111110111110001101000;
    rom[10007] = 25'b1111111110110110000100111;
    rom[10008] = 25'b1111111110101101111110001;
    rom[10009] = 25'b1111111110100101111000111;
    rom[10010] = 25'b1111111110011101110101001;
    rom[10011] = 25'b1111111110010101110010101;
    rom[10012] = 25'b1111111110001101110001110;
    rom[10013] = 25'b1111111110000101110010011;
    rom[10014] = 25'b1111111101111101110100100;
    rom[10015] = 25'b1111111101110101111000000;
    rom[10016] = 25'b1111111101101101111101001;
    rom[10017] = 25'b1111111101100110000011110;
    rom[10018] = 25'b1111111101011110001011111;
    rom[10019] = 25'b1111111101010110010101101;
    rom[10020] = 25'b1111111101001110100000110;
    rom[10021] = 25'b1111111101000110101101101;
    rom[10022] = 25'b1111111100111110111100001;
    rom[10023] = 25'b1111111100110111001100000;
    rom[10024] = 25'b1111111100101111011101110;
    rom[10025] = 25'b1111111100100111110000111;
    rom[10026] = 25'b1111111100100000000101101;
    rom[10027] = 25'b1111111100011000011100001;
    rom[10028] = 25'b1111111100010000110100010;
    rom[10029] = 25'b1111111100001001001110000;
    rom[10030] = 25'b1111111100000001101001011;
    rom[10031] = 25'b1111111011111010000110100;
    rom[10032] = 25'b1111111011110010100101010;
    rom[10033] = 25'b1111111011101011000101110;
    rom[10034] = 25'b1111111011100011100111111;
    rom[10035] = 25'b1111111011011100001011110;
    rom[10036] = 25'b1111111011010100110001011;
    rom[10037] = 25'b1111111011001101011000110;
    rom[10038] = 25'b1111111011000110000001110;
    rom[10039] = 25'b1111111010111110101100100;
    rom[10040] = 25'b1111111010110111011001000;
    rom[10041] = 25'b1111111010110000000111011;
    rom[10042] = 25'b1111111010101000110111100;
    rom[10043] = 25'b1111111010100001101001011;
    rom[10044] = 25'b1111111010011010011101001;
    rom[10045] = 25'b1111111010010011010010100;
    rom[10046] = 25'b1111111010001100001001111;
    rom[10047] = 25'b1111111010000101000011000;
    rom[10048] = 25'b1111111001111101111101111;
    rom[10049] = 25'b1111111001110110111010110;
    rom[10050] = 25'b1111111001101111111001011;
    rom[10051] = 25'b1111111001101000111001110;
    rom[10052] = 25'b1111111001100001111100001;
    rom[10053] = 25'b1111111001011011000000011;
    rom[10054] = 25'b1111111001010100000110011;
    rom[10055] = 25'b1111111001001101001110100;
    rom[10056] = 25'b1111111001000110011000010;
    rom[10057] = 25'b1111111000111111100100001;
    rom[10058] = 25'b1111111000111000110001110;
    rom[10059] = 25'b1111111000110010000001011;
    rom[10060] = 25'b1111111000101011010011000;
    rom[10061] = 25'b1111111000100100100110011;
    rom[10062] = 25'b1111111000011101111011111;
    rom[10063] = 25'b1111111000010111010011010;
    rom[10064] = 25'b1111111000010000101100101;
    rom[10065] = 25'b1111111000001010000111111;
    rom[10066] = 25'b1111111000000011100101001;
    rom[10067] = 25'b1111110111111101000100011;
    rom[10068] = 25'b1111110111110110100101101;
    rom[10069] = 25'b1111110111110000001000111;
    rom[10070] = 25'b1111110111101001101110001;
    rom[10071] = 25'b1111110111100011010101011;
    rom[10072] = 25'b1111110111011100111110101;
    rom[10073] = 25'b1111110111010110101001111;
    rom[10074] = 25'b1111110111010000010111001;
    rom[10075] = 25'b1111110111001010000110011;
    rom[10076] = 25'b1111110111000011110111111;
    rom[10077] = 25'b1111110110111101101011011;
    rom[10078] = 25'b1111110110110111100000110;
    rom[10079] = 25'b1111110110110001011000010;
    rom[10080] = 25'b1111110110101011010001111;
    rom[10081] = 25'b1111110110100101001101100;
    rom[10082] = 25'b1111110110011111001011011;
    rom[10083] = 25'b1111110110011001001011010;
    rom[10084] = 25'b1111110110010011001101001;
    rom[10085] = 25'b1111110110001101010001001;
    rom[10086] = 25'b1111110110000111010111011;
    rom[10087] = 25'b1111110110000001011111101;
    rom[10088] = 25'b1111110101111011101010000;
    rom[10089] = 25'b1111110101110101110110100;
    rom[10090] = 25'b1111110101110000000101000;
    rom[10091] = 25'b1111110101101010010101111;
    rom[10092] = 25'b1111110101100100101000101;
    rom[10093] = 25'b1111110101011110111101110;
    rom[10094] = 25'b1111110101011001010100111;
    rom[10095] = 25'b1111110101010011101110010;
    rom[10096] = 25'b1111110101001110001001110;
    rom[10097] = 25'b1111110101001000100111011;
    rom[10098] = 25'b1111110101000011000111001;
    rom[10099] = 25'b1111110100111101101001010;
    rom[10100] = 25'b1111110100111000001101011;
    rom[10101] = 25'b1111110100110010110011110;
    rom[10102] = 25'b1111110100101101011100010;
    rom[10103] = 25'b1111110100101000000111000;
    rom[10104] = 25'b1111110100100010110011111;
    rom[10105] = 25'b1111110100011101100011000;
    rom[10106] = 25'b1111110100011000010100011;
    rom[10107] = 25'b1111110100010011000111111;
    rom[10108] = 25'b1111110100001101111101101;
    rom[10109] = 25'b1111110100001000110101100;
    rom[10110] = 25'b1111110100000011101111110;
    rom[10111] = 25'b1111110011111110101100001;
    rom[10112] = 25'b1111110011111001101010110;
    rom[10113] = 25'b1111110011110100101011101;
    rom[10114] = 25'b1111110011101111101110111;
    rom[10115] = 25'b1111110011101010110100001;
    rom[10116] = 25'b1111110011100101111011110;
    rom[10117] = 25'b1111110011100001000101101;
    rom[10118] = 25'b1111110011011100010001110;
    rom[10119] = 25'b1111110011010111100000000;
    rom[10120] = 25'b1111110011010010110000101;
    rom[10121] = 25'b1111110011001110000011100;
    rom[10122] = 25'b1111110011001001011000101;
    rom[10123] = 25'b1111110011000100110000000;
    rom[10124] = 25'b1111110011000000001001101;
    rom[10125] = 25'b1111110010111011100101101;
    rom[10126] = 25'b1111110010110111000011110;
    rom[10127] = 25'b1111110010110010100100010;
    rom[10128] = 25'b1111110010101110000111001;
    rom[10129] = 25'b1111110010101001101100001;
    rom[10130] = 25'b1111110010100101010011100;
    rom[10131] = 25'b1111110010100000111101001;
    rom[10132] = 25'b1111110010011100101001000;
    rom[10133] = 25'b1111110010011000010111010;
    rom[10134] = 25'b1111110010010100000111110;
    rom[10135] = 25'b1111110010001111111010100;
    rom[10136] = 25'b1111110010001011101111110;
    rom[10137] = 25'b1111110010000111100111001;
    rom[10138] = 25'b1111110010000011100000110;
    rom[10139] = 25'b1111110001111111011100111;
    rom[10140] = 25'b1111110001111011011011001;
    rom[10141] = 25'b1111110001110111011011110;
    rom[10142] = 25'b1111110001110011011110110;
    rom[10143] = 25'b1111110001101111100100000;
    rom[10144] = 25'b1111110001101011101011100;
    rom[10145] = 25'b1111110001100111110101011;
    rom[10146] = 25'b1111110001100100000001101;
    rom[10147] = 25'b1111110001100000010000010;
    rom[10148] = 25'b1111110001011100100001000;
    rom[10149] = 25'b1111110001011000110100010;
    rom[10150] = 25'b1111110001010101001001110;
    rom[10151] = 25'b1111110001010001100001100;
    rom[10152] = 25'b1111110001001101111011110;
    rom[10153] = 25'b1111110001001010011000010;
    rom[10154] = 25'b1111110001000110110110111;
    rom[10155] = 25'b1111110001000011011000001;
    rom[10156] = 25'b1111110000111111111011100;
    rom[10157] = 25'b1111110000111100100001010;
    rom[10158] = 25'b1111110000111001001001011;
    rom[10159] = 25'b1111110000110101110011111;
    rom[10160] = 25'b1111110000110010100000101;
    rom[10161] = 25'b1111110000101111001111110;
    rom[10162] = 25'b1111110000101100000001000;
    rom[10163] = 25'b1111110000101000110100110;
    rom[10164] = 25'b1111110000100101101010111;
    rom[10165] = 25'b1111110000100010100011011;
    rom[10166] = 25'b1111110000011111011110000;
    rom[10167] = 25'b1111110000011100011011001;
    rom[10168] = 25'b1111110000011001011010100;
    rom[10169] = 25'b1111110000010110011100010;
    rom[10170] = 25'b1111110000010011100000010;
    rom[10171] = 25'b1111110000010000100110110;
    rom[10172] = 25'b1111110000001101101111100;
    rom[10173] = 25'b1111110000001010111010100;
    rom[10174] = 25'b1111110000001000000111111;
    rom[10175] = 25'b1111110000000101010111100;
    rom[10176] = 25'b1111110000000010101001101;
    rom[10177] = 25'b1111101111111111111101111;
    rom[10178] = 25'b1111101111111101010100101;
    rom[10179] = 25'b1111101111111010101101101;
    rom[10180] = 25'b1111101111111000001001000;
    rom[10181] = 25'b1111101111110101100110101;
    rom[10182] = 25'b1111101111110011000110101;
    rom[10183] = 25'b1111101111110000101000111;
    rom[10184] = 25'b1111101111101110001101101;
    rom[10185] = 25'b1111101111101011110100100;
    rom[10186] = 25'b1111101111101001011101110;
    rom[10187] = 25'b1111101111100111001001010;
    rom[10188] = 25'b1111101111100100110111001;
    rom[10189] = 25'b1111101111100010100111011;
    rom[10190] = 25'b1111101111100000011001111;
    rom[10191] = 25'b1111101111011110001110101;
    rom[10192] = 25'b1111101111011100000101110;
    rom[10193] = 25'b1111101111011001111111010;
    rom[10194] = 25'b1111101111010111111011000;
    rom[10195] = 25'b1111101111010101111001000;
    rom[10196] = 25'b1111101111010011111001010;
    rom[10197] = 25'b1111101111010001111011111;
    rom[10198] = 25'b1111101111010000000000110;
    rom[10199] = 25'b1111101111001110001000000;
    rom[10200] = 25'b1111101111001100010001101;
    rom[10201] = 25'b1111101111001010011101011;
    rom[10202] = 25'b1111101111001000101011100;
    rom[10203] = 25'b1111101111000110111011110;
    rom[10204] = 25'b1111101111000101001110100;
    rom[10205] = 25'b1111101111000011100011011;
    rom[10206] = 25'b1111101111000001111010101;
    rom[10207] = 25'b1111101111000000010100000;
    rom[10208] = 25'b1111101110111110101111110;
    rom[10209] = 25'b1111101110111101001101111;
    rom[10210] = 25'b1111101110111011101110001;
    rom[10211] = 25'b1111101110111010010000101;
    rom[10212] = 25'b1111101110111000110101100;
    rom[10213] = 25'b1111101110110111011100100;
    rom[10214] = 25'b1111101110110110000101111;
    rom[10215] = 25'b1111101110110100110001100;
    rom[10216] = 25'b1111101110110011011111011;
    rom[10217] = 25'b1111101110110010001111011;
    rom[10218] = 25'b1111101110110001000001101;
    rom[10219] = 25'b1111101110101111110110001;
    rom[10220] = 25'b1111101110101110101101000;
    rom[10221] = 25'b1111101110101101100110000;
    rom[10222] = 25'b1111101110101100100001010;
    rom[10223] = 25'b1111101110101011011110101;
    rom[10224] = 25'b1111101110101010011110011;
    rom[10225] = 25'b1111101110101001100000010;
    rom[10226] = 25'b1111101110101000100100011;
    rom[10227] = 25'b1111101110100111101010110;
    rom[10228] = 25'b1111101110100110110011010;
    rom[10229] = 25'b1111101110100101111110000;
    rom[10230] = 25'b1111101110100101001010111;
    rom[10231] = 25'b1111101110100100011010000;
    rom[10232] = 25'b1111101110100011101011011;
    rom[10233] = 25'b1111101110100010111110110;
    rom[10234] = 25'b1111101110100010010100100;
    rom[10235] = 25'b1111101110100001101100010;
    rom[10236] = 25'b1111101110100001000110011;
    rom[10237] = 25'b1111101110100000100010100;
    rom[10238] = 25'b1111101110100000000000111;
    rom[10239] = 25'b1111101110011111100001100;
    rom[10240] = 25'b1111101110011111000100001;
    rom[10241] = 25'b1111101110011110101000111;
    rom[10242] = 25'b1111101110011110001111111;
    rom[10243] = 25'b1111101110011101111001000;
    rom[10244] = 25'b1111101110011101100100010;
    rom[10245] = 25'b1111101110011101010001101;
    rom[10246] = 25'b1111101110011101000001001;
    rom[10247] = 25'b1111101110011100110010101;
    rom[10248] = 25'b1111101110011100100110100;
    rom[10249] = 25'b1111101110011100011100011;
    rom[10250] = 25'b1111101110011100010100010;
    rom[10251] = 25'b1111101110011100001110010;
    rom[10252] = 25'b1111101110011100001010100;
    rom[10253] = 25'b1111101110011100001000110;
    rom[10254] = 25'b1111101110011100001001001;
    rom[10255] = 25'b1111101110011100001011100;
    rom[10256] = 25'b1111101110011100010000000;
    rom[10257] = 25'b1111101110011100010110100;
    rom[10258] = 25'b1111101110011100011111010;
    rom[10259] = 25'b1111101110011100101001111;
    rom[10260] = 25'b1111101110011100110110101;
    rom[10261] = 25'b1111101110011101000101011;
    rom[10262] = 25'b1111101110011101010110010;
    rom[10263] = 25'b1111101110011101101001001;
    rom[10264] = 25'b1111101110011101111110000;
    rom[10265] = 25'b1111101110011110010101000;
    rom[10266] = 25'b1111101110011110101101111;
    rom[10267] = 25'b1111101110011111001000111;
    rom[10268] = 25'b1111101110011111100101110;
    rom[10269] = 25'b1111101110100000000100111;
    rom[10270] = 25'b1111101110100000100101110;
    rom[10271] = 25'b1111101110100001001000110;
    rom[10272] = 25'b1111101110100001101101101;
    rom[10273] = 25'b1111101110100010010100110;
    rom[10274] = 25'b1111101110100010111101100;
    rom[10275] = 25'b1111101110100011101000100;
    rom[10276] = 25'b1111101110100100010101010;
    rom[10277] = 25'b1111101110100101000100000;
    rom[10278] = 25'b1111101110100101110100110;
    rom[10279] = 25'b1111101110100110100111011;
    rom[10280] = 25'b1111101110100111011100000;
    rom[10281] = 25'b1111101110101000010010100;
    rom[10282] = 25'b1111101110101001001011000;
    rom[10283] = 25'b1111101110101010000101011;
    rom[10284] = 25'b1111101110101011000001110;
    rom[10285] = 25'b1111101110101011111111111;
    rom[10286] = 25'b1111101110101101000000000;
    rom[10287] = 25'b1111101110101110000010000;
    rom[10288] = 25'b1111101110101111000101110;
    rom[10289] = 25'b1111101110110000001011100;
    rom[10290] = 25'b1111101110110001010011001;
    rom[10291] = 25'b1111101110110010011100100;
    rom[10292] = 25'b1111101110110011100111111;
    rom[10293] = 25'b1111101110110100110101001;
    rom[10294] = 25'b1111101110110110000100001;
    rom[10295] = 25'b1111101110110111010100111;
    rom[10296] = 25'b1111101110111000100111101;
    rom[10297] = 25'b1111101110111001111100001;
    rom[10298] = 25'b1111101110111011010010100;
    rom[10299] = 25'b1111101110111100101010100;
    rom[10300] = 25'b1111101110111110000100011;
    rom[10301] = 25'b1111101110111111100000001;
    rom[10302] = 25'b1111101111000000111101101;
    rom[10303] = 25'b1111101111000010011100111;
    rom[10304] = 25'b1111101111000011111101111;
    rom[10305] = 25'b1111101111000101100000110;
    rom[10306] = 25'b1111101111000111000101010;
    rom[10307] = 25'b1111101111001000101011101;
    rom[10308] = 25'b1111101111001010010011101;
    rom[10309] = 25'b1111101111001011111101011;
    rom[10310] = 25'b1111101111001101101001000;
    rom[10311] = 25'b1111101111001111010110001;
    rom[10312] = 25'b1111101111010001000101000;
    rom[10313] = 25'b1111101111010010110101110;
    rom[10314] = 25'b1111101111010100101000000;
    rom[10315] = 25'b1111101111010110011100001;
    rom[10316] = 25'b1111101111011000010001111;
    rom[10317] = 25'b1111101111011010001001010;
    rom[10318] = 25'b1111101111011100000010010;
    rom[10319] = 25'b1111101111011101111101000;
    rom[10320] = 25'b1111101111011111111001010;
    rom[10321] = 25'b1111101111100001110111010;
    rom[10322] = 25'b1111101111100011110110111;
    rom[10323] = 25'b1111101111100101111000010;
    rom[10324] = 25'b1111101111100111111011001;
    rom[10325] = 25'b1111101111101001111111100;
    rom[10326] = 25'b1111101111101100000101101;
    rom[10327] = 25'b1111101111101110001101010;
    rom[10328] = 25'b1111101111110000010110101;
    rom[10329] = 25'b1111101111110010100001100;
    rom[10330] = 25'b1111101111110100101101110;
    rom[10331] = 25'b1111101111110110111011110;
    rom[10332] = 25'b1111101111111001001011011;
    rom[10333] = 25'b1111101111111011011100100;
    rom[10334] = 25'b1111101111111101101111000;
    rom[10335] = 25'b1111110000000000000011001;
    rom[10336] = 25'b1111110000000010011000111;
    rom[10337] = 25'b1111110000000100110000000;
    rom[10338] = 25'b1111110000000111001000101;
    rom[10339] = 25'b1111110000001001100010111;
    rom[10340] = 25'b1111110000001011111110101;
    rom[10341] = 25'b1111110000001110011011110;
    rom[10342] = 25'b1111110000010000111010011;
    rom[10343] = 25'b1111110000010011011010011;
    rom[10344] = 25'b1111110000010101111011111;
    rom[10345] = 25'b1111110000011000011110111;
    rom[10346] = 25'b1111110000011011000011011;
    rom[10347] = 25'b1111110000011101101001010;
    rom[10348] = 25'b1111110000100000010000011;
    rom[10349] = 25'b1111110000100010111001001;
    rom[10350] = 25'b1111110000100101100011010;
    rom[10351] = 25'b1111110000101000001110110;
    rom[10352] = 25'b1111110000101010111011101;
    rom[10353] = 25'b1111110000101101101001111;
    rom[10354] = 25'b1111110000110000011001100;
    rom[10355] = 25'b1111110000110011001010100;
    rom[10356] = 25'b1111110000110101111100110;
    rom[10357] = 25'b1111110000111000110000011;
    rom[10358] = 25'b1111110000111011100101100;
    rom[10359] = 25'b1111110000111110011011110;
    rom[10360] = 25'b1111110001000001010011100;
    rom[10361] = 25'b1111110001000100001100100;
    rom[10362] = 25'b1111110001000111000110110;
    rom[10363] = 25'b1111110001001010000010010;
    rom[10364] = 25'b1111110001001100111111001;
    rom[10365] = 25'b1111110001001111111101010;
    rom[10366] = 25'b1111110001010010111100101;
    rom[10367] = 25'b1111110001010101111101010;
    rom[10368] = 25'b1111110001011000111111001;
    rom[10369] = 25'b1111110001011100000010010;
    rom[10370] = 25'b1111110001011111000110101;
    rom[10371] = 25'b1111110001100010001100001;
    rom[10372] = 25'b1111110001100101010011000;
    rom[10373] = 25'b1111110001101000011011000;
    rom[10374] = 25'b1111110001101011100100001;
    rom[10375] = 25'b1111110001101110101110100;
    rom[10376] = 25'b1111110001110001111010001;
    rom[10377] = 25'b1111110001110101000110110;
    rom[10378] = 25'b1111110001111000010100101;
    rom[10379] = 25'b1111110001111011100011101;
    rom[10380] = 25'b1111110001111110110011111;
    rom[10381] = 25'b1111110010000010000101000;
    rom[10382] = 25'b1111110010000101010111100;
    rom[10383] = 25'b1111110010001000101011000;
    rom[10384] = 25'b1111110010001011111111101;
    rom[10385] = 25'b1111110010001111010101011;
    rom[10386] = 25'b1111110010010010101100001;
    rom[10387] = 25'b1111110010010110000100001;
    rom[10388] = 25'b1111110010011001011101001;
    rom[10389] = 25'b1111110010011100110111000;
    rom[10390] = 25'b1111110010100000010010001;
    rom[10391] = 25'b1111110010100011101110010;
    rom[10392] = 25'b1111110010100111001011011;
    rom[10393] = 25'b1111110010101010101001100;
    rom[10394] = 25'b1111110010101110001000101;
    rom[10395] = 25'b1111110010110001101000111;
    rom[10396] = 25'b1111110010110101001010000;
    rom[10397] = 25'b1111110010111000101100001;
    rom[10398] = 25'b1111110010111100001111011;
    rom[10399] = 25'b1111110010111111110011011;
    rom[10400] = 25'b1111110011000011011000100;
    rom[10401] = 25'b1111110011000110111110100;
    rom[10402] = 25'b1111110011001010100101100;
    rom[10403] = 25'b1111110011001110001101011;
    rom[10404] = 25'b1111110011010001110110001;
    rom[10405] = 25'b1111110011010101011111111;
    rom[10406] = 25'b1111110011011001001010100;
    rom[10407] = 25'b1111110011011100110110000;
    rom[10408] = 25'b1111110011100000100010011;
    rom[10409] = 25'b1111110011100100001111101;
    rom[10410] = 25'b1111110011100111111101111;
    rom[10411] = 25'b1111110011101011101100111;
    rom[10412] = 25'b1111110011101111011100101;
    rom[10413] = 25'b1111110011110011001101011;
    rom[10414] = 25'b1111110011110110111110110;
    rom[10415] = 25'b1111110011111010110001001;
    rom[10416] = 25'b1111110011111110100100010;
    rom[10417] = 25'b1111110100000010011000010;
    rom[10418] = 25'b1111110100000110001100111;
    rom[10419] = 25'b1111110100001010000010100;
    rom[10420] = 25'b1111110100001101111000111;
    rom[10421] = 25'b1111110100010001101111111;
    rom[10422] = 25'b1111110100010101100111110;
    rom[10423] = 25'b1111110100011001100000010;
    rom[10424] = 25'b1111110100011101011001101;
    rom[10425] = 25'b1111110100100001010011100;
    rom[10426] = 25'b1111110100100101001110010;
    rom[10427] = 25'b1111110100101001001001110;
    rom[10428] = 25'b1111110100101101000101111;
    rom[10429] = 25'b1111110100110001000010111;
    rom[10430] = 25'b1111110100110101000000010;
    rom[10431] = 25'b1111110100111000111110101;
    rom[10432] = 25'b1111110100111100111101011;
    rom[10433] = 25'b1111110101000000111100111;
    rom[10434] = 25'b1111110101000100111101001;
    rom[10435] = 25'b1111110101001000111101111;
    rom[10436] = 25'b1111110101001100111111010;
    rom[10437] = 25'b1111110101010001000001011;
    rom[10438] = 25'b1111110101010101000100001;
    rom[10439] = 25'b1111110101011001000111010;
    rom[10440] = 25'b1111110101011101001011001;
    rom[10441] = 25'b1111110101100001001111101;
    rom[10442] = 25'b1111110101100101010100101;
    rom[10443] = 25'b1111110101101001011010010;
    rom[10444] = 25'b1111110101101101100000010;
    rom[10445] = 25'b1111110101110001100111000;
    rom[10446] = 25'b1111110101110101101110010;
    rom[10447] = 25'b1111110101111001110101111;
    rom[10448] = 25'b1111110101111101111110001;
    rom[10449] = 25'b1111110110000010000110111;
    rom[10450] = 25'b1111110110000110010000001;
    rom[10451] = 25'b1111110110001010011001111;
    rom[10452] = 25'b1111110110001110100100001;
    rom[10453] = 25'b1111110110010010101110111;
    rom[10454] = 25'b1111110110010110111010000;
    rom[10455] = 25'b1111110110011011000101101;
    rom[10456] = 25'b1111110110011111010001110;
    rom[10457] = 25'b1111110110100011011110001;
    rom[10458] = 25'b1111110110100111101011001;
    rom[10459] = 25'b1111110110101011111000011;
    rom[10460] = 25'b1111110110110000000110001;
    rom[10461] = 25'b1111110110110100010100011;
    rom[10462] = 25'b1111110110111000100010111;
    rom[10463] = 25'b1111110110111100110001110;
    rom[10464] = 25'b1111110111000001000001001;
    rom[10465] = 25'b1111110111000101010000110;
    rom[10466] = 25'b1111110111001001100000110;
    rom[10467] = 25'b1111110111001101110001001;
    rom[10468] = 25'b1111110111010010000001111;
    rom[10469] = 25'b1111110111010110010010111;
    rom[10470] = 25'b1111110111011010100100010;
    rom[10471] = 25'b1111110111011110110101111;
    rom[10472] = 25'b1111110111100011000111111;
    rom[10473] = 25'b1111110111100111011010001;
    rom[10474] = 25'b1111110111101011101100101;
    rom[10475] = 25'b1111110111101111111111011;
    rom[10476] = 25'b1111110111110100010010100;
    rom[10477] = 25'b1111110111111000100101110;
    rom[10478] = 25'b1111110111111100111001100;
    rom[10479] = 25'b1111111000000001001101010;
    rom[10480] = 25'b1111111000000101100001011;
    rom[10481] = 25'b1111111000001001110101101;
    rom[10482] = 25'b1111111000001110001010000;
    rom[10483] = 25'b1111111000010010011110110;
    rom[10484] = 25'b1111111000010110110011110;
    rom[10485] = 25'b1111111000011011001000110;
    rom[10486] = 25'b1111111000011111011110000;
    rom[10487] = 25'b1111111000100011110011100;
    rom[10488] = 25'b1111111000101000001001001;
    rom[10489] = 25'b1111111000101100011110111;
    rom[10490] = 25'b1111111000110000110100110;
    rom[10491] = 25'b1111111000110101001010110;
    rom[10492] = 25'b1111111000111001100001000;
    rom[10493] = 25'b1111111000111101110111010;
    rom[10494] = 25'b1111111001000010001101101;
    rom[10495] = 25'b1111111001000110100100001;
    rom[10496] = 25'b1111111001001010111010110;
    rom[10497] = 25'b1111111001001111010001011;
    rom[10498] = 25'b1111111001010011101000001;
    rom[10499] = 25'b1111111001010111111111000;
    rom[10500] = 25'b1111111001011100010101111;
    rom[10501] = 25'b1111111001100000101100110;
    rom[10502] = 25'b1111111001100101000011110;
    rom[10503] = 25'b1111111001101001011010111;
    rom[10504] = 25'b1111111001101101110001111;
    rom[10505] = 25'b1111111001110010001000111;
    rom[10506] = 25'b1111111001110110100000000;
    rom[10507] = 25'b1111111001111010110111001;
    rom[10508] = 25'b1111111001111111001110010;
    rom[10509] = 25'b1111111010000011100101001;
    rom[10510] = 25'b1111111010000111111100010;
    rom[10511] = 25'b1111111010001100010011010;
    rom[10512] = 25'b1111111010010000101010010;
    rom[10513] = 25'b1111111010010101000001001;
    rom[10514] = 25'b1111111010011001011000000;
    rom[10515] = 25'b1111111010011101101110111;
    rom[10516] = 25'b1111111010100010000101101;
    rom[10517] = 25'b1111111010100110011100010;
    rom[10518] = 25'b1111111010101010110010110;
    rom[10519] = 25'b1111111010101111001001010;
    rom[10520] = 25'b1111111010110011011111101;
    rom[10521] = 25'b1111111010110111110101111;
    rom[10522] = 25'b1111111010111100001100000;
    rom[10523] = 25'b1111111011000000100010000;
    rom[10524] = 25'b1111111011000100110111111;
    rom[10525] = 25'b1111111011001001001101101;
    rom[10526] = 25'b1111111011001101100011010;
    rom[10527] = 25'b1111111011010001111000101;
    rom[10528] = 25'b1111111011010110001101111;
    rom[10529] = 25'b1111111011011010100011000;
    rom[10530] = 25'b1111111011011110110111111;
    rom[10531] = 25'b1111111011100011001100101;
    rom[10532] = 25'b1111111011100111100001001;
    rom[10533] = 25'b1111111011101011110101011;
    rom[10534] = 25'b1111111011110000001001101;
    rom[10535] = 25'b1111111011110100011101100;
    rom[10536] = 25'b1111111011111000110001001;
    rom[10537] = 25'b1111111011111101000100100;
    rom[10538] = 25'b1111111100000001010111110;
    rom[10539] = 25'b1111111100000101101010101;
    rom[10540] = 25'b1111111100001001111101011;
    rom[10541] = 25'b1111111100001110001111110;
    rom[10542] = 25'b1111111100010010100010000;
    rom[10543] = 25'b1111111100010110110011111;
    rom[10544] = 25'b1111111100011011000101011;
    rom[10545] = 25'b1111111100011111010110110;
    rom[10546] = 25'b1111111100100011100111110;
    rom[10547] = 25'b1111111100100111111000011;
    rom[10548] = 25'b1111111100101100001000101;
    rom[10549] = 25'b1111111100110000011000110;
    rom[10550] = 25'b1111111100110100101000100;
    rom[10551] = 25'b1111111100111000110111111;
    rom[10552] = 25'b1111111100111101000110111;
    rom[10553] = 25'b1111111101000001010101100;
    rom[10554] = 25'b1111111101000101100011111;
    rom[10555] = 25'b1111111101001001110001110;
    rom[10556] = 25'b1111111101001101111111011;
    rom[10557] = 25'b1111111101010010001100101;
    rom[10558] = 25'b1111111101010110011001100;
    rom[10559] = 25'b1111111101011010100101111;
    rom[10560] = 25'b1111111101011110110001111;
    rom[10561] = 25'b1111111101100010111101100;
    rom[10562] = 25'b1111111101100111001000110;
    rom[10563] = 25'b1111111101101011010011100;
    rom[10564] = 25'b1111111101101111011101111;
    rom[10565] = 25'b1111111101110011100111110;
    rom[10566] = 25'b1111111101110111110001010;
    rom[10567] = 25'b1111111101111011111010010;
    rom[10568] = 25'b1111111110000000000010111;
    rom[10569] = 25'b1111111110000100001011001;
    rom[10570] = 25'b1111111110001000010010110;
    rom[10571] = 25'b1111111110001100011001111;
    rom[10572] = 25'b1111111110010000100000101;
    rom[10573] = 25'b1111111110010100100110111;
    rom[10574] = 25'b1111111110011000101100101;
    rom[10575] = 25'b1111111110011100110001110;
    rom[10576] = 25'b1111111110100000110110100;
    rom[10577] = 25'b1111111110100100111010110;
    rom[10578] = 25'b1111111110101000111110100;
    rom[10579] = 25'b1111111110101101000001100;
    rom[10580] = 25'b1111111110110001000100010;
    rom[10581] = 25'b1111111110110101000110011;
    rom[10582] = 25'b1111111110111001000111110;
    rom[10583] = 25'b1111111110111101001000111;
    rom[10584] = 25'b1111111111000001001001010;
    rom[10585] = 25'b1111111111000101001001010;
    rom[10586] = 25'b1111111111001001001000100;
    rom[10587] = 25'b1111111111001101000111010;
    rom[10588] = 25'b1111111111010001000101011;
    rom[10589] = 25'b1111111111010101000011000;
    rom[10590] = 25'b1111111111011001000000000;
    rom[10591] = 25'b1111111111011100111100011;
    rom[10592] = 25'b1111111111100000111000001;
    rom[10593] = 25'b1111111111100100110011010;
    rom[10594] = 25'b1111111111101000101101111;
    rom[10595] = 25'b1111111111101100100111110;
    rom[10596] = 25'b1111111111110000100001001;
    rom[10597] = 25'b1111111111110100011001110;
    rom[10598] = 25'b1111111111111000010001110;
    rom[10599] = 25'b1111111111111100001001010;
    rom[10600] = 25'b0000000000000000000000000;
    rom[10601] = 25'b0000000000000011110110000;
    rom[10602] = 25'b0000000000000111101011011;
    rom[10603] = 25'b0000000000001011100000001;
    rom[10604] = 25'b0000000000001111010100010;
    rom[10605] = 25'b0000000000010011000111110;
    rom[10606] = 25'b0000000000010110111010011;
    rom[10607] = 25'b0000000000011010101100100;
    rom[10608] = 25'b0000000000011110011101110;
    rom[10609] = 25'b0000000000100010001110100;
    rom[10610] = 25'b0000000000100101111110100;
    rom[10611] = 25'b0000000000101001101101101;
    rom[10612] = 25'b0000000000101101011100010;
    rom[10613] = 25'b0000000000110001001001111;
    rom[10614] = 25'b0000000000110100110111001;
    rom[10615] = 25'b0000000000111000100011100;
    rom[10616] = 25'b0000000000111100001111000;
    rom[10617] = 25'b0000000000111111111001111;
    rom[10618] = 25'b0000000001000011100100001;
    rom[10619] = 25'b0000000001000111001101100;
    rom[10620] = 25'b0000000001001010110110000;
    rom[10621] = 25'b0000000001001110011101111;
    rom[10622] = 25'b0000000001010010000101000;
    rom[10623] = 25'b0000000001010101101011011;
    rom[10624] = 25'b0000000001011001010001000;
    rom[10625] = 25'b0000000001011100110101110;
    rom[10626] = 25'b0000000001100000011001101;
    rom[10627] = 25'b0000000001100011111101000;
    rom[10628] = 25'b0000000001100111011111010;
    rom[10629] = 25'b0000000001101011000001000;
    rom[10630] = 25'b0000000001101110100001110;
    rom[10631] = 25'b0000000001110010000001111;
    rom[10632] = 25'b0000000001110101100001000;
    rom[10633] = 25'b0000000001111000111111011;
    rom[10634] = 25'b0000000001111100011101000;
    rom[10635] = 25'b0000000001111111111001110;
    rom[10636] = 25'b0000000010000011010101101;
    rom[10637] = 25'b0000000010000110110000110;
    rom[10638] = 25'b0000000010001010001011000;
    rom[10639] = 25'b0000000010001101100100011;
    rom[10640] = 25'b0000000010010000111101000;
    rom[10641] = 25'b0000000010010100010100101;
    rom[10642] = 25'b0000000010010111101011100;
    rom[10643] = 25'b0000000010011011000001100;
    rom[10644] = 25'b0000000010011110010110101;
    rom[10645] = 25'b0000000010100001101010111;
    rom[10646] = 25'b0000000010100100111110011;
    rom[10647] = 25'b0000000010101000010000111;
    rom[10648] = 25'b0000000010101011100010100;
    rom[10649] = 25'b0000000010101110110011010;
    rom[10650] = 25'b0000000010110010000011001;
    rom[10651] = 25'b0000000010110101010010001;
    rom[10652] = 25'b0000000010111000100000010;
    rom[10653] = 25'b0000000010111011101101011;
    rom[10654] = 25'b0000000010111110111001110;
    rom[10655] = 25'b0000000011000010000101001;
    rom[10656] = 25'b0000000011000101001111101;
    rom[10657] = 25'b0000000011001000011001010;
    rom[10658] = 25'b0000000011001011100010000;
    rom[10659] = 25'b0000000011001110101001110;
    rom[10660] = 25'b0000000011010001110000100;
    rom[10661] = 25'b0000000011010100110110011;
    rom[10662] = 25'b0000000011010111111011011;
    rom[10663] = 25'b0000000011011010111111011;
    rom[10664] = 25'b0000000011011110000010100;
    rom[10665] = 25'b0000000011100001000100110;
    rom[10666] = 25'b0000000011100100000101111;
    rom[10667] = 25'b0000000011100111000110010;
    rom[10668] = 25'b0000000011101010000101101;
    rom[10669] = 25'b0000000011101101000100000;
    rom[10670] = 25'b0000000011110000000001011;
    rom[10671] = 25'b0000000011110010111101110;
    rom[10672] = 25'b0000000011110101111001011;
    rom[10673] = 25'b0000000011111000110011111;
    rom[10674] = 25'b0000000011111011101101011;
    rom[10675] = 25'b0000000011111110100110001;
    rom[10676] = 25'b0000000100000001011101110;
    rom[10677] = 25'b0000000100000100010100011;
    rom[10678] = 25'b0000000100000111001010000;
    rom[10679] = 25'b0000000100001001111110110;
    rom[10680] = 25'b0000000100001100110010100;
    rom[10681] = 25'b0000000100001111100101010;
    rom[10682] = 25'b0000000100010010010111000;
    rom[10683] = 25'b0000000100010101000111110;
    rom[10684] = 25'b0000000100010111110111100;
    rom[10685] = 25'b0000000100011010100110010;
    rom[10686] = 25'b0000000100011101010100000;
    rom[10687] = 25'b0000000100100000000000110;
    rom[10688] = 25'b0000000100100010101100101;
    rom[10689] = 25'b0000000100100101010111011;
    rom[10690] = 25'b0000000100101000000001001;
    rom[10691] = 25'b0000000100101010101001111;
    rom[10692] = 25'b0000000100101101010001101;
    rom[10693] = 25'b0000000100101111111000010;
    rom[10694] = 25'b0000000100110010011101111;
    rom[10695] = 25'b0000000100110101000010101;
    rom[10696] = 25'b0000000100110111100110010;
    rom[10697] = 25'b0000000100111010001000111;
    rom[10698] = 25'b0000000100111100101010100;
    rom[10699] = 25'b0000000100111111001011000;
    rom[10700] = 25'b0000000101000001101010101;
    rom[10701] = 25'b0000000101000100001001001;
    rom[10702] = 25'b0000000101000110100110100;
    rom[10703] = 25'b0000000101001001000011000;
    rom[10704] = 25'b0000000101001011011110011;
    rom[10705] = 25'b0000000101001101111000110;
    rom[10706] = 25'b0000000101010000010010000;
    rom[10707] = 25'b0000000101010010101010011;
    rom[10708] = 25'b0000000101010101000001100;
    rom[10709] = 25'b0000000101010111010111110;
    rom[10710] = 25'b0000000101011001101100111;
    rom[10711] = 25'b0000000101011100000000111;
    rom[10712] = 25'b0000000101011110010011111;
    rom[10713] = 25'b0000000101100000100110000;
    rom[10714] = 25'b0000000101100010110110111;
    rom[10715] = 25'b0000000101100101000110110;
    rom[10716] = 25'b0000000101100111010101100;
    rom[10717] = 25'b0000000101101001100011011;
    rom[10718] = 25'b0000000101101011110000000;
    rom[10719] = 25'b0000000101101101111011101;
    rom[10720] = 25'b0000000101110000000110010;
    rom[10721] = 25'b0000000101110010001111101;
    rom[10722] = 25'b0000000101110100011000001;
    rom[10723] = 25'b0000000101110110011111100;
    rom[10724] = 25'b0000000101111000100101110;
    rom[10725] = 25'b0000000101111010101011000;
    rom[10726] = 25'b0000000101111100101111001;
    rom[10727] = 25'b0000000101111110110010010;
    rom[10728] = 25'b0000000110000000110100010;
    rom[10729] = 25'b0000000110000010110101010;
    rom[10730] = 25'b0000000110000100110101001;
    rom[10731] = 25'b0000000110000110110011111;
    rom[10732] = 25'b0000000110001000110001101;
    rom[10733] = 25'b0000000110001010101110010;
    rom[10734] = 25'b0000000110001100101001111;
    rom[10735] = 25'b0000000110001110100100010;
    rom[10736] = 25'b0000000110010000011101110;
    rom[10737] = 25'b0000000110010010010110000;
    rom[10738] = 25'b0000000110010100001101011;
    rom[10739] = 25'b0000000110010110000011100;
    rom[10740] = 25'b0000000110010111111000101;
    rom[10741] = 25'b0000000110011001101100101;
    rom[10742] = 25'b0000000110011011011111100;
    rom[10743] = 25'b0000000110011101010001011;
    rom[10744] = 25'b0000000110011111000010000;
    rom[10745] = 25'b0000000110100000110001110;
    rom[10746] = 25'b0000000110100010100000011;
    rom[10747] = 25'b0000000110100100001101111;
    rom[10748] = 25'b0000000110100101111010010;
    rom[10749] = 25'b0000000110100111100101101;
    rom[10750] = 25'b0000000110101001001111111;
    rom[10751] = 25'b0000000110101010111001000;
    rom[10752] = 25'b0000000110101100100001001;
    rom[10753] = 25'b0000000110101110001000001;
    rom[10754] = 25'b0000000110101111101110000;
    rom[10755] = 25'b0000000110110001010010110;
    rom[10756] = 25'b0000000110110010110110101;
    rom[10757] = 25'b0000000110110100011001001;
    rom[10758] = 25'b0000000110110101111010110;
    rom[10759] = 25'b0000000110110111011011001;
    rom[10760] = 25'b0000000110111000111010101;
    rom[10761] = 25'b0000000110111010011000111;
    rom[10762] = 25'b0000000110111011110110000;
    rom[10763] = 25'b0000000110111101010010010;
    rom[10764] = 25'b0000000110111110101101010;
    rom[10765] = 25'b0000000111000000000111010;
    rom[10766] = 25'b0000000111000001100000001;
    rom[10767] = 25'b0000000111000010110111111;
    rom[10768] = 25'b0000000111000100001110101;
    rom[10769] = 25'b0000000111000101100100001;
    rom[10770] = 25'b0000000111000110111000110;
    rom[10771] = 25'b0000000111001000001100001;
    rom[10772] = 25'b0000000111001001011110100;
    rom[10773] = 25'b0000000111001010101111111;
    rom[10774] = 25'b0000000111001100000000000;
    rom[10775] = 25'b0000000111001101001111001;
    rom[10776] = 25'b0000000111001110011101001;
    rom[10777] = 25'b0000000111001111101010001;
    rom[10778] = 25'b0000000111010000110110000;
    rom[10779] = 25'b0000000111010010000000110;
    rom[10780] = 25'b0000000111010011001010100;
    rom[10781] = 25'b0000000111010100010011001;
    rom[10782] = 25'b0000000111010101011010110;
    rom[10783] = 25'b0000000111010110100001010;
    rom[10784] = 25'b0000000111010111100110101;
    rom[10785] = 25'b0000000111011000101011000;
    rom[10786] = 25'b0000000111011001101110010;
    rom[10787] = 25'b0000000111011010110000100;
    rom[10788] = 25'b0000000111011011110001101;
    rom[10789] = 25'b0000000111011100110001101;
    rom[10790] = 25'b0000000111011101110000101;
    rom[10791] = 25'b0000000111011110101110101;
    rom[10792] = 25'b0000000111011111101011011;
    rom[10793] = 25'b0000000111100000100111001;
    rom[10794] = 25'b0000000111100001100010000;
    rom[10795] = 25'b0000000111100010011011101;
    rom[10796] = 25'b0000000111100011010100001;
    rom[10797] = 25'b0000000111100100001011110;
    rom[10798] = 25'b0000000111100101000010001;
    rom[10799] = 25'b0000000111100101110111100;
    rom[10800] = 25'b0000000111100110101100000;
    rom[10801] = 25'b0000000111100111011111001;
    rom[10802] = 25'b0000000111101000010001100;
    rom[10803] = 25'b0000000111101001000010110;
    rom[10804] = 25'b0000000111101001110010110;
    rom[10805] = 25'b0000000111101010100001111;
    rom[10806] = 25'b0000000111101011001111111;
    rom[10807] = 25'b0000000111101011111100111;
    rom[10808] = 25'b0000000111101100101000111;
    rom[10809] = 25'b0000000111101101010011110;
    rom[10810] = 25'b0000000111101101111101101;
    rom[10811] = 25'b0000000111101110100110010;
    rom[10812] = 25'b0000000111101111001110001;
    rom[10813] = 25'b0000000111101111110100111;
    rom[10814] = 25'b0000000111110000011010100;
    rom[10815] = 25'b0000000111110000111111001;
    rom[10816] = 25'b0000000111110001100010110;
    rom[10817] = 25'b0000000111110010000101100;
    rom[10818] = 25'b0000000111110010100111000;
    rom[10819] = 25'b0000000111110011000111100;
    rom[10820] = 25'b0000000111110011100111000;
    rom[10821] = 25'b0000000111110100000101100;
    rom[10822] = 25'b0000000111110100100010111;
    rom[10823] = 25'b0000000111110100111111011;
    rom[10824] = 25'b0000000111110101011010111;
    rom[10825] = 25'b0000000111110101110101010;
    rom[10826] = 25'b0000000111110110001110101;
    rom[10827] = 25'b0000000111110110100111000;
    rom[10828] = 25'b0000000111110110111110011;
    rom[10829] = 25'b0000000111110111010100101;
    rom[10830] = 25'b0000000111110111101010000;
    rom[10831] = 25'b0000000111110111111110100;
    rom[10832] = 25'b0000000111111000010001110;
    rom[10833] = 25'b0000000111111000100100001;
    rom[10834] = 25'b0000000111111000110101011;
    rom[10835] = 25'b0000000111111001000101110;
    rom[10836] = 25'b0000000111111001010101001;
    rom[10837] = 25'b0000000111111001100011100;
    rom[10838] = 25'b0000000111111001110000111;
    rom[10839] = 25'b0000000111111001111101010;
    rom[10840] = 25'b0000000111111010001000101;
    rom[10841] = 25'b0000000111111010010011001;
    rom[10842] = 25'b0000000111111010011100100;
    rom[10843] = 25'b0000000111111010100101000;
    rom[10844] = 25'b0000000111111010101100100;
    rom[10845] = 25'b0000000111111010110011000;
    rom[10846] = 25'b0000000111111010111000101;
    rom[10847] = 25'b0000000111111010111101001;
    rom[10848] = 25'b0000000111111011000000110;
    rom[10849] = 25'b0000000111111011000011011;
    rom[10850] = 25'b0000000111111011000101001;
    rom[10851] = 25'b0000000111111011000101111;
    rom[10852] = 25'b0000000111111011000101101;
    rom[10853] = 25'b0000000111111011000100100;
    rom[10854] = 25'b0000000111111011000010011;
    rom[10855] = 25'b0000000111111010111111010;
    rom[10856] = 25'b0000000111111010111011010;
    rom[10857] = 25'b0000000111111010110110011;
    rom[10858] = 25'b0000000111111010110000011;
    rom[10859] = 25'b0000000111111010101001101;
    rom[10860] = 25'b0000000111111010100001111;
    rom[10861] = 25'b0000000111111010011001001;
    rom[10862] = 25'b0000000111111010001111100;
    rom[10863] = 25'b0000000111111010000101000;
    rom[10864] = 25'b0000000111111001111001100;
    rom[10865] = 25'b0000000111111001101101001;
    rom[10866] = 25'b0000000111111001011111111;
    rom[10867] = 25'b0000000111111001010001101;
    rom[10868] = 25'b0000000111111001000010100;
    rom[10869] = 25'b0000000111111000110010100;
    rom[10870] = 25'b0000000111111000100001100;
    rom[10871] = 25'b0000000111111000001111110;
    rom[10872] = 25'b0000000111110111111101000;
    rom[10873] = 25'b0000000111110111101001011;
    rom[10874] = 25'b0000000111110111010100111;
    rom[10875] = 25'b0000000111110110111111100;
    rom[10876] = 25'b0000000111110110101001001;
    rom[10877] = 25'b0000000111110110010010000;
    rom[10878] = 25'b0000000111110101111010000;
    rom[10879] = 25'b0000000111110101100001000;
    rom[10880] = 25'b0000000111110101000111001;
    rom[10881] = 25'b0000000111110100101100100;
    rom[10882] = 25'b0000000111110100010001000;
    rom[10883] = 25'b0000000111110011110100100;
    rom[10884] = 25'b0000000111110011010111011;
    rom[10885] = 25'b0000000111110010111001010;
    rom[10886] = 25'b0000000111110010011010010;
    rom[10887] = 25'b0000000111110001111010011;
    rom[10888] = 25'b0000000111110001011001101;
    rom[10889] = 25'b0000000111110000111000001;
    rom[10890] = 25'b0000000111110000010101111;
    rom[10891] = 25'b0000000111101111110010101;
    rom[10892] = 25'b0000000111101111001110101;
    rom[10893] = 25'b0000000111101110101001110;
    rom[10894] = 25'b0000000111101110000100001;
    rom[10895] = 25'b0000000111101101011101100;
    rom[10896] = 25'b0000000111101100110110001;
    rom[10897] = 25'b0000000111101100001110001;
    rom[10898] = 25'b0000000111101011100101000;
    rom[10899] = 25'b0000000111101010111011010;
    rom[10900] = 25'b0000000111101010010000110;
    rom[10901] = 25'b0000000111101001100101011;
    rom[10902] = 25'b0000000111101000111001001;
    rom[10903] = 25'b0000000111101000001100001;
    rom[10904] = 25'b0000000111100111011110011;
    rom[10905] = 25'b0000000111100110101111110;
    rom[10906] = 25'b0000000111100110000000100;
    rom[10907] = 25'b0000000111100101010000010;
    rom[10908] = 25'b0000000111100100011111011;
    rom[10909] = 25'b0000000111100011101101110;
    rom[10910] = 25'b0000000111100010111011010;
    rom[10911] = 25'b0000000111100010001000000;
    rom[10912] = 25'b0000000111100001010100000;
    rom[10913] = 25'b0000000111100000011111010;
    rom[10914] = 25'b0000000111011111101001111;
    rom[10915] = 25'b0000000111011110110011100;
    rom[10916] = 25'b0000000111011101111100100;
    rom[10917] = 25'b0000000111011101000100110;
    rom[10918] = 25'b0000000111011100001100010;
    rom[10919] = 25'b0000000111011011010011001;
    rom[10920] = 25'b0000000111011010011001000;
    rom[10921] = 25'b0000000111011001011110011;
    rom[10922] = 25'b0000000111011000100010111;
    rom[10923] = 25'b0000000111010111100110111;
    rom[10924] = 25'b0000000111010110101001111;
    rom[10925] = 25'b0000000111010101101100011;
    rom[10926] = 25'b0000000111010100101110001;
    rom[10927] = 25'b0000000111010011101111000;
    rom[10928] = 25'b0000000111010010101111011;
    rom[10929] = 25'b0000000111010001101110111;
    rom[10930] = 25'b0000000111010000101101111;
    rom[10931] = 25'b0000000111001111101100000;
    rom[10932] = 25'b0000000111001110101001101;
    rom[10933] = 25'b0000000111001101100110011;
    rom[10934] = 25'b0000000111001100100010101;
    rom[10935] = 25'b0000000111001011011110000;
    rom[10936] = 25'b0000000111001010011000110;
    rom[10937] = 25'b0000000111001001010011000;
    rom[10938] = 25'b0000000111001000001100100;
    rom[10939] = 25'b0000000111000111000101010;
    rom[10940] = 25'b0000000111000101111101100;
    rom[10941] = 25'b0000000111000100110101000;
    rom[10942] = 25'b0000000111000011101011111;
    rom[10943] = 25'b0000000111000010100010000;
    rom[10944] = 25'b0000000111000001010111100;
    rom[10945] = 25'b0000000111000000001100100;
    rom[10946] = 25'b0000000110111111000000110;
    rom[10947] = 25'b0000000110111101110100100;
    rom[10948] = 25'b0000000110111100100111100;
    rom[10949] = 25'b0000000110111011011010000;
    rom[10950] = 25'b0000000110111010001011110;
    rom[10951] = 25'b0000000110111000111101000;
    rom[10952] = 25'b0000000110110111101101100;
    rom[10953] = 25'b0000000110110110011101100;
    rom[10954] = 25'b0000000110110101001100111;
    rom[10955] = 25'b0000000110110011111011101;
    rom[10956] = 25'b0000000110110010101001111;
    rom[10957] = 25'b0000000110110001010111011;
    rom[10958] = 25'b0000000110110000000100100;
    rom[10959] = 25'b0000000110101110110001000;
    rom[10960] = 25'b0000000110101101011100110;
    rom[10961] = 25'b0000000110101100001000001;
    rom[10962] = 25'b0000000110101010110010111;
    rom[10963] = 25'b0000000110101001011101000;
    rom[10964] = 25'b0000000110101000000110100;
    rom[10965] = 25'b0000000110100110101111101;
    rom[10966] = 25'b0000000110100101011000001;
    rom[10967] = 25'b0000000110100100000000000;
    rom[10968] = 25'b0000000110100010100111100;
    rom[10969] = 25'b0000000110100001001110011;
    rom[10970] = 25'b0000000110011111110100101;
    rom[10971] = 25'b0000000110011110011010100;
    rom[10972] = 25'b0000000110011100111111110;
    rom[10973] = 25'b0000000110011011100100100;
    rom[10974] = 25'b0000000110011010001000110;
    rom[10975] = 25'b0000000110011000101100100;
    rom[10976] = 25'b0000000110010111001111101;
    rom[10977] = 25'b0000000110010101110010011;
    rom[10978] = 25'b0000000110010100010100100;
    rom[10979] = 25'b0000000110010010110110010;
    rom[10980] = 25'b0000000110010001010111100;
    rom[10981] = 25'b0000000110001111111000010;
    rom[10982] = 25'b0000000110001110011000100;
    rom[10983] = 25'b0000000110001100111000010;
    rom[10984] = 25'b0000000110001011010111100;
    rom[10985] = 25'b0000000110001001110110011;
    rom[10986] = 25'b0000000110001000010100110;
    rom[10987] = 25'b0000000110000110110010101;
    rom[10988] = 25'b0000000110000101010000001;
    rom[10989] = 25'b0000000110000011101101000;
    rom[10990] = 25'b0000000110000010001001101;
    rom[10991] = 25'b0000000110000000100101101;
    rom[10992] = 25'b0000000101111111000001011;
    rom[10993] = 25'b0000000101111101011100100;
    rom[10994] = 25'b0000000101111011110111010;
    rom[10995] = 25'b0000000101111010010001101;
    rom[10996] = 25'b0000000101111000101011100;
    rom[10997] = 25'b0000000101110111000101000;
    rom[10998] = 25'b0000000101110101011110000;
    rom[10999] = 25'b0000000101110011110110101;
    rom[11000] = 25'b0000000101110010001111000;
    rom[11001] = 25'b0000000101110000100110111;
    rom[11002] = 25'b0000000101101110111110011;
    rom[11003] = 25'b0000000101101101010101011;
    rom[11004] = 25'b0000000101101011101100000;
    rom[11005] = 25'b0000000101101010000010010;
    rom[11006] = 25'b0000000101101000011000001;
    rom[11007] = 25'b0000000101100110101101110;
    rom[11008] = 25'b0000000101100101000010111;
    rom[11009] = 25'b0000000101100011010111101;
    rom[11010] = 25'b0000000101100001101100000;
    rom[11011] = 25'b0000000101100000000000001;
    rom[11012] = 25'b0000000101011110010011110;
    rom[11013] = 25'b0000000101011100100111001;
    rom[11014] = 25'b0000000101011010111010010;
    rom[11015] = 25'b0000000101011001001100110;
    rom[11016] = 25'b0000000101010111011111001;
    rom[11017] = 25'b0000000101010101110001000;
    rom[11018] = 25'b0000000101010100000010110;
    rom[11019] = 25'b0000000101010010010100000;
    rom[11020] = 25'b0000000101010000100101000;
    rom[11021] = 25'b0000000101001110110101110;
    rom[11022] = 25'b0000000101001101000110001;
    rom[11023] = 25'b0000000101001011010110001;
    rom[11024] = 25'b0000000101001001100101111;
    rom[11025] = 25'b0000000101000111110101010;
    rom[11026] = 25'b0000000101000110000100011;
    rom[11027] = 25'b0000000101000100010011010;
    rom[11028] = 25'b0000000101000010100001111;
    rom[11029] = 25'b0000000101000000110000001;
    rom[11030] = 25'b0000000100111110111110001;
    rom[11031] = 25'b0000000100111101001011111;
    rom[11032] = 25'b0000000100111011011001010;
    rom[11033] = 25'b0000000100111001100110011;
    rom[11034] = 25'b0000000100110111110011011;
    rom[11035] = 25'b0000000100110110000000000;
    rom[11036] = 25'b0000000100110100001100100;
    rom[11037] = 25'b0000000100110010011000101;
    rom[11038] = 25'b0000000100110000100100100;
    rom[11039] = 25'b0000000100101110110000001;
    rom[11040] = 25'b0000000100101100111011101;
    rom[11041] = 25'b0000000100101011000110110;
    rom[11042] = 25'b0000000100101001010001101;
    rom[11043] = 25'b0000000100100111011100011;
    rom[11044] = 25'b0000000100100101100111000;
    rom[11045] = 25'b0000000100100011110001010;
    rom[11046] = 25'b0000000100100001111011010;
    rom[11047] = 25'b0000000100100000000101001;
    rom[11048] = 25'b0000000100011110001110111;
    rom[11049] = 25'b0000000100011100011000010;
    rom[11050] = 25'b0000000100011010100001100;
    rom[11051] = 25'b0000000100011000101010101;
    rom[11052] = 25'b0000000100010110110011100;
    rom[11053] = 25'b0000000100010100111100001;
    rom[11054] = 25'b0000000100010011000100101;
    rom[11055] = 25'b0000000100010001001101000;
    rom[11056] = 25'b0000000100001111010101010;
    rom[11057] = 25'b0000000100001101011101001;
    rom[11058] = 25'b0000000100001011100100111;
    rom[11059] = 25'b0000000100001001101100110;
    rom[11060] = 25'b0000000100000111110100001;
    rom[11061] = 25'b0000000100000101111011100;
    rom[11062] = 25'b0000000100000100000010110;
    rom[11063] = 25'b0000000100000010001001111;
    rom[11064] = 25'b0000000100000000010000110;
    rom[11065] = 25'b0000000011111110010111100;
    rom[11066] = 25'b0000000011111100011110001;
    rom[11067] = 25'b0000000011111010100100110;
    rom[11068] = 25'b0000000011111000101011001;
    rom[11069] = 25'b0000000011110110110001011;
    rom[11070] = 25'b0000000011110100110111100;
    rom[11071] = 25'b0000000011110010111101101;
    rom[11072] = 25'b0000000011110001000011100;
    rom[11073] = 25'b0000000011101111001001011;
    rom[11074] = 25'b0000000011101101001111001;
    rom[11075] = 25'b0000000011101011010100110;
    rom[11076] = 25'b0000000011101001011010010;
    rom[11077] = 25'b0000000011100111011111111;
    rom[11078] = 25'b0000000011100101100101001;
    rom[11079] = 25'b0000000011100011101010100;
    rom[11080] = 25'b0000000011100001101111101;
    rom[11081] = 25'b0000000011011111110100110;
    rom[11082] = 25'b0000000011011101111001111;
    rom[11083] = 25'b0000000011011011111110111;
    rom[11084] = 25'b0000000011011010000011111;
    rom[11085] = 25'b0000000011011000001000110;
    rom[11086] = 25'b0000000011010110001101101;
    rom[11087] = 25'b0000000011010100010010011;
    rom[11088] = 25'b0000000011010010010111001;
    rom[11089] = 25'b0000000011010000011011111;
    rom[11090] = 25'b0000000011001110100000100;
    rom[11091] = 25'b0000000011001100100101001;
    rom[11092] = 25'b0000000011001010101001110;
    rom[11093] = 25'b0000000011001000101110010;
    rom[11094] = 25'b0000000011000110110010111;
    rom[11095] = 25'b0000000011000100110111011;
    rom[11096] = 25'b0000000011000010111011111;
    rom[11097] = 25'b0000000011000001000000100;
    rom[11098] = 25'b0000000010111111000100111;
    rom[11099] = 25'b0000000010111101001001011;
    rom[11100] = 25'b0000000010111011001101111;
    rom[11101] = 25'b0000000010111001010010011;
    rom[11102] = 25'b0000000010110111010110111;
    rom[11103] = 25'b0000000010110101011011011;
    rom[11104] = 25'b0000000010110011011111111;
    rom[11105] = 25'b0000000010110001100100100;
    rom[11106] = 25'b0000000010101111101001001;
    rom[11107] = 25'b0000000010101101101101101;
    rom[11108] = 25'b0000000010101011110010010;
    rom[11109] = 25'b0000000010101001110110111;
    rom[11110] = 25'b0000000010100111111011101;
    rom[11111] = 25'b0000000010100110000000011;
    rom[11112] = 25'b0000000010100100000101000;
    rom[11113] = 25'b0000000010100010001001111;
    rom[11114] = 25'b0000000010100000001110111;
    rom[11115] = 25'b0000000010011110010011110;
    rom[11116] = 25'b0000000010011100011000110;
    rom[11117] = 25'b0000000010011010011101110;
    rom[11118] = 25'b0000000010011000100010110;
    rom[11119] = 25'b0000000010010110101000000;
    rom[11120] = 25'b0000000010010100101101010;
    rom[11121] = 25'b0000000010010010110010100;
    rom[11122] = 25'b0000000010010000111000000;
    rom[11123] = 25'b0000000010001110111101011;
    rom[11124] = 25'b0000000010001101000011000;
    rom[11125] = 25'b0000000010001011001000101;
    rom[11126] = 25'b0000000010001001001110011;
    rom[11127] = 25'b0000000010000111010100010;
    rom[11128] = 25'b0000000010000101011010001;
    rom[11129] = 25'b0000000010000011100000001;
    rom[11130] = 25'b0000000010000001100110011;
    rom[11131] = 25'b0000000001111111101100101;
    rom[11132] = 25'b0000000001111101110011000;
    rom[11133] = 25'b0000000001111011111001100;
    rom[11134] = 25'b0000000001111010000000000;
    rom[11135] = 25'b0000000001111000000110110;
    rom[11136] = 25'b0000000001110110001101100;
    rom[11137] = 25'b0000000001110100010100100;
    rom[11138] = 25'b0000000001110010011011101;
    rom[11139] = 25'b0000000001110000100010111;
    rom[11140] = 25'b0000000001101110101010011;
    rom[11141] = 25'b0000000001101100110001110;
    rom[11142] = 25'b0000000001101010111001100;
    rom[11143] = 25'b0000000001101001000001011;
    rom[11144] = 25'b0000000001100111001001010;
    rom[11145] = 25'b0000000001100101010001011;
    rom[11146] = 25'b0000000001100011011001101;
    rom[11147] = 25'b0000000001100001100010001;
    rom[11148] = 25'b0000000001011111101010110;
    rom[11149] = 25'b0000000001011101110011100;
    rom[11150] = 25'b0000000001011011111100011;
    rom[11151] = 25'b0000000001011010000101101;
    rom[11152] = 25'b0000000001011000001110111;
    rom[11153] = 25'b0000000001010110011000011;
    rom[11154] = 25'b0000000001010100100010000;
    rom[11155] = 25'b0000000001010010101011111;
    rom[11156] = 25'b0000000001010000110101111;
    rom[11157] = 25'b0000000001001111000000000;
    rom[11158] = 25'b0000000001001101001010100;
    rom[11159] = 25'b0000000001001011010101001;
    rom[11160] = 25'b0000000001001001011111111;
    rom[11161] = 25'b0000000001000111101011000;
    rom[11162] = 25'b0000000001000101110110001;
    rom[11163] = 25'b0000000001000100000001101;
    rom[11164] = 25'b0000000001000010001101010;
    rom[11165] = 25'b0000000001000000011001001;
    rom[11166] = 25'b0000000000111110100101001;
    rom[11167] = 25'b0000000000111100110001100;
    rom[11168] = 25'b0000000000111010111110000;
    rom[11169] = 25'b0000000000111001001010110;
    rom[11170] = 25'b0000000000110111010111110;
    rom[11171] = 25'b0000000000110101100100111;
    rom[11172] = 25'b0000000000110011110010011;
    rom[11173] = 25'b0000000000110010000000000;
    rom[11174] = 25'b0000000000110000001110000;
    rom[11175] = 25'b0000000000101110011100001;
    rom[11176] = 25'b0000000000101100101010101;
    rom[11177] = 25'b0000000000101010111001001;
    rom[11178] = 25'b0000000000101001001000001;
    rom[11179] = 25'b0000000000100111010111010;
    rom[11180] = 25'b0000000000100101100110101;
    rom[11181] = 25'b0000000000100011110110011;
    rom[11182] = 25'b0000000000100010000110011;
    rom[11183] = 25'b0000000000100000010110100;
    rom[11184] = 25'b0000000000011110100111000;
    rom[11185] = 25'b0000000000011100110111101;
    rom[11186] = 25'b0000000000011011001000101;
    rom[11187] = 25'b0000000000011001011010000;
    rom[11188] = 25'b0000000000010111101011100;
    rom[11189] = 25'b0000000000010101111101011;
    rom[11190] = 25'b0000000000010100001111101;
    rom[11191] = 25'b0000000000010010100010000;
    rom[11192] = 25'b0000000000010000110100101;
    rom[11193] = 25'b0000000000001111000111101;
    rom[11194] = 25'b0000000000001101011010111;
    rom[11195] = 25'b0000000000001011101110100;
    rom[11196] = 25'b0000000000001010000010010;
    rom[11197] = 25'b0000000000001000010110100;
    rom[11198] = 25'b0000000000000110101011000;
    rom[11199] = 25'b0000000000000100111111110;
    rom[11200] = 25'b0000000000000011010100110;
    rom[11201] = 25'b0000000000000001101010001;
    rom[11202] = 25'b0000000000000000000000000;
    rom[11203] = 25'b1111111111111110010110000;
    rom[11204] = 25'b1111111111111100101100011;
    rom[11205] = 25'b1111111111111011000011000;
    rom[11206] = 25'b1111111111111001011010000;
    rom[11207] = 25'b1111111111110111110001010;
    rom[11208] = 25'b1111111111110110001000111;
    rom[11209] = 25'b1111111111110100100000110;
    rom[11210] = 25'b1111111111110010111001000;
    rom[11211] = 25'b1111111111110001010001101;
    rom[11212] = 25'b1111111111101111101010101;
    rom[11213] = 25'b1111111111101110000011111;
    rom[11214] = 25'b1111111111101100011101011;
    rom[11215] = 25'b1111111111101010110111011;
    rom[11216] = 25'b1111111111101001010001110;
    rom[11217] = 25'b1111111111100111101100010;
    rom[11218] = 25'b1111111111100110000111010;
    rom[11219] = 25'b1111111111100100100010101;
    rom[11220] = 25'b1111111111100010111110010;
    rom[11221] = 25'b1111111111100001011010010;
    rom[11222] = 25'b1111111111011111110110101;
    rom[11223] = 25'b1111111111011110010011011;
    rom[11224] = 25'b1111111111011100110000011;
    rom[11225] = 25'b1111111111011011001101111;
    rom[11226] = 25'b1111111111011001101011110;
    rom[11227] = 25'b1111111111011000001001111;
    rom[11228] = 25'b1111111111010110101000100;
    rom[11229] = 25'b1111111111010101000111010;
    rom[11230] = 25'b1111111111010011100110100;
    rom[11231] = 25'b1111111111010010000110010;
    rom[11232] = 25'b1111111111010000100110010;
    rom[11233] = 25'b1111111111001111000110101;
    rom[11234] = 25'b1111111111001101100111011;
    rom[11235] = 25'b1111111111001100001000100;
    rom[11236] = 25'b1111111111001010101010000;
    rom[11237] = 25'b1111111111001001001100000;
    rom[11238] = 25'b1111111111000111101110001;
    rom[11239] = 25'b1111111111000110010001000;
    rom[11240] = 25'b1111111111000100110011111;
    rom[11241] = 25'b1111111111000011010111011;
    rom[11242] = 25'b1111111111000001111011010;
    rom[11243] = 25'b1111111111000000011111011;
    rom[11244] = 25'b1111111110111111000100001;
    rom[11245] = 25'b1111111110111101101001001;
    rom[11246] = 25'b1111111110111100001110100;
    rom[11247] = 25'b1111111110111010110100011;
    rom[11248] = 25'b1111111110111001011010100;
    rom[11249] = 25'b1111111110111000000001001;
    rom[11250] = 25'b1111111110110110101000001;
    rom[11251] = 25'b1111111110110101001111101;
    rom[11252] = 25'b1111111110110011110111011;
    rom[11253] = 25'b1111111110110010011111101;
    rom[11254] = 25'b1111111110110001001000010;
    rom[11255] = 25'b1111111110101111110001010;
    rom[11256] = 25'b1111111110101110011010110;
    rom[11257] = 25'b1111111110101101000100101;
    rom[11258] = 25'b1111111110101011101110111;
    rom[11259] = 25'b1111111110101010011001100;
    rom[11260] = 25'b1111111110101001000100110;
    rom[11261] = 25'b1111111110100111110000010;
    rom[11262] = 25'b1111111110100110011100001;
    rom[11263] = 25'b1111111110100101001000100;
    rom[11264] = 25'b1111111110100011110101010;
    rom[11265] = 25'b1111111110100010100010100;
    rom[11266] = 25'b1111111110100001010000010;
    rom[11267] = 25'b1111111110011111111110010;
    rom[11268] = 25'b1111111110011110101100110;
    rom[11269] = 25'b1111111110011101011011101;
    rom[11270] = 25'b1111111110011100001011000;
    rom[11271] = 25'b1111111110011010111010110;
    rom[11272] = 25'b1111111110011001101011000;
    rom[11273] = 25'b1111111110011000011011101;
    rom[11274] = 25'b1111111110010111001100110;
    rom[11275] = 25'b1111111110010101111110010;
    rom[11276] = 25'b1111111110010100110000001;
    rom[11277] = 25'b1111111110010011100010100;
    rom[11278] = 25'b1111111110010010010101010;
    rom[11279] = 25'b1111111110010001001000100;
    rom[11280] = 25'b1111111110001111111100011;
    rom[11281] = 25'b1111111110001110110000011;
    rom[11282] = 25'b1111111110001101100101000;
    rom[11283] = 25'b1111111110001100011010001;
    rom[11284] = 25'b1111111110001011001111101;
    rom[11285] = 25'b1111111110001010000101100;
    rom[11286] = 25'b1111111110001000111011110;
    rom[11287] = 25'b1111111110000111110010101;
    rom[11288] = 25'b1111111110000110101001111;
    rom[11289] = 25'b1111111110000101100001100;
    rom[11290] = 25'b1111111110000100011001101;
    rom[11291] = 25'b1111111110000011010010011;
    rom[11292] = 25'b1111111110000010001011011;
    rom[11293] = 25'b1111111110000001000100111;
    rom[11294] = 25'b1111111101111111111110110;
    rom[11295] = 25'b1111111101111110111001010;
    rom[11296] = 25'b1111111101111101110100001;
    rom[11297] = 25'b1111111101111100101111100;
    rom[11298] = 25'b1111111101111011101011010;
    rom[11299] = 25'b1111111101111010100111011;
    rom[11300] = 25'b1111111101111001100100001;
    rom[11301] = 25'b1111111101111000100001010;
    rom[11302] = 25'b1111111101110111011110111;
    rom[11303] = 25'b1111111101110110011101000;
    rom[11304] = 25'b1111111101110101011011100;
    rom[11305] = 25'b1111111101110100011010011;
    rom[11306] = 25'b1111111101110011011001111;
    rom[11307] = 25'b1111111101110010011001110;
    rom[11308] = 25'b1111111101110001011010001;
    rom[11309] = 25'b1111111101110000011011000;
    rom[11310] = 25'b1111111101101111011100010;
    rom[11311] = 25'b1111111101101110011110000;
    rom[11312] = 25'b1111111101101101100000010;
    rom[11313] = 25'b1111111101101100100010111;
    rom[11314] = 25'b1111111101101011100110000;
    rom[11315] = 25'b1111111101101010101001101;
    rom[11316] = 25'b1111111101101001101101110;
    rom[11317] = 25'b1111111101101000110010011;
    rom[11318] = 25'b1111111101100111110111011;
    rom[11319] = 25'b1111111101100110111100110;
    rom[11320] = 25'b1111111101100110000010110;
    rom[11321] = 25'b1111111101100101001001001;
    rom[11322] = 25'b1111111101100100010000000;
    rom[11323] = 25'b1111111101100011010111011;
    rom[11324] = 25'b1111111101100010011111010;
    rom[11325] = 25'b1111111101100001100111100;
    rom[11326] = 25'b1111111101100000110000010;
    rom[11327] = 25'b1111111101011111111001100;
    rom[11328] = 25'b1111111101011111000011001;
    rom[11329] = 25'b1111111101011110001101011;
    rom[11330] = 25'b1111111101011101011000000;
    rom[11331] = 25'b1111111101011100100011000;
    rom[11332] = 25'b1111111101011011101110101;
    rom[11333] = 25'b1111111101011010111010110;
    rom[11334] = 25'b1111111101011010000111001;
    rom[11335] = 25'b1111111101011001010100001;
    rom[11336] = 25'b1111111101011000100001101;
    rom[11337] = 25'b1111111101010111101111101;
    rom[11338] = 25'b1111111101010110111110000;
    rom[11339] = 25'b1111111101010110001100111;
    rom[11340] = 25'b1111111101010101011100010;
    rom[11341] = 25'b1111111101010100101100000;
    rom[11342] = 25'b1111111101010011111100011;
    rom[11343] = 25'b1111111101010011001101001;
    rom[11344] = 25'b1111111101010010011110011;
    rom[11345] = 25'b1111111101010001110000000;
    rom[11346] = 25'b1111111101010001000010001;
    rom[11347] = 25'b1111111101010000010100111;
    rom[11348] = 25'b1111111101001111101000000;
    rom[11349] = 25'b1111111101001110111011101;
    rom[11350] = 25'b1111111101001110001111101;
    rom[11351] = 25'b1111111101001101100100010;
    rom[11352] = 25'b1111111101001100111001010;
    rom[11353] = 25'b1111111101001100001110110;
    rom[11354] = 25'b1111111101001011100100101;
    rom[11355] = 25'b1111111101001010111011000;
    rom[11356] = 25'b1111111101001010010001111;
    rom[11357] = 25'b1111111101001001101001010;
    rom[11358] = 25'b1111111101001001000001001;
    rom[11359] = 25'b1111111101001000011001100;
    rom[11360] = 25'b1111111101000111110010010;
    rom[11361] = 25'b1111111101000111001011100;
    rom[11362] = 25'b1111111101000110100101001;
    rom[11363] = 25'b1111111101000101111111011;
    rom[11364] = 25'b1111111101000101011010000;
    rom[11365] = 25'b1111111101000100110101010;
    rom[11366] = 25'b1111111101000100010000110;
    rom[11367] = 25'b1111111101000011101100110;
    rom[11368] = 25'b1111111101000011001001010;
    rom[11369] = 25'b1111111101000010100110011;
    rom[11370] = 25'b1111111101000010000011110;
    rom[11371] = 25'b1111111101000001100001110;
    rom[11372] = 25'b1111111101000001000000001;
    rom[11373] = 25'b1111111101000000011111000;
    rom[11374] = 25'b1111111100111111111110011;
    rom[11375] = 25'b1111111100111111011110001;
    rom[11376] = 25'b1111111100111110111110011;
    rom[11377] = 25'b1111111100111110011111001;
    rom[11378] = 25'b1111111100111110000000010;
    rom[11379] = 25'b1111111100111101100010000;
    rom[11380] = 25'b1111111100111101000100001;
    rom[11381] = 25'b1111111100111100100110101;
    rom[11382] = 25'b1111111100111100001001101;
    rom[11383] = 25'b1111111100111011101101001;
    rom[11384] = 25'b1111111100111011010001001;
    rom[11385] = 25'b1111111100111010110101100;
    rom[11386] = 25'b1111111100111010011010011;
    rom[11387] = 25'b1111111100111001111111110;
    rom[11388] = 25'b1111111100111001100101101;
    rom[11389] = 25'b1111111100111001001011111;
    rom[11390] = 25'b1111111100111000110010100;
    rom[11391] = 25'b1111111100111000011001101;
    rom[11392] = 25'b1111111100111000000001011;
    rom[11393] = 25'b1111111100110111101001011;
    rom[11394] = 25'b1111111100110111010010000;
    rom[11395] = 25'b1111111100110110111011000;
    rom[11396] = 25'b1111111100110110100100011;
    rom[11397] = 25'b1111111100110110001110010;
    rom[11398] = 25'b1111111100110101111000110;
    rom[11399] = 25'b1111111100110101100011100;
    rom[11400] = 25'b1111111100110101001110110;
    rom[11401] = 25'b1111111100110100111010011;
    rom[11402] = 25'b1111111100110100100110101;
    rom[11403] = 25'b1111111100110100010011001;
    rom[11404] = 25'b1111111100110100000000010;
    rom[11405] = 25'b1111111100110011101101110;
    rom[11406] = 25'b1111111100110011011011110;
    rom[11407] = 25'b1111111100110011001010001;
    rom[11408] = 25'b1111111100110010111000111;
    rom[11409] = 25'b1111111100110010101000010;
    rom[11410] = 25'b1111111100110010011000000;
    rom[11411] = 25'b1111111100110010001000001;
    rom[11412] = 25'b1111111100110001111000110;
    rom[11413] = 25'b1111111100110001101001110;
    rom[11414] = 25'b1111111100110001011011010;
    rom[11415] = 25'b1111111100110001001101001;
    rom[11416] = 25'b1111111100110000111111100;
    rom[11417] = 25'b1111111100110000110010011;
    rom[11418] = 25'b1111111100110000100101101;
    rom[11419] = 25'b1111111100110000011001010;
    rom[11420] = 25'b1111111100110000001101011;
    rom[11421] = 25'b1111111100110000000001111;
    rom[11422] = 25'b1111111100101111110110111;
    rom[11423] = 25'b1111111100101111101100010;
    rom[11424] = 25'b1111111100101111100010001;
    rom[11425] = 25'b1111111100101111011000011;
    rom[11426] = 25'b1111111100101111001111000;
    rom[11427] = 25'b1111111100101111000110010;
    rom[11428] = 25'b1111111100101110111101110;
    rom[11429] = 25'b1111111100101110110101101;
    rom[11430] = 25'b1111111100101110101110001;
    rom[11431] = 25'b1111111100101110100110111;
    rom[11432] = 25'b1111111100101110100000001;
    rom[11433] = 25'b1111111100101110011001110;
    rom[11434] = 25'b1111111100101110010011111;
    rom[11435] = 25'b1111111100101110001110011;
    rom[11436] = 25'b1111111100101110001001010;
    rom[11437] = 25'b1111111100101110000100101;
    rom[11438] = 25'b1111111100101110000000011;
    rom[11439] = 25'b1111111100101101111100100;
    rom[11440] = 25'b1111111100101101111001001;
    rom[11441] = 25'b1111111100101101110110000;
    rom[11442] = 25'b1111111100101101110011100;
    rom[11443] = 25'b1111111100101101110001010;
    rom[11444] = 25'b1111111100101101101111100;
    rom[11445] = 25'b1111111100101101101110001;
    rom[11446] = 25'b1111111100101101101101001;
    rom[11447] = 25'b1111111100101101101100101;
    rom[11448] = 25'b1111111100101101101100011;
    rom[11449] = 25'b1111111100101101101100101;
    rom[11450] = 25'b1111111100101101101101010;
    rom[11451] = 25'b1111111100101101101110010;
    rom[11452] = 25'b1111111100101101101111110;
    rom[11453] = 25'b1111111100101101110001101;
    rom[11454] = 25'b1111111100101101110011111;
    rom[11455] = 25'b1111111100101101110110100;
    rom[11456] = 25'b1111111100101101111001100;
    rom[11457] = 25'b1111111100101101111100111;
    rom[11458] = 25'b1111111100101110000000101;
    rom[11459] = 25'b1111111100101110000100111;
    rom[11460] = 25'b1111111100101110001001011;
    rom[11461] = 25'b1111111100101110001110011;
    rom[11462] = 25'b1111111100101110010011111;
    rom[11463] = 25'b1111111100101110011001101;
    rom[11464] = 25'b1111111100101110011111101;
    rom[11465] = 25'b1111111100101110100110001;
    rom[11466] = 25'b1111111100101110101101000;
    rom[11467] = 25'b1111111100101110110100010;
    rom[11468] = 25'b1111111100101110111011111;
    rom[11469] = 25'b1111111100101111000011111;
    rom[11470] = 25'b1111111100101111001100010;
    rom[11471] = 25'b1111111100101111010101001;
    rom[11472] = 25'b1111111100101111011110010;
    rom[11473] = 25'b1111111100101111100111110;
    rom[11474] = 25'b1111111100101111110001101;
    rom[11475] = 25'b1111111100101111111011110;
    rom[11476] = 25'b1111111100110000000110011;
    rom[11477] = 25'b1111111100110000010001011;
    rom[11478] = 25'b1111111100110000011100110;
    rom[11479] = 25'b1111111100110000101000100;
    rom[11480] = 25'b1111111100110000110100100;
    rom[11481] = 25'b1111111100110001000000111;
    rom[11482] = 25'b1111111100110001001101101;
    rom[11483] = 25'b1111111100110001011010111;
    rom[11484] = 25'b1111111100110001101000011;
    rom[11485] = 25'b1111111100110001110110001;
    rom[11486] = 25'b1111111100110010000100010;
    rom[11487] = 25'b1111111100110010010010111;
    rom[11488] = 25'b1111111100110010100001110;
    rom[11489] = 25'b1111111100110010110001000;
    rom[11490] = 25'b1111111100110011000000101;
    rom[11491] = 25'b1111111100110011010000100;
    rom[11492] = 25'b1111111100110011100000110;
    rom[11493] = 25'b1111111100110011110001011;
    rom[11494] = 25'b1111111100110100000010010;
    rom[11495] = 25'b1111111100110100010011101;
    rom[11496] = 25'b1111111100110100100101001;
    rom[11497] = 25'b1111111100110100110111001;
    rom[11498] = 25'b1111111100110101001001011;
    rom[11499] = 25'b1111111100110101011100000;
    rom[11500] = 25'b1111111100110101101111000;
    rom[11501] = 25'b1111111100110110000010010;
    rom[11502] = 25'b1111111100110110010101111;
    rom[11503] = 25'b1111111100110110101001111;
    rom[11504] = 25'b1111111100110110111110000;
    rom[11505] = 25'b1111111100110111010010101;
    rom[11506] = 25'b1111111100110111100111100;
    rom[11507] = 25'b1111111100110111111100110;
    rom[11508] = 25'b1111111100111000010010010;
    rom[11509] = 25'b1111111100111000101000001;
    rom[11510] = 25'b1111111100111000111110010;
    rom[11511] = 25'b1111111100111001010100101;
    rom[11512] = 25'b1111111100111001101011100;
    rom[11513] = 25'b1111111100111010000010101;
    rom[11514] = 25'b1111111100111010011010000;
    rom[11515] = 25'b1111111100111010110001110;
    rom[11516] = 25'b1111111100111011001001110;
    rom[11517] = 25'b1111111100111011100010000;
    rom[11518] = 25'b1111111100111011111010101;
    rom[11519] = 25'b1111111100111100010011100;
    rom[11520] = 25'b1111111100111100101100110;
    rom[11521] = 25'b1111111100111101000110010;
    rom[11522] = 25'b1111111100111101100000000;
    rom[11523] = 25'b1111111100111101111010001;
    rom[11524] = 25'b1111111100111110010100100;
    rom[11525] = 25'b1111111100111110101111001;
    rom[11526] = 25'b1111111100111111001010000;
    rom[11527] = 25'b1111111100111111100101010;
    rom[11528] = 25'b1111111101000000000000110;
    rom[11529] = 25'b1111111101000000011100101;
    rom[11530] = 25'b1111111101000000111000110;
    rom[11531] = 25'b1111111101000001010101000;
    rom[11532] = 25'b1111111101000001110001110;
    rom[11533] = 25'b1111111101000010001110101;
    rom[11534] = 25'b1111111101000010101011110;
    rom[11535] = 25'b1111111101000011001001010;
    rom[11536] = 25'b1111111101000011100111000;
    rom[11537] = 25'b1111111101000100000101000;
    rom[11538] = 25'b1111111101000100100011001;
    rom[11539] = 25'b1111111101000101000001101;
    rom[11540] = 25'b1111111101000101100000100;
    rom[11541] = 25'b1111111101000101111111100;
    rom[11542] = 25'b1111111101000110011110110;
    rom[11543] = 25'b1111111101000110111110011;
    rom[11544] = 25'b1111111101000111011110001;
    rom[11545] = 25'b1111111101000111111110010;
    rom[11546] = 25'b1111111101001000011110100;
    rom[11547] = 25'b1111111101001000111111001;
    rom[11548] = 25'b1111111101001001100000000;
    rom[11549] = 25'b1111111101001010000001000;
    rom[11550] = 25'b1111111101001010100010011;
    rom[11551] = 25'b1111111101001011000011111;
    rom[11552] = 25'b1111111101001011100101101;
    rom[11553] = 25'b1111111101001100000111110;
    rom[11554] = 25'b1111111101001100101010000;
    rom[11555] = 25'b1111111101001101001100100;
    rom[11556] = 25'b1111111101001101101111010;
    rom[11557] = 25'b1111111101001110010010010;
    rom[11558] = 25'b1111111101001110110101011;
    rom[11559] = 25'b1111111101001111011000111;
    rom[11560] = 25'b1111111101001111111100100;
    rom[11561] = 25'b1111111101010000100000100;
    rom[11562] = 25'b1111111101010001000100100;
    rom[11563] = 25'b1111111101010001101000111;
    rom[11564] = 25'b1111111101010010001101100;
    rom[11565] = 25'b1111111101010010110010010;
    rom[11566] = 25'b1111111101010011010111010;
    rom[11567] = 25'b1111111101010011111100011;
    rom[11568] = 25'b1111111101010100100001111;
    rom[11569] = 25'b1111111101010101000111100;
    rom[11570] = 25'b1111111101010101101101010;
    rom[11571] = 25'b1111111101010110010011010;
    rom[11572] = 25'b1111111101010110111001100;
    rom[11573] = 25'b1111111101010111100000000;
    rom[11574] = 25'b1111111101011000000110101;
    rom[11575] = 25'b1111111101011000101101100;
    rom[11576] = 25'b1111111101011001010100101;
    rom[11577] = 25'b1111111101011001111011110;
    rom[11578] = 25'b1111111101011010100011010;
    rom[11579] = 25'b1111111101011011001010111;
    rom[11580] = 25'b1111111101011011110010110;
    rom[11581] = 25'b1111111101011100011010110;
    rom[11582] = 25'b1111111101011101000011000;
    rom[11583] = 25'b1111111101011101101011011;
    rom[11584] = 25'b1111111101011110010011111;
    rom[11585] = 25'b1111111101011110111100110;
    rom[11586] = 25'b1111111101011111100101101;
    rom[11587] = 25'b1111111101100000001110110;
    rom[11588] = 25'b1111111101100000111000001;
    rom[11589] = 25'b1111111101100001100001100;
    rom[11590] = 25'b1111111101100010001011001;
    rom[11591] = 25'b1111111101100010110101000;
    rom[11592] = 25'b1111111101100011011111000;
    rom[11593] = 25'b1111111101100100001001001;
    rom[11594] = 25'b1111111101100100110011011;
    rom[11595] = 25'b1111111101100101011101111;
    rom[11596] = 25'b1111111101100110001000100;
    rom[11597] = 25'b1111111101100110110011010;
    rom[11598] = 25'b1111111101100111011110010;
    rom[11599] = 25'b1111111101101000001001011;
    rom[11600] = 25'b1111111101101000110100101;
    rom[11601] = 25'b1111111101101001100000000;
    rom[11602] = 25'b1111111101101010001011101;
    rom[11603] = 25'b1111111101101010110111011;
    rom[11604] = 25'b1111111101101011100011010;
    rom[11605] = 25'b1111111101101100001111010;
    rom[11606] = 25'b1111111101101100111011100;
    rom[11607] = 25'b1111111101101101100111110;
    rom[11608] = 25'b1111111101101110010100010;
    rom[11609] = 25'b1111111101101111000000110;
    rom[11610] = 25'b1111111101101111101101100;
    rom[11611] = 25'b1111111101110000011010011;
    rom[11612] = 25'b1111111101110001000111011;
    rom[11613] = 25'b1111111101110001110100100;
    rom[11614] = 25'b1111111101110010100001110;
    rom[11615] = 25'b1111111101110011001111001;
    rom[11616] = 25'b1111111101110011111100101;
    rom[11617] = 25'b1111111101110100101010010;
    rom[11618] = 25'b1111111101110101011000000;
    rom[11619] = 25'b1111111101110110000101111;
    rom[11620] = 25'b1111111101110110110011111;
    rom[11621] = 25'b1111111101110111100010000;
    rom[11622] = 25'b1111111101111000010000010;
    rom[11623] = 25'b1111111101111000111110100;
    rom[11624] = 25'b1111111101111001101101000;
    rom[11625] = 25'b1111111101111010011011101;
    rom[11626] = 25'b1111111101111011001010010;
    rom[11627] = 25'b1111111101111011111001000;
    rom[11628] = 25'b1111111101111100100111110;
    rom[11629] = 25'b1111111101111101010110110;
    rom[11630] = 25'b1111111101111110000101111;
    rom[11631] = 25'b1111111101111110110101001;
    rom[11632] = 25'b1111111101111111100100011;
    rom[11633] = 25'b1111111110000000010011111;
    rom[11634] = 25'b1111111110000001000011010;
    rom[11635] = 25'b1111111110000001110010110;
    rom[11636] = 25'b1111111110000010100010100;
    rom[11637] = 25'b1111111110000011010010010;
    rom[11638] = 25'b1111111110000100000010001;
    rom[11639] = 25'b1111111110000100110010000;
    rom[11640] = 25'b1111111110000101100010000;
    rom[11641] = 25'b1111111110000110010010000;
    rom[11642] = 25'b1111111110000111000010001;
    rom[11643] = 25'b1111111110000111110010100;
    rom[11644] = 25'b1111111110001000100010110;
    rom[11645] = 25'b1111111110001001010011001;
    rom[11646] = 25'b1111111110001010000011101;
    rom[11647] = 25'b1111111110001010110100001;
    rom[11648] = 25'b1111111110001011100100111;
    rom[11649] = 25'b1111111110001100010101100;
    rom[11650] = 25'b1111111110001101000110010;
    rom[11651] = 25'b1111111110001101110111000;
    rom[11652] = 25'b1111111110001110100111111;
    rom[11653] = 25'b1111111110001111011000111;
    rom[11654] = 25'b1111111110010000001001111;
    rom[11655] = 25'b1111111110010000111011000;
    rom[11656] = 25'b1111111110010001101100000;
    rom[11657] = 25'b1111111110010010011101001;
    rom[11658] = 25'b1111111110010011001110011;
    rom[11659] = 25'b1111111110010011111111101;
    rom[11660] = 25'b1111111110010100110001000;
    rom[11661] = 25'b1111111110010101100010011;
    rom[11662] = 25'b1111111110010110010011111;
    rom[11663] = 25'b1111111110010111000101010;
    rom[11664] = 25'b1111111110010111110110110;
    rom[11665] = 25'b1111111110011000101000010;
    rom[11666] = 25'b1111111110011001011001111;
    rom[11667] = 25'b1111111110011010001011100;
    rom[11668] = 25'b1111111110011010111101001;
    rom[11669] = 25'b1111111110011011101110111;
    rom[11670] = 25'b1111111110011100100000101;
    rom[11671] = 25'b1111111110011101010010011;
    rom[11672] = 25'b1111111110011110000100001;
    rom[11673] = 25'b1111111110011110110110000;
    rom[11674] = 25'b1111111110011111100111110;
    rom[11675] = 25'b1111111110100000011001101;
    rom[11676] = 25'b1111111110100001001011100;
    rom[11677] = 25'b1111111110100001111101100;
    rom[11678] = 25'b1111111110100010101111100;
    rom[11679] = 25'b1111111110100011100001011;
    rom[11680] = 25'b1111111110100100010011011;
    rom[11681] = 25'b1111111110100101000101011;
    rom[11682] = 25'b1111111110100101110111011;
    rom[11683] = 25'b1111111110100110101001011;
    rom[11684] = 25'b1111111110100111011011011;
    rom[11685] = 25'b1111111110101000001101100;
    rom[11686] = 25'b1111111110101000111111100;
    rom[11687] = 25'b1111111110101001110001100;
    rom[11688] = 25'b1111111110101010100011100;
    rom[11689] = 25'b1111111110101011010101101;
    rom[11690] = 25'b1111111110101100000111110;
    rom[11691] = 25'b1111111110101100111001110;
    rom[11692] = 25'b1111111110101101101011111;
    rom[11693] = 25'b1111111110101110011101111;
    rom[11694] = 25'b1111111110101111001111111;
    rom[11695] = 25'b1111111110110000000010000;
    rom[11696] = 25'b1111111110110000110100000;
    rom[11697] = 25'b1111111110110001100110000;
    rom[11698] = 25'b1111111110110010011000001;
    rom[11699] = 25'b1111111110110011001010000;
    rom[11700] = 25'b1111111110110011111100001;
    rom[11701] = 25'b1111111110110100101110001;
    rom[11702] = 25'b1111111110110101100000000;
    rom[11703] = 25'b1111111110110110010010000;
    rom[11704] = 25'b1111111110110111000011111;
    rom[11705] = 25'b1111111110110111110101111;
    rom[11706] = 25'b1111111110111000100111110;
    rom[11707] = 25'b1111111110111001011001100;
    rom[11708] = 25'b1111111110111010001011011;
    rom[11709] = 25'b1111111110111010111101001;
    rom[11710] = 25'b1111111110111011101110111;
    rom[11711] = 25'b1111111110111100100000101;
    rom[11712] = 25'b1111111110111101010010011;
    rom[11713] = 25'b1111111110111110000100001;
    rom[11714] = 25'b1111111110111110110101110;
    rom[11715] = 25'b1111111110111111100111011;
    rom[11716] = 25'b1111111111000000011001000;
    rom[11717] = 25'b1111111111000001001010101;
    rom[11718] = 25'b1111111111000001111100000;
    rom[11719] = 25'b1111111111000010101101100;
    rom[11720] = 25'b1111111111000011011110111;
    rom[11721] = 25'b1111111111000100010000010;
    rom[11722] = 25'b1111111111000101000001101;
    rom[11723] = 25'b1111111111000101110011000;
    rom[11724] = 25'b1111111111000110100100010;
    rom[11725] = 25'b1111111111000111010101010;
    rom[11726] = 25'b1111111111001000000110100;
    rom[11727] = 25'b1111111111001000110111100;
    rom[11728] = 25'b1111111111001001101000101;
    rom[11729] = 25'b1111111111001010011001100;
    rom[11730] = 25'b1111111111001011001010101;
    rom[11731] = 25'b1111111111001011111011011;
    rom[11732] = 25'b1111111111001100101100001;
    rom[11733] = 25'b1111111111001101011101000;
    rom[11734] = 25'b1111111111001110001101101;
    rom[11735] = 25'b1111111111001110111110010;
    rom[11736] = 25'b1111111111001111101110111;
    rom[11737] = 25'b1111111111010000011111010;
    rom[11738] = 25'b1111111111010001001111110;
    rom[11739] = 25'b1111111111010010000000001;
    rom[11740] = 25'b1111111111010010110000011;
    rom[11741] = 25'b1111111111010011100000101;
    rom[11742] = 25'b1111111111010100010000111;
    rom[11743] = 25'b1111111111010101000000111;
    rom[11744] = 25'b1111111111010101110001000;
    rom[11745] = 25'b1111111111010110100000111;
    rom[11746] = 25'b1111111111010111010000110;
    rom[11747] = 25'b1111111111011000000000100;
    rom[11748] = 25'b1111111111011000110000010;
    rom[11749] = 25'b1111111111011001011111111;
    rom[11750] = 25'b1111111111011010001111011;
    rom[11751] = 25'b1111111111011010111110111;
    rom[11752] = 25'b1111111111011011101110001;
    rom[11753] = 25'b1111111111011100011101100;
    rom[11754] = 25'b1111111111011101001100110;
    rom[11755] = 25'b1111111111011101111011111;
    rom[11756] = 25'b1111111111011110101010111;
    rom[11757] = 25'b1111111111011111011001111;
    rom[11758] = 25'b1111111111100000001000101;
    rom[11759] = 25'b1111111111100000110111011;
    rom[11760] = 25'b1111111111100001100110001;
    rom[11761] = 25'b1111111111100010010100101;
    rom[11762] = 25'b1111111111100011000011010;
    rom[11763] = 25'b1111111111100011110001101;
    rom[11764] = 25'b1111111111100100011111111;
    rom[11765] = 25'b1111111111100101001110001;
    rom[11766] = 25'b1111111111100101111100001;
    rom[11767] = 25'b1111111111100110101010001;
    rom[11768] = 25'b1111111111100111011000001;
    rom[11769] = 25'b1111111111101000000101110;
    rom[11770] = 25'b1111111111101000110011100;
    rom[11771] = 25'b1111111111101001100001001;
    rom[11772] = 25'b1111111111101010001110101;
    rom[11773] = 25'b1111111111101010111011111;
    rom[11774] = 25'b1111111111101011101001001;
    rom[11775] = 25'b1111111111101100010110011;
    rom[11776] = 25'b1111111111101101000011011;
    rom[11777] = 25'b1111111111101101110000010;
    rom[11778] = 25'b1111111111101110011101001;
    rom[11779] = 25'b1111111111101111001001111;
    rom[11780] = 25'b1111111111101111110110100;
    rom[11781] = 25'b1111111111110000100010111;
    rom[11782] = 25'b1111111111110001001111010;
    rom[11783] = 25'b1111111111110001111011100;
    rom[11784] = 25'b1111111111110010100111110;
    rom[11785] = 25'b1111111111110011010011101;
    rom[11786] = 25'b1111111111110011111111100;
    rom[11787] = 25'b1111111111110100101011011;
    rom[11788] = 25'b1111111111110101010111000;
    rom[11789] = 25'b1111111111110110000010100;
    rom[11790] = 25'b1111111111110110101101111;
    rom[11791] = 25'b1111111111110111011001001;
    rom[11792] = 25'b1111111111111000000100010;
    rom[11793] = 25'b1111111111111000101111011;
    rom[11794] = 25'b1111111111111001011010010;
    rom[11795] = 25'b1111111111111010000101000;
    rom[11796] = 25'b1111111111111010101111101;
    rom[11797] = 25'b1111111111111011011010001;
    rom[11798] = 25'b1111111111111100000100100;
    rom[11799] = 25'b1111111111111100101110110;
    rom[11800] = 25'b1111111111111101011000111;
    rom[11801] = 25'b1111111111111110000010110;
    rom[11802] = 25'b1111111111111110101100110;
    rom[11803] = 25'b1111111111111111010110011;
    rom[11804] = 25'b0000000000000000000000000;
    rom[11805] = 25'b0000000000000000101001010;
    rom[11806] = 25'b0000000000000001010010101;
    rom[11807] = 25'b0000000000000001111011110;
    rom[11808] = 25'b0000000000000010100100111;
    rom[11809] = 25'b0000000000000011001101101;
    rom[11810] = 25'b0000000000000011110110100;
    rom[11811] = 25'b0000000000000100011111000;
    rom[11812] = 25'b0000000000000101000111100;
    rom[11813] = 25'b0000000000000101101111110;
    rom[11814] = 25'b0000000000000110011000000;
    rom[11815] = 25'b0000000000000111000000000;
    rom[11816] = 25'b0000000000000111100111111;
    rom[11817] = 25'b0000000000001000001111101;
    rom[11818] = 25'b0000000000001000110111010;
    rom[11819] = 25'b0000000000001001011110101;
    rom[11820] = 25'b0000000000001010000101111;
    rom[11821] = 25'b0000000000001010101101001;
    rom[11822] = 25'b0000000000001011010100000;
    rom[11823] = 25'b0000000000001011111011000;
    rom[11824] = 25'b0000000000001100100001101;
    rom[11825] = 25'b0000000000001101001000001;
    rom[11826] = 25'b0000000000001101101110100;
    rom[11827] = 25'b0000000000001110010100110;
    rom[11828] = 25'b0000000000001110111010111;
    rom[11829] = 25'b0000000000001111100000110;
    rom[11830] = 25'b0000000000010000000110100;
    rom[11831] = 25'b0000000000010000101100001;
    rom[11832] = 25'b0000000000010001010001101;
    rom[11833] = 25'b0000000000010001110110111;
    rom[11834] = 25'b0000000000010010011100000;
    rom[11835] = 25'b0000000000010011000001000;
    rom[11836] = 25'b0000000000010011100101110;
    rom[11837] = 25'b0000000000010100001010100;
    rom[11838] = 25'b0000000000010100101111000;
    rom[11839] = 25'b0000000000010101010011010;
    rom[11840] = 25'b0000000000010101110111100;
    rom[11841] = 25'b0000000000010110011011100;
    rom[11842] = 25'b0000000000010110111111011;
    rom[11843] = 25'b0000000000010111100011000;
    rom[11844] = 25'b0000000000011000000110101;
    rom[11845] = 25'b0000000000011000101001111;
    rom[11846] = 25'b0000000000011001001101001;
    rom[11847] = 25'b0000000000011001110000010;
    rom[11848] = 25'b0000000000011010010011001;
    rom[11849] = 25'b0000000000011010110101110;
    rom[11850] = 25'b0000000000011011011000010;
    rom[11851] = 25'b0000000000011011111010101;
    rom[11852] = 25'b0000000000011100011100111;
    rom[11853] = 25'b0000000000011100111110111;
    rom[11854] = 25'b0000000000011101100000101;
    rom[11855] = 25'b0000000000011110000010011;
    rom[11856] = 25'b0000000000011110100100000;
    rom[11857] = 25'b0000000000011111000101010;
    rom[11858] = 25'b0000000000011111100110011;
    rom[11859] = 25'b0000000000100000000111100;
    rom[11860] = 25'b0000000000100000101000011;
    rom[11861] = 25'b0000000000100001001001000;
    rom[11862] = 25'b0000000000100001101001100;
    rom[11863] = 25'b0000000000100010001001111;
    rom[11864] = 25'b0000000000100010101001111;
    rom[11865] = 25'b0000000000100011001001111;
    rom[11866] = 25'b0000000000100011101001110;
    rom[11867] = 25'b0000000000100100001001010;
    rom[11868] = 25'b0000000000100100101000110;
    rom[11869] = 25'b0000000000100101001000000;
    rom[11870] = 25'b0000000000100101100111000;
    rom[11871] = 25'b0000000000100110000110000;
    rom[11872] = 25'b0000000000100110100100110;
    rom[11873] = 25'b0000000000100111000011011;
    rom[11874] = 25'b0000000000100111100001110;
    rom[11875] = 25'b0000000000100111111111111;
    rom[11876] = 25'b0000000000101000011101111;
    rom[11877] = 25'b0000000000101000111011110;
    rom[11878] = 25'b0000000000101001011001100;
    rom[11879] = 25'b0000000000101001110110111;
    rom[11880] = 25'b0000000000101010010100010;
    rom[11881] = 25'b0000000000101010110001011;
    rom[11882] = 25'b0000000000101011001110010;
    rom[11883] = 25'b0000000000101011101011001;
    rom[11884] = 25'b0000000000101100000111110;
    rom[11885] = 25'b0000000000101100100100001;
    rom[11886] = 25'b0000000000101101000000011;
    rom[11887] = 25'b0000000000101101011100011;
    rom[11888] = 25'b0000000000101101111000010;
    rom[11889] = 25'b0000000000101110010011111;
    rom[11890] = 25'b0000000000101110101111100;
    rom[11891] = 25'b0000000000101111001010110;
    rom[11892] = 25'b0000000000101111100101111;
    rom[11893] = 25'b0000000000110000000000111;
    rom[11894] = 25'b0000000000110000011011101;
    rom[11895] = 25'b0000000000110000110110001;
    rom[11896] = 25'b0000000000110001010000101;
    rom[11897] = 25'b0000000000110001101010110;
    rom[11898] = 25'b0000000000110010000100111;
    rom[11899] = 25'b0000000000110010011110101;
    rom[11900] = 25'b0000000000110010111000011;
    rom[11901] = 25'b0000000000110011010001110;
    rom[11902] = 25'b0000000000110011101011001;
    rom[11903] = 25'b0000000000110100000100010;
    rom[11904] = 25'b0000000000110100011101001;
    rom[11905] = 25'b0000000000110100110110000;
    rom[11906] = 25'b0000000000110101001110100;
    rom[11907] = 25'b0000000000110101100110111;
    rom[11908] = 25'b0000000000110101111111000;
    rom[11909] = 25'b0000000000110110010111000;
    rom[11910] = 25'b0000000000110110101110111;
    rom[11911] = 25'b0000000000110111000110011;
    rom[11912] = 25'b0000000000110111011101111;
    rom[11913] = 25'b0000000000110111110101010;
    rom[11914] = 25'b0000000000111000001100010;
    rom[11915] = 25'b0000000000111000100011001;
    rom[11916] = 25'b0000000000111000111001110;
    rom[11917] = 25'b0000000000111001010000010;
    rom[11918] = 25'b0000000000111001100110101;
    rom[11919] = 25'b0000000000111001111100110;
    rom[11920] = 25'b0000000000111010010010110;
    rom[11921] = 25'b0000000000111010101000100;
    rom[11922] = 25'b0000000000111010111110000;
    rom[11923] = 25'b0000000000111011010011011;
    rom[11924] = 25'b0000000000111011101000101;
    rom[11925] = 25'b0000000000111011111101101;
    rom[11926] = 25'b0000000000111100010010011;
    rom[11927] = 25'b0000000000111100100111000;
    rom[11928] = 25'b0000000000111100111011101;
    rom[11929] = 25'b0000000000111101001111110;
    rom[11930] = 25'b0000000000111101100011111;
    rom[11931] = 25'b0000000000111101110111110;
    rom[11932] = 25'b0000000000111110001011100;
    rom[11933] = 25'b0000000000111110011111000;
    rom[11934] = 25'b0000000000111110110010011;
    rom[11935] = 25'b0000000000111111000101100;
    rom[11936] = 25'b0000000000111111011000011;
    rom[11937] = 25'b0000000000111111101011010;
    rom[11938] = 25'b0000000000111111111101110;
    rom[11939] = 25'b0000000001000000010000010;
    rom[11940] = 25'b0000000001000000100010011;
    rom[11941] = 25'b0000000001000000110100011;
    rom[11942] = 25'b0000000001000001000110010;
    rom[11943] = 25'b0000000001000001010111111;
    rom[11944] = 25'b0000000001000001101001010;
    rom[11945] = 25'b0000000001000001111010101;
    rom[11946] = 25'b0000000001000010001011110;
    rom[11947] = 25'b0000000001000010011100101;
    rom[11948] = 25'b0000000001000010101101011;
    rom[11949] = 25'b0000000001000010111101110;
    rom[11950] = 25'b0000000001000011001110001;
    rom[11951] = 25'b0000000001000011011110011;
    rom[11952] = 25'b0000000001000011101110010;
    rom[11953] = 25'b0000000001000011111110001;
    rom[11954] = 25'b0000000001000100001101101;
    rom[11955] = 25'b0000000001000100011101001;
    rom[11956] = 25'b0000000001000100101100011;
    rom[11957] = 25'b0000000001000100111011011;
    rom[11958] = 25'b0000000001000101001010010;
    rom[11959] = 25'b0000000001000101011000111;
    rom[11960] = 25'b0000000001000101100111011;
    rom[11961] = 25'b0000000001000101110101110;
    rom[11962] = 25'b0000000001000110000011111;
    rom[11963] = 25'b0000000001000110010001110;
    rom[11964] = 25'b0000000001000110011111100;
    rom[11965] = 25'b0000000001000110101101001;
    rom[11966] = 25'b0000000001000110111010100;
    rom[11967] = 25'b0000000001000111000111110;
    rom[11968] = 25'b0000000001000111010100101;
    rom[11969] = 25'b0000000001000111100001100;
    rom[11970] = 25'b0000000001000111101110001;
    rom[11971] = 25'b0000000001000111111010101;
    rom[11972] = 25'b0000000001001000000111000;
    rom[11973] = 25'b0000000001001000010011001;
    rom[11974] = 25'b0000000001001000011111000;
    rom[11975] = 25'b0000000001001000101010110;
    rom[11976] = 25'b0000000001001000110110010;
    rom[11977] = 25'b0000000001001001000001101;
    rom[11978] = 25'b0000000001001001001100111;
    rom[11979] = 25'b0000000001001001011000000;
    rom[11980] = 25'b0000000001001001100010110;
    rom[11981] = 25'b0000000001001001101101100;
    rom[11982] = 25'b0000000001001001110111111;
    rom[11983] = 25'b0000000001001010000010001;
    rom[11984] = 25'b0000000001001010001100011;
    rom[11985] = 25'b0000000001001010010110010;
    rom[11986] = 25'b0000000001001010100000000;
    rom[11987] = 25'b0000000001001010101001101;
    rom[11988] = 25'b0000000001001010110011001;
    rom[11989] = 25'b0000000001001010111100011;
    rom[11990] = 25'b0000000001001011000101011;
    rom[11991] = 25'b0000000001001011001110001;
    rom[11992] = 25'b0000000001001011010110111;
    rom[11993] = 25'b0000000001001011011111011;
    rom[11994] = 25'b0000000001001011100111110;
    rom[11995] = 25'b0000000001001011110000000;
    rom[11996] = 25'b0000000001001011111000000;
    rom[11997] = 25'b0000000001001011111111111;
    rom[11998] = 25'b0000000001001100000111100;
    rom[11999] = 25'b0000000001001100001110111;
    rom[12000] = 25'b0000000001001100010110010;
    rom[12001] = 25'b0000000001001100011101011;
    rom[12002] = 25'b0000000001001100100100010;
    rom[12003] = 25'b0000000001001100101011001;
    rom[12004] = 25'b0000000001001100110001110;
    rom[12005] = 25'b0000000001001100111000001;
    rom[12006] = 25'b0000000001001100111110100;
    rom[12007] = 25'b0000000001001101000100100;
    rom[12008] = 25'b0000000001001101001010100;
    rom[12009] = 25'b0000000001001101010000010;
    rom[12010] = 25'b0000000001001101010101110;
    rom[12011] = 25'b0000000001001101011011001;
    rom[12012] = 25'b0000000001001101100000100;
    rom[12013] = 25'b0000000001001101100101100;
    rom[12014] = 25'b0000000001001101101010100;
    rom[12015] = 25'b0000000001001101101111001;
    rom[12016] = 25'b0000000001001101110011110;
    rom[12017] = 25'b0000000001001101111000001;
    rom[12018] = 25'b0000000001001101111100011;
    rom[12019] = 25'b0000000001001110000000100;
    rom[12020] = 25'b0000000001001110000100011;
    rom[12021] = 25'b0000000001001110001000001;
    rom[12022] = 25'b0000000001001110001011101;
    rom[12023] = 25'b0000000001001110001111000;
    rom[12024] = 25'b0000000001001110010010011;
    rom[12025] = 25'b0000000001001110010101011;
    rom[12026] = 25'b0000000001001110011000010;
    rom[12027] = 25'b0000000001001110011011000;
    rom[12028] = 25'b0000000001001110011101110;
    rom[12029] = 25'b0000000001001110100000001;
    rom[12030] = 25'b0000000001001110100010011;
    rom[12031] = 25'b0000000001001110100100100;
    rom[12032] = 25'b0000000001001110100110011;
    rom[12033] = 25'b0000000001001110101000010;
    rom[12034] = 25'b0000000001001110101001111;
    rom[12035] = 25'b0000000001001110101011010;
    rom[12036] = 25'b0000000001001110101100110;
    rom[12037] = 25'b0000000001001110101101111;
    rom[12038] = 25'b0000000001001110101110111;
    rom[12039] = 25'b0000000001001110101111101;
    rom[12040] = 25'b0000000001001110110000010;
    rom[12041] = 25'b0000000001001110110000111;
    rom[12042] = 25'b0000000001001110110001010;
    rom[12043] = 25'b0000000001001110110001100;
    rom[12044] = 25'b0000000001001110110001101;
    rom[12045] = 25'b0000000001001110110001100;
    rom[12046] = 25'b0000000001001110110001010;
    rom[12047] = 25'b0000000001001110110000111;
    rom[12048] = 25'b0000000001001110110000010;
    rom[12049] = 25'b0000000001001110101111101;
    rom[12050] = 25'b0000000001001110101110110;
    rom[12051] = 25'b0000000001001110101101110;
    rom[12052] = 25'b0000000001001110101100101;
    rom[12053] = 25'b0000000001001110101011010;
    rom[12054] = 25'b0000000001001110101001111;
    rom[12055] = 25'b0000000001001110101000010;
    rom[12056] = 25'b0000000001001110100110100;
    rom[12057] = 25'b0000000001001110100100101;
    rom[12058] = 25'b0000000001001110100010101;
    rom[12059] = 25'b0000000001001110100000011;
    rom[12060] = 25'b0000000001001110011110000;
    rom[12061] = 25'b0000000001001110011011101;
    rom[12062] = 25'b0000000001001110011000111;
    rom[12063] = 25'b0000000001001110010110001;
    rom[12064] = 25'b0000000001001110010011010;
    rom[12065] = 25'b0000000001001110010000010;
    rom[12066] = 25'b0000000001001110001101000;
    rom[12067] = 25'b0000000001001110001001110;
    rom[12068] = 25'b0000000001001110000110010;
    rom[12069] = 25'b0000000001001110000010101;
    rom[12070] = 25'b0000000001001101111110111;
    rom[12071] = 25'b0000000001001101111011000;
    rom[12072] = 25'b0000000001001101110111000;
    rom[12073] = 25'b0000000001001101110010110;
    rom[12074] = 25'b0000000001001101101110100;
    rom[12075] = 25'b0000000001001101101010000;
    rom[12076] = 25'b0000000001001101100101100;
    rom[12077] = 25'b0000000001001101100000110;
    rom[12078] = 25'b0000000001001101011011111;
    rom[12079] = 25'b0000000001001101010110111;
    rom[12080] = 25'b0000000001001101010001110;
    rom[12081] = 25'b0000000001001101001100100;
    rom[12082] = 25'b0000000001001101000111001;
    rom[12083] = 25'b0000000001001101000001101;
    rom[12084] = 25'b0000000001001100111100000;
    rom[12085] = 25'b0000000001001100110110001;
    rom[12086] = 25'b0000000001001100110000010;
    rom[12087] = 25'b0000000001001100101010010;
    rom[12088] = 25'b0000000001001100100100001;
    rom[12089] = 25'b0000000001001100011101110;
    rom[12090] = 25'b0000000001001100010111011;
    rom[12091] = 25'b0000000001001100010000111;
    rom[12092] = 25'b0000000001001100001010001;
    rom[12093] = 25'b0000000001001100000011011;
    rom[12094] = 25'b0000000001001011111100011;
    rom[12095] = 25'b0000000001001011110101011;
    rom[12096] = 25'b0000000001001011101110001;
    rom[12097] = 25'b0000000001001011100111000;
    rom[12098] = 25'b0000000001001011011111100;
    rom[12099] = 25'b0000000001001011011000000;
    rom[12100] = 25'b0000000001001011010000010;
    rom[12101] = 25'b0000000001001011001000100;
    rom[12102] = 25'b0000000001001011000000101;
    rom[12103] = 25'b0000000001001010111000101;
    rom[12104] = 25'b0000000001001010110000011;
    rom[12105] = 25'b0000000001001010101000010;
    rom[12106] = 25'b0000000001001010011111111;
    rom[12107] = 25'b0000000001001010010111011;
    rom[12108] = 25'b0000000001001010001110110;
    rom[12109] = 25'b0000000001001010000110000;
    rom[12110] = 25'b0000000001001001111101001;
    rom[12111] = 25'b0000000001001001110100010;
    rom[12112] = 25'b0000000001001001101011010;
    rom[12113] = 25'b0000000001001001100010000;
    rom[12114] = 25'b0000000001001001011000110;
    rom[12115] = 25'b0000000001001001001111010;
    rom[12116] = 25'b0000000001001001000101110;
    rom[12117] = 25'b0000000001001000111100010;
    rom[12118] = 25'b0000000001001000110010011;
    rom[12119] = 25'b0000000001001000101000101;
    rom[12120] = 25'b0000000001001000011110101;
    rom[12121] = 25'b0000000001001000010100100;
    rom[12122] = 25'b0000000001001000001010100;
    rom[12123] = 25'b0000000001001000000000001;
    rom[12124] = 25'b0000000001000111110101111;
    rom[12125] = 25'b0000000001000111101011010;
    rom[12126] = 25'b0000000001000111100000110;
    rom[12127] = 25'b0000000001000111010110000;
    rom[12128] = 25'b0000000001000111001011010;
    rom[12129] = 25'b0000000001000111000000100;
    rom[12130] = 25'b0000000001000110110101011;
    rom[12131] = 25'b0000000001000110101010011;
    rom[12132] = 25'b0000000001000110011111010;
    rom[12133] = 25'b0000000001000110010011111;
    rom[12134] = 25'b0000000001000110001000100;
    rom[12135] = 25'b0000000001000101111101001;
    rom[12136] = 25'b0000000001000101110001100;
    rom[12137] = 25'b0000000001000101100101110;
    rom[12138] = 25'b0000000001000101011010001;
    rom[12139] = 25'b0000000001000101001110001;
    rom[12140] = 25'b0000000001000101000010010;
    rom[12141] = 25'b0000000001000100110110001;
    rom[12142] = 25'b0000000001000100101010000;
    rom[12143] = 25'b0000000001000100011101110;
    rom[12144] = 25'b0000000001000100010001100;
    rom[12145] = 25'b0000000001000100000101000;
    rom[12146] = 25'b0000000001000011111000101;
    rom[12147] = 25'b0000000001000011101100000;
    rom[12148] = 25'b0000000001000011011111010;
    rom[12149] = 25'b0000000001000011010010100;
    rom[12150] = 25'b0000000001000011000101101;
    rom[12151] = 25'b0000000001000010111000110;
    rom[12152] = 25'b0000000001000010101011110;
    rom[12153] = 25'b0000000001000010011110101;
    rom[12154] = 25'b0000000001000010010001011;
    rom[12155] = 25'b0000000001000010000100010;
    rom[12156] = 25'b0000000001000001110110110;
    rom[12157] = 25'b0000000001000001101001010;
    rom[12158] = 25'b0000000001000001011011110;
    rom[12159] = 25'b0000000001000001001110001;
    rom[12160] = 25'b0000000001000001000000101;
    rom[12161] = 25'b0000000001000000110010110;
    rom[12162] = 25'b0000000001000000100100111;
    rom[12163] = 25'b0000000001000000010111000;
    rom[12164] = 25'b0000000001000000001001000;
    rom[12165] = 25'b0000000000111111111011000;
    rom[12166] = 25'b0000000000111111101100110;
    rom[12167] = 25'b0000000000111111011110100;
    rom[12168] = 25'b0000000000111111010000010;
    rom[12169] = 25'b0000000000111111000001111;
    rom[12170] = 25'b0000000000111110110011011;
    rom[12171] = 25'b0000000000111110100100111;
    rom[12172] = 25'b0000000000111110010110011;
    rom[12173] = 25'b0000000000111110000111110;
    rom[12174] = 25'b0000000000111101111000111;
    rom[12175] = 25'b0000000000111101101010001;
    rom[12176] = 25'b0000000000111101011011010;
    rom[12177] = 25'b0000000000111101001100011;
    rom[12178] = 25'b0000000000111100111101010;
    rom[12179] = 25'b0000000000111100101110010;
    rom[12180] = 25'b0000000000111100011111001;
    rom[12181] = 25'b0000000000111100001111111;
    rom[12182] = 25'b0000000000111100000000101;
    rom[12183] = 25'b0000000000111011110001011;
    rom[12184] = 25'b0000000000111011100010000;
    rom[12185] = 25'b0000000000111011010010011;
    rom[12186] = 25'b0000000000111011000010111;
    rom[12187] = 25'b0000000000111010110011011;
    rom[12188] = 25'b0000000000111010100011110;
    rom[12189] = 25'b0000000000111010010100000;
    rom[12190] = 25'b0000000000111010000100010;
    rom[12191] = 25'b0000000000111001110100100;
    rom[12192] = 25'b0000000000111001100100101;
    rom[12193] = 25'b0000000000111001010100101;
    rom[12194] = 25'b0000000000111001000100110;
    rom[12195] = 25'b0000000000111000110100101;
    rom[12196] = 25'b0000000000111000100100100;
    rom[12197] = 25'b0000000000111000010100100;
    rom[12198] = 25'b0000000000111000000100010;
    rom[12199] = 25'b0000000000110111110011111;
    rom[12200] = 25'b0000000000110111100011101;
    rom[12201] = 25'b0000000000110111010011010;
    rom[12202] = 25'b0000000000110111000010111;
    rom[12203] = 25'b0000000000110110110010011;
    rom[12204] = 25'b0000000000110110100010000;
    rom[12205] = 25'b0000000000110110010001011;
    rom[12206] = 25'b0000000000110110000000110;
    rom[12207] = 25'b0000000000110101110000001;
    rom[12208] = 25'b0000000000110101011111011;
    rom[12209] = 25'b0000000000110101001110101;
    rom[12210] = 25'b0000000000110100111101111;
    rom[12211] = 25'b0000000000110100101101000;
    rom[12212] = 25'b0000000000110100011100001;
    rom[12213] = 25'b0000000000110100001011010;
    rom[12214] = 25'b0000000000110011111010010;
    rom[12215] = 25'b0000000000110011101001010;
    rom[12216] = 25'b0000000000110011011000001;
    rom[12217] = 25'b0000000000110011000111001;
    rom[12218] = 25'b0000000000110010110110000;
    rom[12219] = 25'b0000000000110010100100111;
    rom[12220] = 25'b0000000000110010010011101;
    rom[12221] = 25'b0000000000110010000010011;
    rom[12222] = 25'b0000000000110001110001001;
    rom[12223] = 25'b0000000000110001011111111;
    rom[12224] = 25'b0000000000110001001110100;
    rom[12225] = 25'b0000000000110000111101001;
    rom[12226] = 25'b0000000000110000101011101;
    rom[12227] = 25'b0000000000110000011010010;
    rom[12228] = 25'b0000000000110000001000110;
    rom[12229] = 25'b0000000000101111110111010;
    rom[12230] = 25'b0000000000101111100101101;
    rom[12231] = 25'b0000000000101111010100001;
    rom[12232] = 25'b0000000000101111000010100;
    rom[12233] = 25'b0000000000101110110000111;
    rom[12234] = 25'b0000000000101110011111010;
    rom[12235] = 25'b0000000000101110001101100;
    rom[12236] = 25'b0000000000101101111011110;
    rom[12237] = 25'b0000000000101101101010000;
    rom[12238] = 25'b0000000000101101011000001;
    rom[12239] = 25'b0000000000101101000110011;
    rom[12240] = 25'b0000000000101100110100100;
    rom[12241] = 25'b0000000000101100100010110;
    rom[12242] = 25'b0000000000101100010000111;
    rom[12243] = 25'b0000000000101011111111000;
    rom[12244] = 25'b0000000000101011101101000;
    rom[12245] = 25'b0000000000101011011011000;
    rom[12246] = 25'b0000000000101011001001001;
    rom[12247] = 25'b0000000000101010110111001;
    rom[12248] = 25'b0000000000101010100101001;
    rom[12249] = 25'b0000000000101010010011001;
    rom[12250] = 25'b0000000000101010000001000;
    rom[12251] = 25'b0000000000101001101110111;
    rom[12252] = 25'b0000000000101001011100111;
    rom[12253] = 25'b0000000000101001001010110;
    rom[12254] = 25'b0000000000101000111000110;
    rom[12255] = 25'b0000000000101000100110100;
    rom[12256] = 25'b0000000000101000010100011;
    rom[12257] = 25'b0000000000101000000010010;
    rom[12258] = 25'b0000000000100111110000001;
    rom[12259] = 25'b0000000000100111011101111;
    rom[12260] = 25'b0000000000100111001011101;
    rom[12261] = 25'b0000000000100110111001100;
    rom[12262] = 25'b0000000000100110100111010;
    rom[12263] = 25'b0000000000100110010101000;
    rom[12264] = 25'b0000000000100110000010110;
    rom[12265] = 25'b0000000000100101110000100;
    rom[12266] = 25'b0000000000100101011110010;
    rom[12267] = 25'b0000000000100101001100000;
    rom[12268] = 25'b0000000000100100111001101;
    rom[12269] = 25'b0000000000100100100111011;
    rom[12270] = 25'b0000000000100100010101001;
    rom[12271] = 25'b0000000000100100000010110;
    rom[12272] = 25'b0000000000100011110000100;
    rom[12273] = 25'b0000000000100011011110010;
    rom[12274] = 25'b0000000000100011001100000;
    rom[12275] = 25'b0000000000100010111001100;
    rom[12276] = 25'b0000000000100010100111010;
    rom[12277] = 25'b0000000000100010010101000;
    rom[12278] = 25'b0000000000100010000010101;
    rom[12279] = 25'b0000000000100001110000010;
    rom[12280] = 25'b0000000000100001011110000;
    rom[12281] = 25'b0000000000100001001011101;
    rom[12282] = 25'b0000000000100000111001011;
    rom[12283] = 25'b0000000000100000100111000;
    rom[12284] = 25'b0000000000100000010100101;
    rom[12285] = 25'b0000000000100000000010011;
    rom[12286] = 25'b0000000000011111110000000;
    rom[12287] = 25'b0000000000011111011101110;
    rom[12288] = 25'b0000000000011111001011011;
    rom[12289] = 25'b0000000000011110111001001;
    rom[12290] = 25'b0000000000011110100110111;
    rom[12291] = 25'b0000000000011110010100100;
    rom[12292] = 25'b0000000000011110000010010;
    rom[12293] = 25'b0000000000011101110000000;
    rom[12294] = 25'b0000000000011101011101110;
    rom[12295] = 25'b0000000000011101001011011;
    rom[12296] = 25'b0000000000011100111001001;
    rom[12297] = 25'b0000000000011100100110111;
    rom[12298] = 25'b0000000000011100010100101;
    rom[12299] = 25'b0000000000011100000010011;
    rom[12300] = 25'b0000000000011011110000010;
    rom[12301] = 25'b0000000000011011011110000;
    rom[12302] = 25'b0000000000011011001011111;
    rom[12303] = 25'b0000000000011010111001100;
    rom[12304] = 25'b0000000000011010100111100;
    rom[12305] = 25'b0000000000011010010101010;
    rom[12306] = 25'b0000000000011010000011001;
    rom[12307] = 25'b0000000000011001110001000;
    rom[12308] = 25'b0000000000011001011110111;
    rom[12309] = 25'b0000000000011001001100110;
    rom[12310] = 25'b0000000000011000111010110;
    rom[12311] = 25'b0000000000011000101000101;
    rom[12312] = 25'b0000000000011000010110101;
    rom[12313] = 25'b0000000000011000000100100;
    rom[12314] = 25'b0000000000010111110010100;
    rom[12315] = 25'b0000000000010111100000100;
    rom[12316] = 25'b0000000000010111001110100;
    rom[12317] = 25'b0000000000010110111100100;
    rom[12318] = 25'b0000000000010110101010101;
    rom[12319] = 25'b0000000000010110011000110;
    rom[12320] = 25'b0000000000010110000110110;
    rom[12321] = 25'b0000000000010101110100111;
    rom[12322] = 25'b0000000000010101100011000;
    rom[12323] = 25'b0000000000010101010001001;
    rom[12324] = 25'b0000000000010100111111011;
    rom[12325] = 25'b0000000000010100101101100;
    rom[12326] = 25'b0000000000010100011011110;
    rom[12327] = 25'b0000000000010100001010000;
    rom[12328] = 25'b0000000000010011111000011;
    rom[12329] = 25'b0000000000010011100110101;
    rom[12330] = 25'b0000000000010011010101000;
    rom[12331] = 25'b0000000000010011000011011;
    rom[12332] = 25'b0000000000010010110001110;
    rom[12333] = 25'b0000000000010010100000001;
    rom[12334] = 25'b0000000000010010001110101;
    rom[12335] = 25'b0000000000010001111101001;
    rom[12336] = 25'b0000000000010001101011100;
    rom[12337] = 25'b0000000000010001011010001;
    rom[12338] = 25'b0000000000010001001000101;
    rom[12339] = 25'b0000000000010000110111010;
    rom[12340] = 25'b0000000000010000100101110;
    rom[12341] = 25'b0000000000010000010100100;
    rom[12342] = 25'b0000000000010000000011001;
    rom[12343] = 25'b0000000000001111110001110;
    rom[12344] = 25'b0000000000001111100000101;
    rom[12345] = 25'b0000000000001111001111010;
    rom[12346] = 25'b0000000000001110111110001;
    rom[12347] = 25'b0000000000001110101100111;
    rom[12348] = 25'b0000000000001110011011110;
    rom[12349] = 25'b0000000000001110001010101;
    rom[12350] = 25'b0000000000001101111001101;
    rom[12351] = 25'b0000000000001101101000100;
    rom[12352] = 25'b0000000000001101010111100;
    rom[12353] = 25'b0000000000001101000110101;
    rom[12354] = 25'b0000000000001100110101110;
    rom[12355] = 25'b0000000000001100100100111;
    rom[12356] = 25'b0000000000001100010011111;
    rom[12357] = 25'b0000000000001100000011001;
    rom[12358] = 25'b0000000000001011110010011;
    rom[12359] = 25'b0000000000001011100001101;
    rom[12360] = 25'b0000000000001011010001000;
    rom[12361] = 25'b0000000000001011000000010;
    rom[12362] = 25'b0000000000001010101111101;
    rom[12363] = 25'b0000000000001010011111000;
    rom[12364] = 25'b0000000000001010001110100;
    rom[12365] = 25'b0000000000001001111101111;
    rom[12366] = 25'b0000000000001001101101100;
    rom[12367] = 25'b0000000000001001011101001;
    rom[12368] = 25'b0000000000001001001100110;
    rom[12369] = 25'b0000000000001000111100011;
    rom[12370] = 25'b0000000000001000101100000;
    rom[12371] = 25'b0000000000001000011011110;
    rom[12372] = 25'b0000000000001000001011100;
    rom[12373] = 25'b0000000000000111111011011;
    rom[12374] = 25'b0000000000000111101011010;
    rom[12375] = 25'b0000000000000111011011001;
    rom[12376] = 25'b0000000000000111001011001;
    rom[12377] = 25'b0000000000000110111011001;
    rom[12378] = 25'b0000000000000110101011010;
    rom[12379] = 25'b0000000000000110011011010;
    rom[12380] = 25'b0000000000000110001011011;
    rom[12381] = 25'b0000000000000101111011101;
    rom[12382] = 25'b0000000000000101101011111;
    rom[12383] = 25'b0000000000000101011100001;
    rom[12384] = 25'b0000000000000101001100011;
    rom[12385] = 25'b0000000000000100111100110;
    rom[12386] = 25'b0000000000000100101101001;
    rom[12387] = 25'b0000000000000100011101101;
    rom[12388] = 25'b0000000000000100001110001;
    rom[12389] = 25'b0000000000000011111110101;
    rom[12390] = 25'b0000000000000011101111011;
    rom[12391] = 25'b0000000000000011011111111;
    rom[12392] = 25'b0000000000000011010000101;
    rom[12393] = 25'b0000000000000011000001011;
    rom[12394] = 25'b0000000000000010110010010;
    rom[12395] = 25'b0000000000000010100011001;
    rom[12396] = 25'b0000000000000010010100000;
    rom[12397] = 25'b0000000000000010000100111;
    rom[12398] = 25'b0000000000000001110110000;
    rom[12399] = 25'b0000000000000001100111000;
    rom[12400] = 25'b0000000000000001011000001;
    rom[12401] = 25'b0000000000000001001001010;
    rom[12402] = 25'b0000000000000000111010100;
    rom[12403] = 25'b0000000000000000101011110;
    rom[12404] = 25'b0000000000000000011101001;
    rom[12405] = 25'b0000000000000000001110100;
    rom[12406] = 25'b0000000000000000000000000;
    rom[12407] = 25'b1111111111111111110001100;
    rom[12408] = 25'b1111111111111111100011000;
    rom[12409] = 25'b1111111111111111010100100;
    rom[12410] = 25'b1111111111111111000110010;
    rom[12411] = 25'b1111111111111110111000000;
    rom[12412] = 25'b1111111111111110101001110;
    rom[12413] = 25'b1111111111111110011011100;
    rom[12414] = 25'b1111111111111110001101011;
    rom[12415] = 25'b1111111111111101111111010;
    rom[12416] = 25'b1111111111111101110001010;
    rom[12417] = 25'b1111111111111101100011010;
    rom[12418] = 25'b1111111111111101010101010;
    rom[12419] = 25'b1111111111111101000111100;
    rom[12420] = 25'b1111111111111100111001101;
    rom[12421] = 25'b1111111111111100101100000;
    rom[12422] = 25'b1111111111111100011110010;
    rom[12423] = 25'b1111111111111100010000101;
    rom[12424] = 25'b1111111111111100000011000;
    rom[12425] = 25'b1111111111111011110101100;
    rom[12426] = 25'b1111111111111011101000000;
    rom[12427] = 25'b1111111111111011011010101;
    rom[12428] = 25'b1111111111111011001101011;
    rom[12429] = 25'b1111111111111011000000000;
    rom[12430] = 25'b1111111111111010110010110;
    rom[12431] = 25'b1111111111111010100101101;
    rom[12432] = 25'b1111111111111010011000100;
    rom[12433] = 25'b1111111111111010001011011;
    rom[12434] = 25'b1111111111111001111110100;
    rom[12435] = 25'b1111111111111001110001101;
    rom[12436] = 25'b1111111111111001100100110;
    rom[12437] = 25'b1111111111111001010111111;
    rom[12438] = 25'b1111111111111001001011001;
    rom[12439] = 25'b1111111111111000111110100;
    rom[12440] = 25'b1111111111111000110001110;
    rom[12441] = 25'b1111111111111000100101010;
    rom[12442] = 25'b1111111111111000011000110;
    rom[12443] = 25'b1111111111111000001100010;
    rom[12444] = 25'b1111111111111000000000000;
    rom[12445] = 25'b1111111111110111110011101;
    rom[12446] = 25'b1111111111110111100111011;
    rom[12447] = 25'b1111111111110111011011001;
    rom[12448] = 25'b1111111111110111001111000;
    rom[12449] = 25'b1111111111110111000010111;
    rom[12450] = 25'b1111111111110110110110111;
    rom[12451] = 25'b1111111111110110101011000;
    rom[12452] = 25'b1111111111110110011111001;
    rom[12453] = 25'b1111111111110110010011010;
    rom[12454] = 25'b1111111111110110000111100;
    rom[12455] = 25'b1111111111110101111011110;
    rom[12456] = 25'b1111111111110101110000010;
    rom[12457] = 25'b1111111111110101100100101;
    rom[12458] = 25'b1111111111110101011001001;
    rom[12459] = 25'b1111111111110101001101101;
    rom[12460] = 25'b1111111111110101000010010;
    rom[12461] = 25'b1111111111110100110111000;
    rom[12462] = 25'b1111111111110100101011110;
    rom[12463] = 25'b1111111111110100100000100;
    rom[12464] = 25'b1111111111110100010101011;
    rom[12465] = 25'b1111111111110100001010011;
    rom[12466] = 25'b1111111111110011111111010;
    rom[12467] = 25'b1111111111110011110100100;
    rom[12468] = 25'b1111111111110011101001100;
    rom[12469] = 25'b1111111111110011011110110;
    rom[12470] = 25'b1111111111110011010100000;
    rom[12471] = 25'b1111111111110011001001010;
    rom[12472] = 25'b1111111111110010111110110;
    rom[12473] = 25'b1111111111110010110100010;
    rom[12474] = 25'b1111111111110010101001110;
    rom[12475] = 25'b1111111111110010011111010;
    rom[12476] = 25'b1111111111110010010101000;
    rom[12477] = 25'b1111111111110010001010101;
    rom[12478] = 25'b1111111111110010000000100;
    rom[12479] = 25'b1111111111110001110110011;
    rom[12480] = 25'b1111111111110001101100010;
    rom[12481] = 25'b1111111111110001100010001;
    rom[12482] = 25'b1111111111110001011000010;
    rom[12483] = 25'b1111111111110001001110011;
    rom[12484] = 25'b1111111111110001000100101;
    rom[12485] = 25'b1111111111110000111010111;
    rom[12486] = 25'b1111111111110000110001001;
    rom[12487] = 25'b1111111111110000100111100;
    rom[12488] = 25'b1111111111110000011101111;
    rom[12489] = 25'b1111111111110000010100100;
    rom[12490] = 25'b1111111111110000001011001;
    rom[12491] = 25'b1111111111110000000001110;
    rom[12492] = 25'b1111111111101111111000011;
    rom[12493] = 25'b1111111111101111101111001;
    rom[12494] = 25'b1111111111101111100110000;
    rom[12495] = 25'b1111111111101111011101000;
    rom[12496] = 25'b1111111111101111010011111;
    rom[12497] = 25'b1111111111101111001011000;
    rom[12498] = 25'b1111111111101111000010001;
    rom[12499] = 25'b1111111111101110111001010;
    rom[12500] = 25'b1111111111101110110000100;
    rom[12501] = 25'b1111111111101110100111110;
    rom[12502] = 25'b1111111111101110011111010;
    rom[12503] = 25'b1111111111101110010110101;
    rom[12504] = 25'b1111111111101110001110001;
    rom[12505] = 25'b1111111111101110000101101;
    rom[12506] = 25'b1111111111101101111101011;
    rom[12507] = 25'b1111111111101101110101001;
    rom[12508] = 25'b1111111111101101101100111;
    rom[12509] = 25'b1111111111101101100100110;
    rom[12510] = 25'b1111111111101101011100101;
    rom[12511] = 25'b1111111111101101010100100;
    rom[12512] = 25'b1111111111101101001100110;
    rom[12513] = 25'b1111111111101101000100110;
    rom[12514] = 25'b1111111111101100111101000;
    rom[12515] = 25'b1111111111101100110101010;
    rom[12516] = 25'b1111111111101100101101100;
    rom[12517] = 25'b1111111111101100100101111;
    rom[12518] = 25'b1111111111101100011110011;
    rom[12519] = 25'b1111111111101100010110111;
    rom[12520] = 25'b1111111111101100001111100;
    rom[12521] = 25'b1111111111101100001000001;
    rom[12522] = 25'b1111111111101100000000110;
    rom[12523] = 25'b1111111111101011111001101;
    rom[12524] = 25'b1111111111101011110010011;
    rom[12525] = 25'b1111111111101011101011011;
    rom[12526] = 25'b1111111111101011100100011;
    rom[12527] = 25'b1111111111101011011101011;
    rom[12528] = 25'b1111111111101011010110101;
    rom[12529] = 25'b1111111111101011001111110;
    rom[12530] = 25'b1111111111101011001001000;
    rom[12531] = 25'b1111111111101011000010010;
    rom[12532] = 25'b1111111111101010111011101;
    rom[12533] = 25'b1111111111101010110101001;
    rom[12534] = 25'b1111111111101010101110101;
    rom[12535] = 25'b1111111111101010101000010;
    rom[12536] = 25'b1111111111101010100001111;
    rom[12537] = 25'b1111111111101010011011101;
    rom[12538] = 25'b1111111111101010010101011;
    rom[12539] = 25'b1111111111101010001111010;
    rom[12540] = 25'b1111111111101010001001001;
    rom[12541] = 25'b1111111111101010000011001;
    rom[12542] = 25'b1111111111101001111101001;
    rom[12543] = 25'b1111111111101001110111011;
    rom[12544] = 25'b1111111111101001110001100;
    rom[12545] = 25'b1111111111101001101011110;
    rom[12546] = 25'b1111111111101001100110001;
    rom[12547] = 25'b1111111111101001100000100;
    rom[12548] = 25'b1111111111101001011011000;
    rom[12549] = 25'b1111111111101001010101011;
    rom[12550] = 25'b1111111111101001010000000;
    rom[12551] = 25'b1111111111101001001010101;
    rom[12552] = 25'b1111111111101001000101011;
    rom[12553] = 25'b1111111111101001000000001;
    rom[12554] = 25'b1111111111101000111011000;
    rom[12555] = 25'b1111111111101000110101111;
    rom[12556] = 25'b1111111111101000110000111;
    rom[12557] = 25'b1111111111101000101011111;
    rom[12558] = 25'b1111111111101000100111000;
    rom[12559] = 25'b1111111111101000100010001;
    rom[12560] = 25'b1111111111101000011101011;
    rom[12561] = 25'b1111111111101000011000110;
    rom[12562] = 25'b1111111111101000010100000;
    rom[12563] = 25'b1111111111101000001111100;
    rom[12564] = 25'b1111111111101000001010111;
    rom[12565] = 25'b1111111111101000000110100;
    rom[12566] = 25'b1111111111101000000010001;
    rom[12567] = 25'b1111111111100111111101110;
    rom[12568] = 25'b1111111111100111111001100;
    rom[12569] = 25'b1111111111100111110101010;
    rom[12570] = 25'b1111111111100111110001010;
    rom[12571] = 25'b1111111111100111101101001;
    rom[12572] = 25'b1111111111100111101001001;
    rom[12573] = 25'b1111111111100111100101010;
    rom[12574] = 25'b1111111111100111100001011;
    rom[12575] = 25'b1111111111100111011101100;
    rom[12576] = 25'b1111111111100111011001110;
    rom[12577] = 25'b1111111111100111010110001;
    rom[12578] = 25'b1111111111100111010010100;
    rom[12579] = 25'b1111111111100111001110111;
    rom[12580] = 25'b1111111111100111001011011;
    rom[12581] = 25'b1111111111100111001000000;
    rom[12582] = 25'b1111111111100111000100101;
    rom[12583] = 25'b1111111111100111000001011;
    rom[12584] = 25'b1111111111100110111110001;
    rom[12585] = 25'b1111111111100110111011000;
    rom[12586] = 25'b1111111111100110110111110;
    rom[12587] = 25'b1111111111100110110100110;
    rom[12588] = 25'b1111111111100110110001110;
    rom[12589] = 25'b1111111111100110101110111;
    rom[12590] = 25'b1111111111100110101100000;
    rom[12591] = 25'b1111111111100110101001001;
    rom[12592] = 25'b1111111111100110100110011;
    rom[12593] = 25'b1111111111100110100011101;
    rom[12594] = 25'b1111111111100110100001000;
    rom[12595] = 25'b1111111111100110011110100;
    rom[12596] = 25'b1111111111100110011100000;
    rom[12597] = 25'b1111111111100110011001100;
    rom[12598] = 25'b1111111111100110010111001;
    rom[12599] = 25'b1111111111100110010100110;
    rom[12600] = 25'b1111111111100110010010100;
    rom[12601] = 25'b1111111111100110010000010;
    rom[12602] = 25'b1111111111100110001110001;
    rom[12603] = 25'b1111111111100110001100000;
    rom[12604] = 25'b1111111111100110001010000;
    rom[12605] = 25'b1111111111100110001000001;
    rom[12606] = 25'b1111111111100110000110010;
    rom[12607] = 25'b1111111111100110000100010;
    rom[12608] = 25'b1111111111100110000010100;
    rom[12609] = 25'b1111111111100110000000110;
    rom[12610] = 25'b1111111111100101111111001;
    rom[12611] = 25'b1111111111100101111101100;
    rom[12612] = 25'b1111111111100101111011111;
    rom[12613] = 25'b1111111111100101111010011;
    rom[12614] = 25'b1111111111100101111001000;
    rom[12615] = 25'b1111111111100101110111101;
    rom[12616] = 25'b1111111111100101110110010;
    rom[12617] = 25'b1111111111100101110101000;
    rom[12618] = 25'b1111111111100101110011111;
    rom[12619] = 25'b1111111111100101110010101;
    rom[12620] = 25'b1111111111100101110001100;
    rom[12621] = 25'b1111111111100101110000100;
    rom[12622] = 25'b1111111111100101101111100;
    rom[12623] = 25'b1111111111100101101110100;
    rom[12624] = 25'b1111111111100101101101101;
    rom[12625] = 25'b1111111111100101101100110;
    rom[12626] = 25'b1111111111100101101100000;
    rom[12627] = 25'b1111111111100101101011011;
    rom[12628] = 25'b1111111111100101101010101;
    rom[12629] = 25'b1111111111100101101010001;
    rom[12630] = 25'b1111111111100101101001101;
    rom[12631] = 25'b1111111111100101101001001;
    rom[12632] = 25'b1111111111100101101000101;
    rom[12633] = 25'b1111111111100101101000010;
    rom[12634] = 25'b1111111111100101100111111;
    rom[12635] = 25'b1111111111100101100111110;
    rom[12636] = 25'b1111111111100101100111100;
    rom[12637] = 25'b1111111111100101100111010;
    rom[12638] = 25'b1111111111100101100111001;
    rom[12639] = 25'b1111111111100101100111000;
    rom[12640] = 25'b1111111111100101100111000;
    rom[12641] = 25'b1111111111100101100111001;
    rom[12642] = 25'b1111111111100101100111010;
    rom[12643] = 25'b1111111111100101100111011;
    rom[12644] = 25'b1111111111100101100111101;
    rom[12645] = 25'b1111111111100101100111110;
    rom[12646] = 25'b1111111111100101101000001;
    rom[12647] = 25'b1111111111100101101000100;
    rom[12648] = 25'b1111111111100101101000111;
    rom[12649] = 25'b1111111111100101101001011;
    rom[12650] = 25'b1111111111100101101001111;
    rom[12651] = 25'b1111111111100101101010100;
    rom[12652] = 25'b1111111111100101101011000;
    rom[12653] = 25'b1111111111100101101011110;
    rom[12654] = 25'b1111111111100101101100011;
    rom[12655] = 25'b1111111111100101101101001;
    rom[12656] = 25'b1111111111100101101110000;
    rom[12657] = 25'b1111111111100101101110111;
    rom[12658] = 25'b1111111111100101101111110;
    rom[12659] = 25'b1111111111100101110000110;
    rom[12660] = 25'b1111111111100101110001110;
    rom[12661] = 25'b1111111111100101110010110;
    rom[12662] = 25'b1111111111100101110011111;
    rom[12663] = 25'b1111111111100101110101000;
    rom[12664] = 25'b1111111111100101110110001;
    rom[12665] = 25'b1111111111100101110111011;
    rom[12666] = 25'b1111111111100101111000110;
    rom[12667] = 25'b1111111111100101111010001;
    rom[12668] = 25'b1111111111100101111011100;
    rom[12669] = 25'b1111111111100101111100111;
    rom[12670] = 25'b1111111111100101111110011;
    rom[12671] = 25'b1111111111100110000000000;
    rom[12672] = 25'b1111111111100110000001100;
    rom[12673] = 25'b1111111111100110000011001;
    rom[12674] = 25'b1111111111100110000100110;
    rom[12675] = 25'b1111111111100110000110100;
    rom[12676] = 25'b1111111111100110001000010;
    rom[12677] = 25'b1111111111100110001010000;
    rom[12678] = 25'b1111111111100110001011111;
    rom[12679] = 25'b1111111111100110001101110;
    rom[12680] = 25'b1111111111100110001111101;
    rom[12681] = 25'b1111111111100110010001110;
    rom[12682] = 25'b1111111111100110010011110;
    rom[12683] = 25'b1111111111100110010101110;
    rom[12684] = 25'b1111111111100110010111111;
    rom[12685] = 25'b1111111111100110011010000;
    rom[12686] = 25'b1111111111100110011100010;
    rom[12687] = 25'b1111111111100110011110100;
    rom[12688] = 25'b1111111111100110100000101;
    rom[12689] = 25'b1111111111100110100011000;
    rom[12690] = 25'b1111111111100110100101100;
    rom[12691] = 25'b1111111111100110100111110;
    rom[12692] = 25'b1111111111100110101010010;
    rom[12693] = 25'b1111111111100110101100110;
    rom[12694] = 25'b1111111111100110101111010;
    rom[12695] = 25'b1111111111100110110001111;
    rom[12696] = 25'b1111111111100110110100100;
    rom[12697] = 25'b1111111111100110110111001;
    rom[12698] = 25'b1111111111100110111001110;
    rom[12699] = 25'b1111111111100110111100100;
    rom[12700] = 25'b1111111111100110111111010;
    rom[12701] = 25'b1111111111100111000010001;
    rom[12702] = 25'b1111111111100111000100111;
    rom[12703] = 25'b1111111111100111000111110;
    rom[12704] = 25'b1111111111100111001010110;
    rom[12705] = 25'b1111111111100111001101110;
    rom[12706] = 25'b1111111111100111010000110;
    rom[12707] = 25'b1111111111100111010011111;
    rom[12708] = 25'b1111111111100111010110111;
    rom[12709] = 25'b1111111111100111011010000;
    rom[12710] = 25'b1111111111100111011101001;
    rom[12711] = 25'b1111111111100111100000010;
    rom[12712] = 25'b1111111111100111100011100;
    rom[12713] = 25'b1111111111100111100110110;
    rom[12714] = 25'b1111111111100111101010001;
    rom[12715] = 25'b1111111111100111101101100;
    rom[12716] = 25'b1111111111100111110000111;
    rom[12717] = 25'b1111111111100111110100010;
    rom[12718] = 25'b1111111111100111110111101;
    rom[12719] = 25'b1111111111100111111011001;
    rom[12720] = 25'b1111111111100111111110101;
    rom[12721] = 25'b1111111111101000000010001;
    rom[12722] = 25'b1111111111101000000101110;
    rom[12723] = 25'b1111111111101000001001011;
    rom[12724] = 25'b1111111111101000001101000;
    rom[12725] = 25'b1111111111101000010000110;
    rom[12726] = 25'b1111111111101000010100011;
    rom[12727] = 25'b1111111111101000011000001;
    rom[12728] = 25'b1111111111101000011011111;
    rom[12729] = 25'b1111111111101000011111110;
    rom[12730] = 25'b1111111111101000100011100;
    rom[12731] = 25'b1111111111101000100111100;
    rom[12732] = 25'b1111111111101000101011011;
    rom[12733] = 25'b1111111111101000101111011;
    rom[12734] = 25'b1111111111101000110011010;
    rom[12735] = 25'b1111111111101000110111011;
    rom[12736] = 25'b1111111111101000111011010;
    rom[12737] = 25'b1111111111101000111111011;
    rom[12738] = 25'b1111111111101001000011100;
    rom[12739] = 25'b1111111111101001000111101;
    rom[12740] = 25'b1111111111101001001011110;
    rom[12741] = 25'b1111111111101001001111111;
    rom[12742] = 25'b1111111111101001010100001;
    rom[12743] = 25'b1111111111101001011000011;
    rom[12744] = 25'b1111111111101001011100101;
    rom[12745] = 25'b1111111111101001100000111;
    rom[12746] = 25'b1111111111101001100101010;
    rom[12747] = 25'b1111111111101001101001101;
    rom[12748] = 25'b1111111111101001101110000;
    rom[12749] = 25'b1111111111101001110010011;
    rom[12750] = 25'b1111111111101001110110111;
    rom[12751] = 25'b1111111111101001111011011;
    rom[12752] = 25'b1111111111101001111111111;
    rom[12753] = 25'b1111111111101010000100010;
    rom[12754] = 25'b1111111111101010001000111;
    rom[12755] = 25'b1111111111101010001101100;
    rom[12756] = 25'b1111111111101010010010000;
    rom[12757] = 25'b1111111111101010010110110;
    rom[12758] = 25'b1111111111101010011011010;
    rom[12759] = 25'b1111111111101010100000000;
    rom[12760] = 25'b1111111111101010100100110;
    rom[12761] = 25'b1111111111101010101001011;
    rom[12762] = 25'b1111111111101010101110001;
    rom[12763] = 25'b1111111111101010110010111;
    rom[12764] = 25'b1111111111101010110111110;
    rom[12765] = 25'b1111111111101010111100100;
    rom[12766] = 25'b1111111111101011000001011;
    rom[12767] = 25'b1111111111101011000110010;
    rom[12768] = 25'b1111111111101011001011001;
    rom[12769] = 25'b1111111111101011010000000;
    rom[12770] = 25'b1111111111101011010101000;
    rom[12771] = 25'b1111111111101011011001111;
    rom[12772] = 25'b1111111111101011011110111;
    rom[12773] = 25'b1111111111101011100011111;
    rom[12774] = 25'b1111111111101011101000111;
    rom[12775] = 25'b1111111111101011101110000;
    rom[12776] = 25'b1111111111101011110011000;
    rom[12777] = 25'b1111111111101011111000001;
    rom[12778] = 25'b1111111111101011111101001;
    rom[12779] = 25'b1111111111101100000010010;
    rom[12780] = 25'b1111111111101100000111100;
    rom[12781] = 25'b1111111111101100001100101;
    rom[12782] = 25'b1111111111101100010001110;
    rom[12783] = 25'b1111111111101100010111000;
    rom[12784] = 25'b1111111111101100011100010;
    rom[12785] = 25'b1111111111101100100001011;
    rom[12786] = 25'b1111111111101100100110110;
    rom[12787] = 25'b1111111111101100101100000;
    rom[12788] = 25'b1111111111101100110001010;
    rom[12789] = 25'b1111111111101100110110101;
    rom[12790] = 25'b1111111111101100111011111;
    rom[12791] = 25'b1111111111101101000001011;
    rom[12792] = 25'b1111111111101101000110101;
    rom[12793] = 25'b1111111111101101001100000;
    rom[12794] = 25'b1111111111101101010001100;
    rom[12795] = 25'b1111111111101101010110111;
    rom[12796] = 25'b1111111111101101011100011;
    rom[12797] = 25'b1111111111101101100001110;
    rom[12798] = 25'b1111111111101101100111001;
    rom[12799] = 25'b1111111111101101101100110;
    rom[12800] = 25'b1111111111101101110010001;
    rom[12801] = 25'b1111111111101101110111101;
    rom[12802] = 25'b1111111111101101111101001;
    rom[12803] = 25'b1111111111101110000010110;
    rom[12804] = 25'b1111111111101110001000011;
    rom[12805] = 25'b1111111111101110001101111;
    rom[12806] = 25'b1111111111101110010011011;
    rom[12807] = 25'b1111111111101110011001000;
    rom[12808] = 25'b1111111111101110011110101;
    rom[12809] = 25'b1111111111101110100100010;
    rom[12810] = 25'b1111111111101110101001111;
    rom[12811] = 25'b1111111111101110101111101;
    rom[12812] = 25'b1111111111101110110101010;
    rom[12813] = 25'b1111111111101110111010111;
    rom[12814] = 25'b1111111111101111000000101;
    rom[12815] = 25'b1111111111101111000110010;
    rom[12816] = 25'b1111111111101111001100000;
    rom[12817] = 25'b1111111111101111010001110;
    rom[12818] = 25'b1111111111101111010111011;
    rom[12819] = 25'b1111111111101111011101001;
    rom[12820] = 25'b1111111111101111100010111;
    rom[12821] = 25'b1111111111101111101000101;
    rom[12822] = 25'b1111111111101111101110011;
    rom[12823] = 25'b1111111111101111110100010;
    rom[12824] = 25'b1111111111101111111010000;
    rom[12825] = 25'b1111111111101111111111111;
    rom[12826] = 25'b1111111111110000000101101;
    rom[12827] = 25'b1111111111110000001011011;
    rom[12828] = 25'b1111111111110000010001010;
    rom[12829] = 25'b1111111111110000010111001;
    rom[12830] = 25'b1111111111110000011101000;
    rom[12831] = 25'b1111111111110000100010110;
    rom[12832] = 25'b1111111111110000101000101;
    rom[12833] = 25'b1111111111110000101110100;
    rom[12834] = 25'b1111111111110000110100011;
    rom[12835] = 25'b1111111111110000111010010;
    rom[12836] = 25'b1111111111110001000000001;
    rom[12837] = 25'b1111111111110001000110000;
    rom[12838] = 25'b1111111111110001001100000;
    rom[12839] = 25'b1111111111110001010001111;
    rom[12840] = 25'b1111111111110001010111110;
    rom[12841] = 25'b1111111111110001011101110;
    rom[12842] = 25'b1111111111110001100011101;
    rom[12843] = 25'b1111111111110001101001100;
    rom[12844] = 25'b1111111111110001101111100;
    rom[12845] = 25'b1111111111110001110101011;
    rom[12846] = 25'b1111111111110001111011011;
    rom[12847] = 25'b1111111111110010000001011;
    rom[12848] = 25'b1111111111110010000111010;
    rom[12849] = 25'b1111111111110010001101010;
    rom[12850] = 25'b1111111111110010010011001;
    rom[12851] = 25'b1111111111110010011001010;
    rom[12852] = 25'b1111111111110010011111010;
    rom[12853] = 25'b1111111111110010100101001;
    rom[12854] = 25'b1111111111110010101011001;
    rom[12855] = 25'b1111111111110010110001001;
    rom[12856] = 25'b1111111111110010110111001;
    rom[12857] = 25'b1111111111110010111101001;
    rom[12858] = 25'b1111111111110011000011001;
    rom[12859] = 25'b1111111111110011001001001;
    rom[12860] = 25'b1111111111110011001111000;
    rom[12861] = 25'b1111111111110011010101001;
    rom[12862] = 25'b1111111111110011011011000;
    rom[12863] = 25'b1111111111110011100001001;
    rom[12864] = 25'b1111111111110011100111000;
    rom[12865] = 25'b1111111111110011101101001;
    rom[12866] = 25'b1111111111110011110011001;
    rom[12867] = 25'b1111111111110011111001001;
    rom[12868] = 25'b1111111111110011111111001;
    rom[12869] = 25'b1111111111110100000101001;
    rom[12870] = 25'b1111111111110100001011001;
    rom[12871] = 25'b1111111111110100010001001;
    rom[12872] = 25'b1111111111110100010111001;
    rom[12873] = 25'b1111111111110100011101001;
    rom[12874] = 25'b1111111111110100100011001;
    rom[12875] = 25'b1111111111110100101001001;
    rom[12876] = 25'b1111111111110100101111001;
    rom[12877] = 25'b1111111111110100110101010;
    rom[12878] = 25'b1111111111110100111011001;
    rom[12879] = 25'b1111111111110101000001010;
    rom[12880] = 25'b1111111111110101000111001;
    rom[12881] = 25'b1111111111110101001101001;
    rom[12882] = 25'b1111111111110101010011001;
    rom[12883] = 25'b1111111111110101011001001;
    rom[12884] = 25'b1111111111110101011111010;
    rom[12885] = 25'b1111111111110101100101001;
    rom[12886] = 25'b1111111111110101101011001;
    rom[12887] = 25'b1111111111110101110001000;
    rom[12888] = 25'b1111111111110101110111001;
    rom[12889] = 25'b1111111111110101111101001;
    rom[12890] = 25'b1111111111110110000011000;
    rom[12891] = 25'b1111111111110110001001000;
    rom[12892] = 25'b1111111111110110001110111;
    rom[12893] = 25'b1111111111110110010100111;
    rom[12894] = 25'b1111111111110110011010111;
    rom[12895] = 25'b1111111111110110100000110;
    rom[12896] = 25'b1111111111110110100110110;
    rom[12897] = 25'b1111111111110110101100110;
    rom[12898] = 25'b1111111111110110110010101;
    rom[12899] = 25'b1111111111110110111000101;
    rom[12900] = 25'b1111111111110110111110100;
    rom[12901] = 25'b1111111111110111000100011;
    rom[12902] = 25'b1111111111110111001010011;
    rom[12903] = 25'b1111111111110111010000010;
    rom[12904] = 25'b1111111111110111010110001;
    rom[12905] = 25'b1111111111110111011100000;
    rom[12906] = 25'b1111111111110111100010000;
    rom[12907] = 25'b1111111111110111100111110;
    rom[12908] = 25'b1111111111110111101101101;
    rom[12909] = 25'b1111111111110111110011101;
    rom[12910] = 25'b1111111111110111111001100;
    rom[12911] = 25'b1111111111110111111111010;
    rom[12912] = 25'b1111111111111000000101001;
    rom[12913] = 25'b1111111111111000001011000;
    rom[12914] = 25'b1111111111111000010000111;
    rom[12915] = 25'b1111111111111000010110110;
    rom[12916] = 25'b1111111111111000011100011;
    rom[12917] = 25'b1111111111111000100010010;
    rom[12918] = 25'b1111111111111000101000001;
    rom[12919] = 25'b1111111111111000101101111;
    rom[12920] = 25'b1111111111111000110011110;
    rom[12921] = 25'b1111111111111000111001100;
    rom[12922] = 25'b1111111111111000111111010;
    rom[12923] = 25'b1111111111111001000100111;
    rom[12924] = 25'b1111111111111001001010101;
    rom[12925] = 25'b1111111111111001010000011;
    rom[12926] = 25'b1111111111111001010110001;
    rom[12927] = 25'b1111111111111001011011111;
    rom[12928] = 25'b1111111111111001100001101;
    rom[12929] = 25'b1111111111111001100111010;
    rom[12930] = 25'b1111111111111001101101000;
    rom[12931] = 25'b1111111111111001110010101;
    rom[12932] = 25'b1111111111111001111000011;
    rom[12933] = 25'b1111111111111001111110000;
    rom[12934] = 25'b1111111111111010000011101;
    rom[12935] = 25'b1111111111111010001001010;
    rom[12936] = 25'b1111111111111010001110111;
    rom[12937] = 25'b1111111111111010010100100;
    rom[12938] = 25'b1111111111111010011010010;
    rom[12939] = 25'b1111111111111010011111111;
    rom[12940] = 25'b1111111111111010100101011;
    rom[12941] = 25'b1111111111111010101010111;
    rom[12942] = 25'b1111111111111010110000100;
    rom[12943] = 25'b1111111111111010110110000;
    rom[12944] = 25'b1111111111111010111011101;
    rom[12945] = 25'b1111111111111011000001001;
    rom[12946] = 25'b1111111111111011000110101;
    rom[12947] = 25'b1111111111111011001100001;
    rom[12948] = 25'b1111111111111011010001101;
    rom[12949] = 25'b1111111111111011010111001;
    rom[12950] = 25'b1111111111111011011100100;
    rom[12951] = 25'b1111111111111011100010001;
    rom[12952] = 25'b1111111111111011100111100;
    rom[12953] = 25'b1111111111111011101100111;
    rom[12954] = 25'b1111111111111011110010011;
    rom[12955] = 25'b1111111111111011110111101;
    rom[12956] = 25'b1111111111111011111101001;
    rom[12957] = 25'b1111111111111100000010100;
    rom[12958] = 25'b1111111111111100000111110;
    rom[12959] = 25'b1111111111111100001101001;
    rom[12960] = 25'b1111111111111100010010011;
    rom[12961] = 25'b1111111111111100010111110;
    rom[12962] = 25'b1111111111111100011101001;
    rom[12963] = 25'b1111111111111100100010011;
    rom[12964] = 25'b1111111111111100100111110;
    rom[12965] = 25'b1111111111111100101100111;
    rom[12966] = 25'b1111111111111100110010010;
    rom[12967] = 25'b1111111111111100110111011;
    rom[12968] = 25'b1111111111111100111100101;
    rom[12969] = 25'b1111111111111101000001111;
    rom[12970] = 25'b1111111111111101000111000;
    rom[12971] = 25'b1111111111111101001100001;
    rom[12972] = 25'b1111111111111101010001011;
    rom[12973] = 25'b1111111111111101010110100;
    rom[12974] = 25'b1111111111111101011011101;
    rom[12975] = 25'b1111111111111101100000101;
    rom[12976] = 25'b1111111111111101100101110;
    rom[12977] = 25'b1111111111111101101010111;
    rom[12978] = 25'b1111111111111101110000000;
    rom[12979] = 25'b1111111111111101110101000;
    rom[12980] = 25'b1111111111111101111010000;
    rom[12981] = 25'b1111111111111101111111000;
    rom[12982] = 25'b1111111111111110000100000;
    rom[12983] = 25'b1111111111111110001001000;
    rom[12984] = 25'b1111111111111110001110000;
    rom[12985] = 25'b1111111111111110010011000;
    rom[12986] = 25'b1111111111111110010111111;
    rom[12987] = 25'b1111111111111110011100110;
    rom[12988] = 25'b1111111111111110100001101;
    rom[12989] = 25'b1111111111111110100110100;
    rom[12990] = 25'b1111111111111110101011011;
    rom[12991] = 25'b1111111111111110110000010;
    rom[12992] = 25'b1111111111111110110101001;
    rom[12993] = 25'b1111111111111110111001111;
    rom[12994] = 25'b1111111111111110111110101;
    rom[12995] = 25'b1111111111111111000011100;
    rom[12996] = 25'b1111111111111111001000010;
    rom[12997] = 25'b1111111111111111001101000;
    rom[12998] = 25'b1111111111111111010001110;
    rom[12999] = 25'b1111111111111111010110100;
    rom[13000] = 25'b1111111111111111011011001;
    rom[13001] = 25'b1111111111111111011111111;
    rom[13002] = 25'b1111111111111111100100011;
    rom[13003] = 25'b1111111111111111101001001;
    rom[13004] = 25'b1111111111111111101101101;
    rom[13005] = 25'b1111111111111111110010011;
    rom[13006] = 25'b1111111111111111110110111;
    rom[13007] = 25'b1111111111111111111011100;
    rom[13008] = 25'b0000000000000000000000000;
    rom[13009] = 25'b0000000000000000000100011;
    rom[13010] = 25'b0000000000000000001001000;
    rom[13011] = 25'b0000000000000000001101100;
    rom[13012] = 25'b0000000000000000010001111;
    rom[13013] = 25'b0000000000000000010110011;
    rom[13014] = 25'b0000000000000000011010110;
    rom[13015] = 25'b0000000000000000011111010;
    rom[13016] = 25'b0000000000000000100011100;
    rom[13017] = 25'b0000000000000000100111111;
    rom[13018] = 25'b0000000000000000101100010;
    rom[13019] = 25'b0000000000000000110000101;
    rom[13020] = 25'b0000000000000000110101000;
    rom[13021] = 25'b0000000000000000111001010;
    rom[13022] = 25'b0000000000000000111101101;
    rom[13023] = 25'b0000000000000001000001111;
    rom[13024] = 25'b0000000000000001000110001;
    rom[13025] = 25'b0000000000000001001010010;
    rom[13026] = 25'b0000000000000001001110100;
    rom[13027] = 25'b0000000000000001010010101;
    rom[13028] = 25'b0000000000000001010110110;
    rom[13029] = 25'b0000000000000001011011000;
    rom[13030] = 25'b0000000000000001011111001;
    rom[13031] = 25'b0000000000000001100011010;
    rom[13032] = 25'b0000000000000001100111010;
    rom[13033] = 25'b0000000000000001101011011;
    rom[13034] = 25'b0000000000000001101111011;
    rom[13035] = 25'b0000000000000001110011011;
    rom[13036] = 25'b0000000000000001110111011;
    rom[13037] = 25'b0000000000000001111011011;
    rom[13038] = 25'b0000000000000001111111011;
    rom[13039] = 25'b0000000000000010000011011;
    rom[13040] = 25'b0000000000000010000111010;
    rom[13041] = 25'b0000000000000010001011001;
    rom[13042] = 25'b0000000000000010001111000;
    rom[13043] = 25'b0000000000000010010010111;
    rom[13044] = 25'b0000000000000010010110110;
    rom[13045] = 25'b0000000000000010011010100;
    rom[13046] = 25'b0000000000000010011110011;
    rom[13047] = 25'b0000000000000010100010001;
    rom[13048] = 25'b0000000000000010100101111;
    rom[13049] = 25'b0000000000000010101001101;
    rom[13050] = 25'b0000000000000010101101011;
    rom[13051] = 25'b0000000000000010110001000;
    rom[13052] = 25'b0000000000000010110100110;
    rom[13053] = 25'b0000000000000010111000011;
    rom[13054] = 25'b0000000000000010111100000;
    rom[13055] = 25'b0000000000000010111111101;
    rom[13056] = 25'b0000000000000011000011010;
    rom[13057] = 25'b0000000000000011000110111;
    rom[13058] = 25'b0000000000000011001010011;
    rom[13059] = 25'b0000000000000011001101111;
    rom[13060] = 25'b0000000000000011010001011;
    rom[13061] = 25'b0000000000000011010100111;
    rom[13062] = 25'b0000000000000011011000011;
    rom[13063] = 25'b0000000000000011011011110;
    rom[13064] = 25'b0000000000000011011111010;
    rom[13065] = 25'b0000000000000011100010101;
    rom[13066] = 25'b0000000000000011100110000;
    rom[13067] = 25'b0000000000000011101001011;
    rom[13068] = 25'b0000000000000011101100110;
    rom[13069] = 25'b0000000000000011110000000;
    rom[13070] = 25'b0000000000000011110011011;
    rom[13071] = 25'b0000000000000011110110101;
    rom[13072] = 25'b0000000000000011111001111;
    rom[13073] = 25'b0000000000000011111101001;
    rom[13074] = 25'b0000000000000100000000011;
    rom[13075] = 25'b0000000000000100000011100;
    rom[13076] = 25'b0000000000000100000110101;
    rom[13077] = 25'b0000000000000100001001111;
    rom[13078] = 25'b0000000000000100001101000;
    rom[13079] = 25'b0000000000000100010000001;
    rom[13080] = 25'b0000000000000100010011001;
    rom[13081] = 25'b0000000000000100010110010;
    rom[13082] = 25'b0000000000000100011001010;
    rom[13083] = 25'b0000000000000100011100011;
    rom[13084] = 25'b0000000000000100011111010;
    rom[13085] = 25'b0000000000000100100010010;
    rom[13086] = 25'b0000000000000100100101010;
    rom[13087] = 25'b0000000000000100101000001;
    rom[13088] = 25'b0000000000000100101011001;
    rom[13089] = 25'b0000000000000100101110000;
    rom[13090] = 25'b0000000000000100110000111;
    rom[13091] = 25'b0000000000000100110011110;
    rom[13092] = 25'b0000000000000100110110100;
    rom[13093] = 25'b0000000000000100111001011;
    rom[13094] = 25'b0000000000000100111100001;
    rom[13095] = 25'b0000000000000100111110111;
    rom[13096] = 25'b0000000000000101000001101;
    rom[13097] = 25'b0000000000000101000100010;
    rom[13098] = 25'b0000000000000101000111000;
    rom[13099] = 25'b0000000000000101001001110;
    rom[13100] = 25'b0000000000000101001100011;
    rom[13101] = 25'b0000000000000101001111000;
    rom[13102] = 25'b0000000000000101010001101;
    rom[13103] = 25'b0000000000000101010100001;
    rom[13104] = 25'b0000000000000101010110110;
    rom[13105] = 25'b0000000000000101011001011;
    rom[13106] = 25'b0000000000000101011011110;
    rom[13107] = 25'b0000000000000101011110011;
    rom[13108] = 25'b0000000000000101100000110;
    rom[13109] = 25'b0000000000000101100011010;
    rom[13110] = 25'b0000000000000101100101101;
    rom[13111] = 25'b0000000000000101101000001;
    rom[13112] = 25'b0000000000000101101010101;
    rom[13113] = 25'b0000000000000101101100111;
    rom[13114] = 25'b0000000000000101101111010;
    rom[13115] = 25'b0000000000000101110001101;
    rom[13116] = 25'b0000000000000101110011111;
    rom[13117] = 25'b0000000000000101110110001;
    rom[13118] = 25'b0000000000000101111000100;
    rom[13119] = 25'b0000000000000101111010110;
    rom[13120] = 25'b0000000000000101111101000;
    rom[13121] = 25'b0000000000000101111111010;
    rom[13122] = 25'b0000000000000110000001011;
    rom[13123] = 25'b0000000000000110000011100;
    rom[13124] = 25'b0000000000000110000101101;
    rom[13125] = 25'b0000000000000110000111110;
    rom[13126] = 25'b0000000000000110001001111;
    rom[13127] = 25'b0000000000000110001100000;
    rom[13128] = 25'b0000000000000110001110000;
    rom[13129] = 25'b0000000000000110010000000;
    rom[13130] = 25'b0000000000000110010010000;
    rom[13131] = 25'b0000000000000110010100000;
    rom[13132] = 25'b0000000000000110010110000;
    rom[13133] = 25'b0000000000000110011000000;
    rom[13134] = 25'b0000000000000110011001111;
    rom[13135] = 25'b0000000000000110011011110;
    rom[13136] = 25'b0000000000000110011101110;
    rom[13137] = 25'b0000000000000110011111100;
    rom[13138] = 25'b0000000000000110100001011;
    rom[13139] = 25'b0000000000000110100011010;
    rom[13140] = 25'b0000000000000110100101000;
    rom[13141] = 25'b0000000000000110100110111;
    rom[13142] = 25'b0000000000000110101000100;
    rom[13143] = 25'b0000000000000110101010010;
    rom[13144] = 25'b0000000000000110101100000;
    rom[13145] = 25'b0000000000000110101101110;
    rom[13146] = 25'b0000000000000110101111011;
    rom[13147] = 25'b0000000000000110110001000;
    rom[13148] = 25'b0000000000000110110010101;
    rom[13149] = 25'b0000000000000110110100011;
    rom[13150] = 25'b0000000000000110110110000;
    rom[13151] = 25'b0000000000000110110111011;
    rom[13152] = 25'b0000000000000110111001000;
    rom[13153] = 25'b0000000000000110111010100;
    rom[13154] = 25'b0000000000000110111100001;
    rom[13155] = 25'b0000000000000110111101101;
    rom[13156] = 25'b0000000000000110111111001;
    rom[13157] = 25'b0000000000000111000000100;
    rom[13158] = 25'b0000000000000111000010000;
    rom[13159] = 25'b0000000000000111000011011;
    rom[13160] = 25'b0000000000000111000100110;
    rom[13161] = 25'b0000000000000111000110001;
    rom[13162] = 25'b0000000000000111000111100;
    rom[13163] = 25'b0000000000000111001000110;
    rom[13164] = 25'b0000000000000111001010001;
    rom[13165] = 25'b0000000000000111001011011;
    rom[13166] = 25'b0000000000000111001100110;
    rom[13167] = 25'b0000000000000111001101111;
    rom[13168] = 25'b0000000000000111001111001;
    rom[13169] = 25'b0000000000000111010000010;
    rom[13170] = 25'b0000000000000111010001101;
    rom[13171] = 25'b0000000000000111010010110;
    rom[13172] = 25'b0000000000000111010011111;
    rom[13173] = 25'b0000000000000111010101000;
    rom[13174] = 25'b0000000000000111010110001;
    rom[13175] = 25'b0000000000000111010111010;
    rom[13176] = 25'b0000000000000111011000010;
    rom[13177] = 25'b0000000000000111011001011;
    rom[13178] = 25'b0000000000000111011010011;
    rom[13179] = 25'b0000000000000111011011011;
    rom[13180] = 25'b0000000000000111011100011;
    rom[13181] = 25'b0000000000000111011101011;
    rom[13182] = 25'b0000000000000111011110011;
    rom[13183] = 25'b0000000000000111011111010;
    rom[13184] = 25'b0000000000000111100000001;
    rom[13185] = 25'b0000000000000111100001001;
    rom[13186] = 25'b0000000000000111100010000;
    rom[13187] = 25'b0000000000000111100010110;
    rom[13188] = 25'b0000000000000111100011101;
    rom[13189] = 25'b0000000000000111100100100;
    rom[13190] = 25'b0000000000000111100101010;
    rom[13191] = 25'b0000000000000111100110000;
    rom[13192] = 25'b0000000000000111100110111;
    rom[13193] = 25'b0000000000000111100111101;
    rom[13194] = 25'b0000000000000111101000011;
    rom[13195] = 25'b0000000000000111101001000;
    rom[13196] = 25'b0000000000000111101001110;
    rom[13197] = 25'b0000000000000111101010011;
    rom[13198] = 25'b0000000000000111101011000;
    rom[13199] = 25'b0000000000000111101011101;
    rom[13200] = 25'b0000000000000111101100010;
    rom[13201] = 25'b0000000000000111101100111;
    rom[13202] = 25'b0000000000000111101101100;
    rom[13203] = 25'b0000000000000111101110000;
    rom[13204] = 25'b0000000000000111101110101;
    rom[13205] = 25'b0000000000000111101111000;
    rom[13206] = 25'b0000000000000111101111101;
    rom[13207] = 25'b0000000000000111110000001;
    rom[13208] = 25'b0000000000000111110000100;
    rom[13209] = 25'b0000000000000111110001000;
    rom[13210] = 25'b0000000000000111110001100;
    rom[13211] = 25'b0000000000000111110001111;
    rom[13212] = 25'b0000000000000111110010010;
    rom[13213] = 25'b0000000000000111110010101;
    rom[13214] = 25'b0000000000000111110011000;
    rom[13215] = 25'b0000000000000111110011011;
    rom[13216] = 25'b0000000000000111110011110;
    rom[13217] = 25'b0000000000000111110100000;
    rom[13218] = 25'b0000000000000111110100011;
    rom[13219] = 25'b0000000000000111110100100;
    rom[13220] = 25'b0000000000000111110100111;
    rom[13221] = 25'b0000000000000111110101001;
    rom[13222] = 25'b0000000000000111110101010;
    rom[13223] = 25'b0000000000000111110101100;
    rom[13224] = 25'b0000000000000111110101110;
    rom[13225] = 25'b0000000000000111110110000;
    rom[13226] = 25'b0000000000000111110110000;
    rom[13227] = 25'b0000000000000111110110010;
    rom[13228] = 25'b0000000000000111110110011;
    rom[13229] = 25'b0000000000000111110110100;
    rom[13230] = 25'b0000000000000111110110101;
    rom[13231] = 25'b0000000000000111110110101;
    rom[13232] = 25'b0000000000000111110110110;
    rom[13233] = 25'b0000000000000111110110110;
    rom[13234] = 25'b0000000000000111110110110;
    rom[13235] = 25'b0000000000000111110110110;
    rom[13236] = 25'b0000000000000111110110110;
    rom[13237] = 25'b0000000000000111110110110;
    rom[13238] = 25'b0000000000000111110110110;
    rom[13239] = 25'b0000000000000111110110110;
    rom[13240] = 25'b0000000000000111110110101;
    rom[13241] = 25'b0000000000000111110110100;
    rom[13242] = 25'b0000000000000111110110011;
    rom[13243] = 25'b0000000000000111110110010;
    rom[13244] = 25'b0000000000000111110110001;
    rom[13245] = 25'b0000000000000111110110000;
    rom[13246] = 25'b0000000000000111110101111;
    rom[13247] = 25'b0000000000000111110101110;
    rom[13248] = 25'b0000000000000111110101100;
    rom[13249] = 25'b0000000000000111110101010;
    rom[13250] = 25'b0000000000000111110101001;
    rom[13251] = 25'b0000000000000111110100111;
    rom[13252] = 25'b0000000000000111110100100;
    rom[13253] = 25'b0000000000000111110100011;
    rom[13254] = 25'b0000000000000111110100000;
    rom[13255] = 25'b0000000000000111110011110;
    rom[13256] = 25'b0000000000000111110011011;
    rom[13257] = 25'b0000000000000111110011001;
    rom[13258] = 25'b0000000000000111110010110;
    rom[13259] = 25'b0000000000000111110010011;
    rom[13260] = 25'b0000000000000111110010000;
    rom[13261] = 25'b0000000000000111110001110;
    rom[13262] = 25'b0000000000000111110001010;
    rom[13263] = 25'b0000000000000111110000111;
    rom[13264] = 25'b0000000000000111110000011;
    rom[13265] = 25'b0000000000000111110000000;
    rom[13266] = 25'b0000000000000111101111100;
    rom[13267] = 25'b0000000000000111101111000;
    rom[13268] = 25'b0000000000000111101110101;
    rom[13269] = 25'b0000000000000111101110001;
    rom[13270] = 25'b0000000000000111101101100;
    rom[13271] = 25'b0000000000000111101101000;
    rom[13272] = 25'b0000000000000111101100100;
    rom[13273] = 25'b0000000000000111101100000;
    rom[13274] = 25'b0000000000000111101011011;
    rom[13275] = 25'b0000000000000111101010110;
    rom[13276] = 25'b0000000000000111101010010;
    rom[13277] = 25'b0000000000000111101001101;
    rom[13278] = 25'b0000000000000111101001000;
    rom[13279] = 25'b0000000000000111101000011;
    rom[13280] = 25'b0000000000000111100111110;
    rom[13281] = 25'b0000000000000111100111000;
    rom[13282] = 25'b0000000000000111100110011;
    rom[13283] = 25'b0000000000000111100101101;
    rom[13284] = 25'b0000000000000111100101000;
    rom[13285] = 25'b0000000000000111100100010;
    rom[13286] = 25'b0000000000000111100011100;
    rom[13287] = 25'b0000000000000111100010110;
    rom[13288] = 25'b0000000000000111100010001;
    rom[13289] = 25'b0000000000000111100001011;
    rom[13290] = 25'b0000000000000111100000101;
    rom[13291] = 25'b0000000000000111011111111;
    rom[13292] = 25'b0000000000000111011111000;
    rom[13293] = 25'b0000000000000111011110010;
    rom[13294] = 25'b0000000000000111011101011;
    rom[13295] = 25'b0000000000000111011100100;
    rom[13296] = 25'b0000000000000111011011101;
    rom[13297] = 25'b0000000000000111011010111;
    rom[13298] = 25'b0000000000000111011010000;
    rom[13299] = 25'b0000000000000111011001001;
    rom[13300] = 25'b0000000000000111011000010;
    rom[13301] = 25'b0000000000000111010111011;
    rom[13302] = 25'b0000000000000111010110100;
    rom[13303] = 25'b0000000000000111010101100;
    rom[13304] = 25'b0000000000000111010100100;
    rom[13305] = 25'b0000000000000111010011101;
    rom[13306] = 25'b0000000000000111010010101;
    rom[13307] = 25'b0000000000000111010001110;
    rom[13308] = 25'b0000000000000111010000110;
    rom[13309] = 25'b0000000000000111001111110;
    rom[13310] = 25'b0000000000000111001110110;
    rom[13311] = 25'b0000000000000111001101110;
    rom[13312] = 25'b0000000000000111001100110;
    rom[13313] = 25'b0000000000000111001011110;
    rom[13314] = 25'b0000000000000111001010101;
    rom[13315] = 25'b0000000000000111001001101;
    rom[13316] = 25'b0000000000000111001000100;
    rom[13317] = 25'b0000000000000111000111100;
    rom[13318] = 25'b0000000000000111000110011;
    rom[13319] = 25'b0000000000000111000101011;
    rom[13320] = 25'b0000000000000111000100010;
    rom[13321] = 25'b0000000000000111000011001;
    rom[13322] = 25'b0000000000000111000010000;
    rom[13323] = 25'b0000000000000111000000111;
    rom[13324] = 25'b0000000000000110111111110;
    rom[13325] = 25'b0000000000000110111110100;
    rom[13326] = 25'b0000000000000110111101011;
    rom[13327] = 25'b0000000000000110111100010;
    rom[13328] = 25'b0000000000000110111011000;
    rom[13329] = 25'b0000000000000110111001111;
    rom[13330] = 25'b0000000000000110111000110;
    rom[13331] = 25'b0000000000000110110111100;
    rom[13332] = 25'b0000000000000110110110010;
    rom[13333] = 25'b0000000000000110110101001;
    rom[13334] = 25'b0000000000000110110011111;
    rom[13335] = 25'b0000000000000110110010100;
    rom[13336] = 25'b0000000000000110110001011;
    rom[13337] = 25'b0000000000000110110000001;
    rom[13338] = 25'b0000000000000110101110111;
    rom[13339] = 25'b0000000000000110101101100;
    rom[13340] = 25'b0000000000000110101100010;
    rom[13341] = 25'b0000000000000110101011000;
    rom[13342] = 25'b0000000000000110101001110;
    rom[13343] = 25'b0000000000000110101000011;
    rom[13344] = 25'b0000000000000110100111000;
    rom[13345] = 25'b0000000000000110100101110;
    rom[13346] = 25'b0000000000000110100100011;
    rom[13347] = 25'b0000000000000110100011001;
    rom[13348] = 25'b0000000000000110100001110;
    rom[13349] = 25'b0000000000000110100000011;
    rom[13350] = 25'b0000000000000110011111000;
    rom[13351] = 25'b0000000000000110011101101;
    rom[13352] = 25'b0000000000000110011100011;
    rom[13353] = 25'b0000000000000110011011000;
    rom[13354] = 25'b0000000000000110011001100;
    rom[13355] = 25'b0000000000000110011000001;
    rom[13356] = 25'b0000000000000110010110110;
    rom[13357] = 25'b0000000000000110010101010;
    rom[13358] = 25'b0000000000000110010011111;
    rom[13359] = 25'b0000000000000110010010011;
    rom[13360] = 25'b0000000000000110010001000;
    rom[13361] = 25'b0000000000000110001111101;
    rom[13362] = 25'b0000000000000110001110001;
    rom[13363] = 25'b0000000000000110001100110;
    rom[13364] = 25'b0000000000000110001011010;
    rom[13365] = 25'b0000000000000110001001110;
    rom[13366] = 25'b0000000000000110001000011;
    rom[13367] = 25'b0000000000000110000110111;
    rom[13368] = 25'b0000000000000110000101011;
    rom[13369] = 25'b0000000000000110000011111;
    rom[13370] = 25'b0000000000000110000010011;
    rom[13371] = 25'b0000000000000110000000110;
    rom[13372] = 25'b0000000000000101111111010;
    rom[13373] = 25'b0000000000000101111101110;
    rom[13374] = 25'b0000000000000101111100011;
    rom[13375] = 25'b0000000000000101111010110;
    rom[13376] = 25'b0000000000000101111001010;
    rom[13377] = 25'b0000000000000101110111110;
    rom[13378] = 25'b0000000000000101110110001;
    rom[13379] = 25'b0000000000000101110100100;
    rom[13380] = 25'b0000000000000101110011001;
    rom[13381] = 25'b0000000000000101110001100;
    rom[13382] = 25'b0000000000000101110000000;
    rom[13383] = 25'b0000000000000101101110011;
    rom[13384] = 25'b0000000000000101101100110;
    rom[13385] = 25'b0000000000000101101011010;
    rom[13386] = 25'b0000000000000101101001101;
    rom[13387] = 25'b0000000000000101101000000;
    rom[13388] = 25'b0000000000000101100110011;
    rom[13389] = 25'b0000000000000101100100111;
    rom[13390] = 25'b0000000000000101100011010;
    rom[13391] = 25'b0000000000000101100001101;
    rom[13392] = 25'b0000000000000101100000000;
    rom[13393] = 25'b0000000000000101011110100;
    rom[13394] = 25'b0000000000000101011100111;
    rom[13395] = 25'b0000000000000101011011001;
    rom[13396] = 25'b0000000000000101011001100;
    rom[13397] = 25'b0000000000000101011000000;
    rom[13398] = 25'b0000000000000101010110010;
    rom[13399] = 25'b0000000000000101010100101;
    rom[13400] = 25'b0000000000000101010011000;
    rom[13401] = 25'b0000000000000101010001011;
    rom[13402] = 25'b0000000000000101001111101;
    rom[13403] = 25'b0000000000000101001110001;
    rom[13404] = 25'b0000000000000101001100011;
    rom[13405] = 25'b0000000000000101001010110;
    rom[13406] = 25'b0000000000000101001001001;
    rom[13407] = 25'b0000000000000101000111011;
    rom[13408] = 25'b0000000000000101000101101;
    rom[13409] = 25'b0000000000000101000100001;
    rom[13410] = 25'b0000000000000101000010011;
    rom[13411] = 25'b0000000000000101000000101;
    rom[13412] = 25'b0000000000000100111111000;
    rom[13413] = 25'b0000000000000100111101010;
    rom[13414] = 25'b0000000000000100111011101;
    rom[13415] = 25'b0000000000000100111010000;
    rom[13416] = 25'b0000000000000100111000010;
    rom[13417] = 25'b0000000000000100110110101;
    rom[13418] = 25'b0000000000000100110100111;
    rom[13419] = 25'b0000000000000100110011001;
    rom[13420] = 25'b0000000000000100110001100;
    rom[13421] = 25'b0000000000000100101111101;
    rom[13422] = 25'b0000000000000100101110000;
    rom[13423] = 25'b0000000000000100101100010;
    rom[13424] = 25'b0000000000000100101010101;
    rom[13425] = 25'b0000000000000100101000111;
    rom[13426] = 25'b0000000000000100100111001;
    rom[13427] = 25'b0000000000000100100101100;
    rom[13428] = 25'b0000000000000100100011101;
    rom[13429] = 25'b0000000000000100100010000;
    rom[13430] = 25'b0000000000000100100000010;
    rom[13431] = 25'b0000000000000100011110100;
    rom[13432] = 25'b0000000000000100011100110;
    rom[13433] = 25'b0000000000000100011011000;
    rom[13434] = 25'b0000000000000100011001011;
    rom[13435] = 25'b0000000000000100010111100;
    rom[13436] = 25'b0000000000000100010101111;
    rom[13437] = 25'b0000000000000100010100001;
    rom[13438] = 25'b0000000000000100010010011;
    rom[13439] = 25'b0000000000000100010000101;
    rom[13440] = 25'b0000000000000100001110111;
    rom[13441] = 25'b0000000000000100001101001;
    rom[13442] = 25'b0000000000000100001011011;
    rom[13443] = 25'b0000000000000100001001101;
    rom[13444] = 25'b0000000000000100000111111;
    rom[13445] = 25'b0000000000000100000110001;
    rom[13446] = 25'b0000000000000100000100011;
    rom[13447] = 25'b0000000000000100000010101;
    rom[13448] = 25'b0000000000000100000000111;
    rom[13449] = 25'b0000000000000011111111010;
    rom[13450] = 25'b0000000000000011111101011;
    rom[13451] = 25'b0000000000000011111011101;
    rom[13452] = 25'b0000000000000011111001111;
    rom[13453] = 25'b0000000000000011111000001;
    rom[13454] = 25'b0000000000000011110110011;
    rom[13455] = 25'b0000000000000011110100101;
    rom[13456] = 25'b0000000000000011110010111;
    rom[13457] = 25'b0000000000000011110001001;
    rom[13458] = 25'b0000000000000011101111011;
    rom[13459] = 25'b0000000000000011101101101;
    rom[13460] = 25'b0000000000000011101011111;
    rom[13461] = 25'b0000000000000011101010001;
    rom[13462] = 25'b0000000000000011101000011;
    rom[13463] = 25'b0000000000000011100110101;
    rom[13464] = 25'b0000000000000011100100111;
    rom[13465] = 25'b0000000000000011100011001;
    rom[13466] = 25'b0000000000000011100001011;
    rom[13467] = 25'b0000000000000011011111101;
    rom[13468] = 25'b0000000000000011011101110;
    rom[13469] = 25'b0000000000000011011100001;
    rom[13470] = 25'b0000000000000011011010010;
    rom[13471] = 25'b0000000000000011011000101;
    rom[13472] = 25'b0000000000000011010110110;
    rom[13473] = 25'b0000000000000011010101001;
    rom[13474] = 25'b0000000000000011010011010;
    rom[13475] = 25'b0000000000000011010001101;
    rom[13476] = 25'b0000000000000011001111110;
    rom[13477] = 25'b0000000000000011001110001;
    rom[13478] = 25'b0000000000000011001100011;
    rom[13479] = 25'b0000000000000011001010101;
    rom[13480] = 25'b0000000000000011001000111;
    rom[13481] = 25'b0000000000000011000111000;
    rom[13482] = 25'b0000000000000011000101011;
    rom[13483] = 25'b0000000000000011000011101;
    rom[13484] = 25'b0000000000000011000001111;
    rom[13485] = 25'b0000000000000011000000001;
    rom[13486] = 25'b0000000000000010111110100;
    rom[13487] = 25'b0000000000000010111100101;
    rom[13488] = 25'b0000000000000010111011000;
    rom[13489] = 25'b0000000000000010111001010;
    rom[13490] = 25'b0000000000000010110111011;
    rom[13491] = 25'b0000000000000010110101110;
    rom[13492] = 25'b0000000000000010110100000;
    rom[13493] = 25'b0000000000000010110010011;
    rom[13494] = 25'b0000000000000010110000101;
    rom[13495] = 25'b0000000000000010101110111;
    rom[13496] = 25'b0000000000000010101101001;
    rom[13497] = 25'b0000000000000010101011011;
    rom[13498] = 25'b0000000000000010101001110;
    rom[13499] = 25'b0000000000000010101000000;
    rom[13500] = 25'b0000000000000010100110011;
    rom[13501] = 25'b0000000000000010100100101;
    rom[13502] = 25'b0000000000000010100010111;
    rom[13503] = 25'b0000000000000010100001010;
    rom[13504] = 25'b0000000000000010011111100;
    rom[13505] = 25'b0000000000000010011101110;
    rom[13506] = 25'b0000000000000010011100001;
    rom[13507] = 25'b0000000000000010011010011;
    rom[13508] = 25'b0000000000000010011000110;
    rom[13509] = 25'b0000000000000010010111000;
    rom[13510] = 25'b0000000000000010010101010;
    rom[13511] = 25'b0000000000000010010011101;
    rom[13512] = 25'b0000000000000010010001111;
    rom[13513] = 25'b0000000000000010010000010;
    rom[13514] = 25'b0000000000000010001110101;
    rom[13515] = 25'b0000000000000010001100111;
    rom[13516] = 25'b0000000000000010001011010;
    rom[13517] = 25'b0000000000000010001001101;
    rom[13518] = 25'b0000000000000010000111111;
    rom[13519] = 25'b0000000000000010000110010;
    rom[13520] = 25'b0000000000000010000100101;
    rom[13521] = 25'b0000000000000010000010111;
    rom[13522] = 25'b0000000000000010000001011;
    rom[13523] = 25'b0000000000000001111111101;
    rom[13524] = 25'b0000000000000001111110000;
    rom[13525] = 25'b0000000000000001111100011;
    rom[13526] = 25'b0000000000000001111010110;
    rom[13527] = 25'b0000000000000001111001000;
    rom[13528] = 25'b0000000000000001110111011;
    rom[13529] = 25'b0000000000000001110101111;
    rom[13530] = 25'b0000000000000001110100001;
    rom[13531] = 25'b0000000000000001110010100;
    rom[13532] = 25'b0000000000000001110001000;
    rom[13533] = 25'b0000000000000001101111011;
    rom[13534] = 25'b0000000000000001101101101;
    rom[13535] = 25'b0000000000000001101100000;
    rom[13536] = 25'b0000000000000001101010100;
    rom[13537] = 25'b0000000000000001101000111;
    rom[13538] = 25'b0000000000000001100111010;
    rom[13539] = 25'b0000000000000001100101101;
    rom[13540] = 25'b0000000000000001100100001;
    rom[13541] = 25'b0000000000000001100010100;
    rom[13542] = 25'b0000000000000001100000111;
    rom[13543] = 25'b0000000000000001011111010;
    rom[13544] = 25'b0000000000000001011101110;
    rom[13545] = 25'b0000000000000001011100010;
    rom[13546] = 25'b0000000000000001011010101;
    rom[13547] = 25'b0000000000000001011001000;
    rom[13548] = 25'b0000000000000001010111100;
    rom[13549] = 25'b0000000000000001010110000;
    rom[13550] = 25'b0000000000000001010100011;
    rom[13551] = 25'b0000000000000001010010111;
    rom[13552] = 25'b0000000000000001010001010;
    rom[13553] = 25'b0000000000000001001111110;
    rom[13554] = 25'b0000000000000001001110001;
    rom[13555] = 25'b0000000000000001001100110;
    rom[13556] = 25'b0000000000000001001011010;
    rom[13557] = 25'b0000000000000001001001101;
    rom[13558] = 25'b0000000000000001001000001;
    rom[13559] = 25'b0000000000000001000110101;
    rom[13560] = 25'b0000000000000001000101001;
    rom[13561] = 25'b0000000000000001000011100;
    rom[13562] = 25'b0000000000000001000010001;
    rom[13563] = 25'b0000000000000001000000101;
    rom[13564] = 25'b0000000000000000111111001;
    rom[13565] = 25'b0000000000000000111101101;
    rom[13566] = 25'b0000000000000000111100001;
    rom[13567] = 25'b0000000000000000111010101;
    rom[13568] = 25'b0000000000000000111001010;
    rom[13569] = 25'b0000000000000000110111110;
    rom[13570] = 25'b0000000000000000110110010;
    rom[13571] = 25'b0000000000000000110100110;
    rom[13572] = 25'b0000000000000000110011011;
    rom[13573] = 25'b0000000000000000110001111;
    rom[13574] = 25'b0000000000000000110000011;
    rom[13575] = 25'b0000000000000000101111000;
    rom[13576] = 25'b0000000000000000101101100;
    rom[13577] = 25'b0000000000000000101100001;
    rom[13578] = 25'b0000000000000000101010101;
    rom[13579] = 25'b0000000000000000101001010;
    rom[13580] = 25'b0000000000000000100111111;
    rom[13581] = 25'b0000000000000000100110100;
    rom[13582] = 25'b0000000000000000100101000;
    rom[13583] = 25'b0000000000000000100011101;
    rom[13584] = 25'b0000000000000000100010010;
    rom[13585] = 25'b0000000000000000100000111;
    rom[13586] = 25'b0000000000000000011111100;
    rom[13587] = 25'b0000000000000000011110001;
    rom[13588] = 25'b0000000000000000011100110;
    rom[13589] = 25'b0000000000000000011011011;
    rom[13590] = 25'b0000000000000000011010000;
    rom[13591] = 25'b0000000000000000011000110;
    rom[13592] = 25'b0000000000000000010111011;
    rom[13593] = 25'b0000000000000000010110000;
    rom[13594] = 25'b0000000000000000010100101;
    rom[13595] = 25'b0000000000000000010011010;
    rom[13596] = 25'b0000000000000000010001111;
    rom[13597] = 25'b0000000000000000010000101;
    rom[13598] = 25'b0000000000000000001111011;
    rom[13599] = 25'b0000000000000000001110000;
    rom[13600] = 25'b0000000000000000001100110;
    rom[13601] = 25'b0000000000000000001011011;
    rom[13602] = 25'b0000000000000000001010000;
    rom[13603] = 25'b0000000000000000001000110;
    rom[13604] = 25'b0000000000000000000111100;
    rom[13605] = 25'b0000000000000000000110010;
    rom[13606] = 25'b0000000000000000000100111;
    rom[13607] = 25'b0000000000000000000011101;
    rom[13608] = 25'b0000000000000000000010011;
    rom[13609] = 25'b0000000000000000000001001;
    rom[13610] = 25'b0000000000000000000000000;
    rom[13611] = 25'b1111111111111111111110110;
    rom[13612] = 25'b1111111111111111111101100;
    rom[13613] = 25'b1111111111111111111100010;
    rom[13614] = 25'b1111111111111111111011000;
    rom[13615] = 25'b1111111111111111111001110;
    rom[13616] = 25'b1111111111111111111000101;
    rom[13617] = 25'b1111111111111111110111011;
    rom[13618] = 25'b1111111111111111110110001;
    rom[13619] = 25'b1111111111111111110101000;
    rom[13620] = 25'b1111111111111111110011110;
    rom[13621] = 25'b1111111111111111110010100;
    rom[13622] = 25'b1111111111111111110001011;
    rom[13623] = 25'b1111111111111111110000010;
    rom[13624] = 25'b1111111111111111101111000;
    rom[13625] = 25'b1111111111111111101101111;
    rom[13626] = 25'b1111111111111111101100110;
    rom[13627] = 25'b1111111111111111101011100;
    rom[13628] = 25'b1111111111111111101010011;
    rom[13629] = 25'b1111111111111111101001001;
    rom[13630] = 25'b1111111111111111101000001;
    rom[13631] = 25'b1111111111111111100111000;
    rom[13632] = 25'b1111111111111111100101110;
    rom[13633] = 25'b1111111111111111100100110;
    rom[13634] = 25'b1111111111111111100011100;
    rom[13635] = 25'b1111111111111111100010100;
    rom[13636] = 25'b1111111111111111100001011;
    rom[13637] = 25'b1111111111111111100000010;
    rom[13638] = 25'b1111111111111111011111010;
    rom[13639] = 25'b1111111111111111011110001;
    rom[13640] = 25'b1111111111111111011101000;
    rom[13641] = 25'b1111111111111111011011111;
    rom[13642] = 25'b1111111111111111011010111;
    rom[13643] = 25'b1111111111111111011001110;
    rom[13644] = 25'b1111111111111111011000110;
    rom[13645] = 25'b1111111111111111010111101;
    rom[13646] = 25'b1111111111111111010110110;
    rom[13647] = 25'b1111111111111111010101101;
    rom[13648] = 25'b1111111111111111010100100;
    rom[13649] = 25'b1111111111111111010011100;
    rom[13650] = 25'b1111111111111111010010100;
    rom[13651] = 25'b1111111111111111010001100;
    rom[13652] = 25'b1111111111111111010000100;
    rom[13653] = 25'b1111111111111111001111100;
    rom[13654] = 25'b1111111111111111001110100;
    rom[13655] = 25'b1111111111111111001101100;
    rom[13656] = 25'b1111111111111111001100100;
    rom[13657] = 25'b1111111111111111001011100;
    rom[13658] = 25'b1111111111111111001010101;
    rom[13659] = 25'b1111111111111111001001101;
    rom[13660] = 25'b1111111111111111001000101;
    rom[13661] = 25'b1111111111111111000111110;
    rom[13662] = 25'b1111111111111111000110110;
    rom[13663] = 25'b1111111111111111000101110;
    rom[13664] = 25'b1111111111111111000100111;
    rom[13665] = 25'b1111111111111111000100000;
    rom[13666] = 25'b1111111111111111000011000;
    rom[13667] = 25'b1111111111111111000010001;
    rom[13668] = 25'b1111111111111111000001010;
    rom[13669] = 25'b1111111111111111000000010;
    rom[13670] = 25'b1111111111111110111111011;
    rom[13671] = 25'b1111111111111110111110100;
    rom[13672] = 25'b1111111111111110111101101;
    rom[13673] = 25'b1111111111111110111100110;
    rom[13674] = 25'b1111111111111110111011111;
    rom[13675] = 25'b1111111111111110111011000;
    rom[13676] = 25'b1111111111111110111010001;
    rom[13677] = 25'b1111111111111110111001010;
    rom[13678] = 25'b1111111111111110111000011;
    rom[13679] = 25'b1111111111111110110111101;
    rom[13680] = 25'b1111111111111110110110110;
    rom[13681] = 25'b1111111111111110110110000;
    rom[13682] = 25'b1111111111111110110101001;
    rom[13683] = 25'b1111111111111110110100010;
    rom[13684] = 25'b1111111111111110110011100;
    rom[13685] = 25'b1111111111111110110010101;
    rom[13686] = 25'b1111111111111110110001111;
    rom[13687] = 25'b1111111111111110110001000;
    rom[13688] = 25'b1111111111111110110000010;
    rom[13689] = 25'b1111111111111110101111100;
    rom[13690] = 25'b1111111111111110101110110;
    rom[13691] = 25'b1111111111111110101110000;
    rom[13692] = 25'b1111111111111110101101010;
    rom[13693] = 25'b1111111111111110101100100;
    rom[13694] = 25'b1111111111111110101011110;
    rom[13695] = 25'b1111111111111110101011000;
    rom[13696] = 25'b1111111111111110101010010;
    rom[13697] = 25'b1111111111111110101001100;
    rom[13698] = 25'b1111111111111110101000110;
    rom[13699] = 25'b1111111111111110101000000;
    rom[13700] = 25'b1111111111111110100111011;
    rom[13701] = 25'b1111111111111110100110101;
    rom[13702] = 25'b1111111111111110100101111;
    rom[13703] = 25'b1111111111111110100101010;
    rom[13704] = 25'b1111111111111110100100100;
    rom[13705] = 25'b1111111111111110100011111;
    rom[13706] = 25'b1111111111111110100011001;
    rom[13707] = 25'b1111111111111110100010100;
    rom[13708] = 25'b1111111111111110100001111;
    rom[13709] = 25'b1111111111111110100001010;
    rom[13710] = 25'b1111111111111110100000101;
    rom[13711] = 25'b1111111111111110100000000;
    rom[13712] = 25'b1111111111111110011111010;
    rom[13713] = 25'b1111111111111110011110101;
    rom[13714] = 25'b1111111111111110011110000;
    rom[13715] = 25'b1111111111111110011101011;
    rom[13716] = 25'b1111111111111110011100110;
    rom[13717] = 25'b1111111111111110011100001;
    rom[13718] = 25'b1111111111111110011011101;
    rom[13719] = 25'b1111111111111110011011000;
    rom[13720] = 25'b1111111111111110011010010;
    rom[13721] = 25'b1111111111111110011001110;
    rom[13722] = 25'b1111111111111110011001001;
    rom[13723] = 25'b1111111111111110011000101;
    rom[13724] = 25'b1111111111111110011000001;
    rom[13725] = 25'b1111111111111110010111011;
    rom[13726] = 25'b1111111111111110010110111;
    rom[13727] = 25'b1111111111111110010110011;
    rom[13728] = 25'b1111111111111110010101111;
    rom[13729] = 25'b1111111111111110010101010;
    rom[13730] = 25'b1111111111111110010100110;
    rom[13731] = 25'b1111111111111110010100010;
    rom[13732] = 25'b1111111111111110010011110;
    rom[13733] = 25'b1111111111111110010011001;
    rom[13734] = 25'b1111111111111110010010101;
    rom[13735] = 25'b1111111111111110010010010;
    rom[13736] = 25'b1111111111111110010001110;
    rom[13737] = 25'b1111111111111110010001001;
    rom[13738] = 25'b1111111111111110010000110;
    rom[13739] = 25'b1111111111111110010000010;
    rom[13740] = 25'b1111111111111110001111110;
    rom[13741] = 25'b1111111111111110001111011;
    rom[13742] = 25'b1111111111111110001110111;
    rom[13743] = 25'b1111111111111110001110011;
    rom[13744] = 25'b1111111111111110001110000;
    rom[13745] = 25'b1111111111111110001101100;
    rom[13746] = 25'b1111111111111110001101000;
    rom[13747] = 25'b1111111111111110001100101;
    rom[13748] = 25'b1111111111111110001100001;
    rom[13749] = 25'b1111111111111110001011110;
    rom[13750] = 25'b1111111111111110001011011;
    rom[13751] = 25'b1111111111111110001011000;
    rom[13752] = 25'b1111111111111110001010101;
    rom[13753] = 25'b1111111111111110001010001;
    rom[13754] = 25'b1111111111111110001001110;
    rom[13755] = 25'b1111111111111110001001011;
    rom[13756] = 25'b1111111111111110001001000;
    rom[13757] = 25'b1111111111111110001000101;
    rom[13758] = 25'b1111111111111110001000010;
    rom[13759] = 25'b1111111111111110000111111;
    rom[13760] = 25'b1111111111111110000111100;
    rom[13761] = 25'b1111111111111110000111001;
    rom[13762] = 25'b1111111111111110000110111;
    rom[13763] = 25'b1111111111111110000110100;
    rom[13764] = 25'b1111111111111110000110001;
    rom[13765] = 25'b1111111111111110000101110;
    rom[13766] = 25'b1111111111111110000101100;
    rom[13767] = 25'b1111111111111110000101001;
    rom[13768] = 25'b1111111111111110000100111;
    rom[13769] = 25'b1111111111111110000100100;
    rom[13770] = 25'b1111111111111110000100010;
    rom[13771] = 25'b1111111111111110000100000;
    rom[13772] = 25'b1111111111111110000011101;
    rom[13773] = 25'b1111111111111110000011011;
    rom[13774] = 25'b1111111111111110000011001;
    rom[13775] = 25'b1111111111111110000010110;
    rom[13776] = 25'b1111111111111110000010100;
    rom[13777] = 25'b1111111111111110000010010;
    rom[13778] = 25'b1111111111111110000010000;
    rom[13779] = 25'b1111111111111110000001110;
    rom[13780] = 25'b1111111111111110000001100;
    rom[13781] = 25'b1111111111111110000001010;
    rom[13782] = 25'b1111111111111110000001000;
    rom[13783] = 25'b1111111111111110000000110;
    rom[13784] = 25'b1111111111111110000000101;
    rom[13785] = 25'b1111111111111110000000011;
    rom[13786] = 25'b1111111111111110000000001;
    rom[13787] = 25'b1111111111111110000000000;
    rom[13788] = 25'b1111111111111101111111110;
    rom[13789] = 25'b1111111111111101111111100;
    rom[13790] = 25'b1111111111111101111111010;
    rom[13791] = 25'b1111111111111101111111001;
    rom[13792] = 25'b1111111111111101111110111;
    rom[13793] = 25'b1111111111111101111110110;
    rom[13794] = 25'b1111111111111101111110100;
    rom[13795] = 25'b1111111111111101111110011;
    rom[13796] = 25'b1111111111111101111110010;
    rom[13797] = 25'b1111111111111101111110000;
    rom[13798] = 25'b1111111111111101111101111;
    rom[13799] = 25'b1111111111111101111101110;
    rom[13800] = 25'b1111111111111101111101101;
    rom[13801] = 25'b1111111111111101111101100;
    rom[13802] = 25'b1111111111111101111101010;
    rom[13803] = 25'b1111111111111101111101001;
    rom[13804] = 25'b1111111111111101111101001;
    rom[13805] = 25'b1111111111111101111101000;
    rom[13806] = 25'b1111111111111101111100111;
    rom[13807] = 25'b1111111111111101111100110;
    rom[13808] = 25'b1111111111111101111100101;
    rom[13809] = 25'b1111111111111101111100100;
    rom[13810] = 25'b1111111111111101111100011;
    rom[13811] = 25'b1111111111111101111100011;
    rom[13812] = 25'b1111111111111101111100010;
    rom[13813] = 25'b1111111111111101111100001;
    rom[13814] = 25'b1111111111111101111100001;
    rom[13815] = 25'b1111111111111101111100000;
    rom[13816] = 25'b1111111111111101111011111;
    rom[13817] = 25'b1111111111111101111011111;
    rom[13818] = 25'b1111111111111101111011110;
    rom[13819] = 25'b1111111111111101111011101;
    rom[13820] = 25'b1111111111111101111011101;
    rom[13821] = 25'b1111111111111101111011101;
    rom[13822] = 25'b1111111111111101111011101;
    rom[13823] = 25'b1111111111111101111011101;
    rom[13824] = 25'b1111111111111101111011101;
    rom[13825] = 25'b1111111111111101111011100;
    rom[13826] = 25'b1111111111111101111011100;
    rom[13827] = 25'b1111111111111101111011100;
    rom[13828] = 25'b1111111111111101111011100;
    rom[13829] = 25'b1111111111111101111011100;
    rom[13830] = 25'b1111111111111101111011100;
    rom[13831] = 25'b1111111111111101111011100;
    rom[13832] = 25'b1111111111111101111011100;
    rom[13833] = 25'b1111111111111101111011100;
    rom[13834] = 25'b1111111111111101111011100;
    rom[13835] = 25'b1111111111111101111011100;
    rom[13836] = 25'b1111111111111101111011100;
    rom[13837] = 25'b1111111111111101111011100;
    rom[13838] = 25'b1111111111111101111011101;
    rom[13839] = 25'b1111111111111101111011101;
    rom[13840] = 25'b1111111111111101111011101;
    rom[13841] = 25'b1111111111111101111011101;
    rom[13842] = 25'b1111111111111101111011101;
    rom[13843] = 25'b1111111111111101111011101;
    rom[13844] = 25'b1111111111111101111011110;
    rom[13845] = 25'b1111111111111101111011111;
    rom[13846] = 25'b1111111111111101111011111;
    rom[13847] = 25'b1111111111111101111100000;
    rom[13848] = 25'b1111111111111101111100000;
    rom[13849] = 25'b1111111111111101111100001;
    rom[13850] = 25'b1111111111111101111100010;
    rom[13851] = 25'b1111111111111101111100011;
    rom[13852] = 25'b1111111111111101111100011;
    rom[13853] = 25'b1111111111111101111100011;
    rom[13854] = 25'b1111111111111101111100100;
    rom[13855] = 25'b1111111111111101111100101;
    rom[13856] = 25'b1111111111111101111100110;
    rom[13857] = 25'b1111111111111101111100111;
    rom[13858] = 25'b1111111111111101111101000;
    rom[13859] = 25'b1111111111111101111101001;
    rom[13860] = 25'b1111111111111101111101001;
    rom[13861] = 25'b1111111111111101111101010;
    rom[13862] = 25'b1111111111111101111101011;
    rom[13863] = 25'b1111111111111101111101101;
    rom[13864] = 25'b1111111111111101111101110;
    rom[13865] = 25'b1111111111111101111101110;
    rom[13866] = 25'b1111111111111101111101111;
    rom[13867] = 25'b1111111111111101111110001;
    rom[13868] = 25'b1111111111111101111110010;
    rom[13869] = 25'b1111111111111101111110100;
    rom[13870] = 25'b1111111111111101111110100;
    rom[13871] = 25'b1111111111111101111110101;
    rom[13872] = 25'b1111111111111101111110111;
    rom[13873] = 25'b1111111111111101111111001;
    rom[13874] = 25'b1111111111111101111111010;
    rom[13875] = 25'b1111111111111101111111011;
    rom[13876] = 25'b1111111111111101111111100;
    rom[13877] = 25'b1111111111111101111111110;
    rom[13878] = 25'b1111111111111110000000000;
    rom[13879] = 25'b1111111111111110000000000;
    rom[13880] = 25'b1111111111111110000000010;
    rom[13881] = 25'b1111111111111110000000100;
    rom[13882] = 25'b1111111111111110000000101;
    rom[13883] = 25'b1111111111111110000000111;
    rom[13884] = 25'b1111111111111110000001001;
    rom[13885] = 25'b1111111111111110000001011;
    rom[13886] = 25'b1111111111111110000001011;
    rom[13887] = 25'b1111111111111110000001101;
    rom[13888] = 25'b1111111111111110000001111;
    rom[13889] = 25'b1111111111111110000010001;
    rom[13890] = 25'b1111111111111110000010011;
    rom[13891] = 25'b1111111111111110000010101;
    rom[13892] = 25'b1111111111111110000010110;
    rom[13893] = 25'b1111111111111110000011000;
    rom[13894] = 25'b1111111111111110000011010;
    rom[13895] = 25'b1111111111111110000011100;
    rom[13896] = 25'b1111111111111110000011110;
    rom[13897] = 25'b1111111111111110000100000;
    rom[13898] = 25'b1111111111111110000100010;
    rom[13899] = 25'b1111111111111110000100100;
    rom[13900] = 25'b1111111111111110000100110;
    rom[13901] = 25'b1111111111111110000100111;
    rom[13902] = 25'b1111111111111110000101010;
    rom[13903] = 25'b1111111111111110000101100;
    rom[13904] = 25'b1111111111111110000101110;
    rom[13905] = 25'b1111111111111110000110000;
    rom[13906] = 25'b1111111111111110000110011;
    rom[13907] = 25'b1111111111111110000110100;
    rom[13908] = 25'b1111111111111110000110111;
    rom[13909] = 25'b1111111111111110000111000;
    rom[13910] = 25'b1111111111111110000111011;
    rom[13911] = 25'b1111111111111110000111110;
    rom[13912] = 25'b1111111111111110000111111;
    rom[13913] = 25'b1111111111111110001000010;
    rom[13914] = 25'b1111111111111110001000100;
    rom[13915] = 25'b1111111111111110001000110;
    rom[13916] = 25'b1111111111111110001001001;
    rom[13917] = 25'b1111111111111110001001011;
    rom[13918] = 25'b1111111111111110001001110;
    rom[13919] = 25'b1111111111111110001010000;
    rom[13920] = 25'b1111111111111110001010010;
    rom[13921] = 25'b1111111111111110001010101;
    rom[13922] = 25'b1111111111111110001010111;
    rom[13923] = 25'b1111111111111110001011010;
    rom[13924] = 25'b1111111111111110001011100;
    rom[13925] = 25'b1111111111111110001011111;
    rom[13926] = 25'b1111111111111110001100001;
    rom[13927] = 25'b1111111111111110001100100;
    rom[13928] = 25'b1111111111111110001100110;
    rom[13929] = 25'b1111111111111110001101001;
    rom[13930] = 25'b1111111111111110001101100;
    rom[13931] = 25'b1111111111111110001101110;
    rom[13932] = 25'b1111111111111110001110001;
    rom[13933] = 25'b1111111111111110001110100;
    rom[13934] = 25'b1111111111111110001110111;
    rom[13935] = 25'b1111111111111110001111001;
    rom[13936] = 25'b1111111111111110001111100;
    rom[13937] = 25'b1111111111111110001111110;
    rom[13938] = 25'b1111111111111110010000010;
    rom[13939] = 25'b1111111111111110010000100;
    rom[13940] = 25'b1111111111111110010000111;
    rom[13941] = 25'b1111111111111110010001010;
    rom[13942] = 25'b1111111111111110010001101;
    rom[13943] = 25'b1111111111111110010001111;
    rom[13944] = 25'b1111111111111110010010011;
    rom[13945] = 25'b1111111111111110010010101;
    rom[13946] = 25'b1111111111111110010011000;
    rom[13947] = 25'b1111111111111110010011011;
    rom[13948] = 25'b1111111111111110010011110;
    rom[13949] = 25'b1111111111111110010100001;
    rom[13950] = 25'b1111111111111110010100100;
    rom[13951] = 25'b1111111111111110010100111;
    rom[13952] = 25'b1111111111111110010101010;
    rom[13953] = 25'b1111111111111110010101101;
    rom[13954] = 25'b1111111111111110010110000;
    rom[13955] = 25'b1111111111111110010110011;
    rom[13956] = 25'b1111111111111110010110110;
    rom[13957] = 25'b1111111111111110010111001;
    rom[13958] = 25'b1111111111111110010111011;
    rom[13959] = 25'b1111111111111110010111111;
    rom[13960] = 25'b1111111111111110011000010;
    rom[13961] = 25'b1111111111111110011000101;
    rom[13962] = 25'b1111111111111110011001000;
    rom[13963] = 25'b1111111111111110011001100;
    rom[13964] = 25'b1111111111111110011001110;
    rom[13965] = 25'b1111111111111110011010010;
    rom[13966] = 25'b1111111111111110011010101;
    rom[13967] = 25'b1111111111111110011011000;
    rom[13968] = 25'b1111111111111110011011011;
    rom[13969] = 25'b1111111111111110011011110;
    rom[13970] = 25'b1111111111111110011100010;
    rom[13971] = 25'b1111111111111110011100101;
    rom[13972] = 25'b1111111111111110011101000;
    rom[13973] = 25'b1111111111111110011101011;
    rom[13974] = 25'b1111111111111110011101110;
    rom[13975] = 25'b1111111111111110011110010;
    rom[13976] = 25'b1111111111111110011110101;
    rom[13977] = 25'b1111111111111110011111001;
    rom[13978] = 25'b1111111111111110011111011;
    rom[13979] = 25'b1111111111111110011111111;
    rom[13980] = 25'b1111111111111110100000010;
    rom[13981] = 25'b1111111111111110100000101;
    rom[13982] = 25'b1111111111111110100001001;
    rom[13983] = 25'b1111111111111110100001100;
    rom[13984] = 25'b1111111111111110100010000;
    rom[13985] = 25'b1111111111111110100010011;
    rom[13986] = 25'b1111111111111110100010110;
    rom[13987] = 25'b1111111111111110100011010;
    rom[13988] = 25'b1111111111111110100011101;
    rom[13989] = 25'b1111111111111110100100001;
    rom[13990] = 25'b1111111111111110100100100;
    rom[13991] = 25'b1111111111111110100100111;
    rom[13992] = 25'b1111111111111110100101011;
    rom[13993] = 25'b1111111111111110100101110;
    rom[13994] = 25'b1111111111111110100110010;
    rom[13995] = 25'b1111111111111110100110101;
    rom[13996] = 25'b1111111111111110100111000;
    rom[13997] = 25'b1111111111111110100111100;
    rom[13998] = 25'b1111111111111110100111111;
    rom[13999] = 25'b1111111111111110101000011;
    rom[14000] = 25'b1111111111111110101000110;
    rom[14001] = 25'b1111111111111110101001001;
    rom[14002] = 25'b1111111111111110101001101;
    rom[14003] = 25'b1111111111111110101010001;
    rom[14004] = 25'b1111111111111110101010101;
    rom[14005] = 25'b1111111111111110101011000;
    rom[14006] = 25'b1111111111111110101011011;
    rom[14007] = 25'b1111111111111110101011111;
    rom[14008] = 25'b1111111111111110101100010;
    rom[14009] = 25'b1111111111111110101100110;
    rom[14010] = 25'b1111111111111110101101010;
    rom[14011] = 25'b1111111111111110101101101;
    rom[14012] = 25'b1111111111111110101110001;
    rom[14013] = 25'b1111111111111110101110100;
    rom[14014] = 25'b1111111111111110101110111;
    rom[14015] = 25'b1111111111111110101111011;
    rom[14016] = 25'b1111111111111110101111111;
    rom[14017] = 25'b1111111111111110110000010;
    rom[14018] = 25'b1111111111111110110000110;
    rom[14019] = 25'b1111111111111110110001001;
    rom[14020] = 25'b1111111111111110110001110;
    rom[14021] = 25'b1111111111111110110010001;
    rom[14022] = 25'b1111111111111110110010100;
    rom[14023] = 25'b1111111111111110110011000;
    rom[14024] = 25'b1111111111111110110011011;
    rom[14025] = 25'b1111111111111110110011111;
    rom[14026] = 25'b1111111111111110110100011;
    rom[14027] = 25'b1111111111111110110100110;
    rom[14028] = 25'b1111111111111110110101010;
    rom[14029] = 25'b1111111111111110110101110;
    rom[14030] = 25'b1111111111111110110110001;
    rom[14031] = 25'b1111111111111110110110101;
    rom[14032] = 25'b1111111111111110110111000;
    rom[14033] = 25'b1111111111111110110111100;
    rom[14034] = 25'b1111111111111110111000000;
    rom[14035] = 25'b1111111111111110111000011;
    rom[14036] = 25'b1111111111111110111000111;
    rom[14037] = 25'b1111111111111110111001011;
    rom[14038] = 25'b1111111111111110111001110;
    rom[14039] = 25'b1111111111111110111010010;
    rom[14040] = 25'b1111111111111110111010110;
    rom[14041] = 25'b1111111111111110111011001;
    rom[14042] = 25'b1111111111111110111011101;
    rom[14043] = 25'b1111111111111110111100000;
    rom[14044] = 25'b1111111111111110111100100;
    rom[14045] = 25'b1111111111111110111101000;
    rom[14046] = 25'b1111111111111110111101011;
    rom[14047] = 25'b1111111111111110111101110;
    rom[14048] = 25'b1111111111111110111110011;
    rom[14049] = 25'b1111111111111110111110110;
    rom[14050] = 25'b1111111111111110111111010;
    rom[14051] = 25'b1111111111111110111111110;
    rom[14052] = 25'b1111111111111111000000001;
    rom[14053] = 25'b1111111111111111000000101;
    rom[14054] = 25'b1111111111111111000001000;
    rom[14055] = 25'b1111111111111111000001100;
    rom[14056] = 25'b1111111111111111000010000;
    rom[14057] = 25'b1111111111111111000010011;
    rom[14058] = 25'b1111111111111111000010110;
    rom[14059] = 25'b1111111111111111000011011;
    rom[14060] = 25'b1111111111111111000011110;
    rom[14061] = 25'b1111111111111111000100010;
    rom[14062] = 25'b1111111111111111000100110;
    rom[14063] = 25'b1111111111111111000101001;
    rom[14064] = 25'b1111111111111111000101101;
    rom[14065] = 25'b1111111111111111000110000;
    rom[14066] = 25'b1111111111111111000110100;
    rom[14067] = 25'b1111111111111111000111000;
    rom[14068] = 25'b1111111111111111000111011;
    rom[14069] = 25'b1111111111111111000111110;
    rom[14070] = 25'b1111111111111111001000011;
    rom[14071] = 25'b1111111111111111001000110;
    rom[14072] = 25'b1111111111111111001001001;
    rom[14073] = 25'b1111111111111111001001101;
    rom[14074] = 25'b1111111111111111001010001;
    rom[14075] = 25'b1111111111111111001010101;
    rom[14076] = 25'b1111111111111111001011000;
    rom[14077] = 25'b1111111111111111001011011;
    rom[14078] = 25'b1111111111111111001011111;
    rom[14079] = 25'b1111111111111111001100011;
    rom[14080] = 25'b1111111111111111001100110;
    rom[14081] = 25'b1111111111111111001101010;
    rom[14082] = 25'b1111111111111111001101101;
    rom[14083] = 25'b1111111111111111001110001;
    rom[14084] = 25'b1111111111111111001110101;
    rom[14085] = 25'b1111111111111111001111000;
    rom[14086] = 25'b1111111111111111001111100;
    rom[14087] = 25'b1111111111111111001111111;
    rom[14088] = 25'b1111111111111111010000010;
    rom[14089] = 25'b1111111111111111010000111;
    rom[14090] = 25'b1111111111111111010001010;
    rom[14091] = 25'b1111111111111111010001110;
    rom[14092] = 25'b1111111111111111010010001;
    rom[14093] = 25'b1111111111111111010010100;
    rom[14094] = 25'b1111111111111111010011000;
    rom[14095] = 25'b1111111111111111010011100;
    rom[14096] = 25'b1111111111111111010011111;
    rom[14097] = 25'b1111111111111111010100011;
    rom[14098] = 25'b1111111111111111010100110;
    rom[14099] = 25'b1111111111111111010101010;
    rom[14100] = 25'b1111111111111111010101101;
    rom[14101] = 25'b1111111111111111010110000;
    rom[14102] = 25'b1111111111111111010110100;
    rom[14103] = 25'b1111111111111111010110111;
    rom[14104] = 25'b1111111111111111010111011;
    rom[14105] = 25'b1111111111111111010111111;
    rom[14106] = 25'b1111111111111111011000010;
    rom[14107] = 25'b1111111111111111011000110;
    rom[14108] = 25'b1111111111111111011001001;
    rom[14109] = 25'b1111111111111111011001100;
    rom[14110] = 25'b1111111111111111011010000;
    rom[14111] = 25'b1111111111111111011010011;
    rom[14112] = 25'b1111111111111111011010111;
    rom[14113] = 25'b1111111111111111011011010;
    rom[14114] = 25'b1111111111111111011011101;
    rom[14115] = 25'b1111111111111111011100001;
    rom[14116] = 25'b1111111111111111011100100;
    rom[14117] = 25'b1111111111111111011101000;
    rom[14118] = 25'b1111111111111111011101011;
    rom[14119] = 25'b1111111111111111011101110;
    rom[14120] = 25'b1111111111111111011110010;
    rom[14121] = 25'b1111111111111111011110101;
    rom[14122] = 25'b1111111111111111011111001;
    rom[14123] = 25'b1111111111111111011111100;
    rom[14124] = 25'b1111111111111111100000000;
    rom[14125] = 25'b1111111111111111100000010;
    rom[14126] = 25'b1111111111111111100000101;
    rom[14127] = 25'b1111111111111111100001001;
    rom[14128] = 25'b1111111111111111100001100;
    rom[14129] = 25'b1111111111111111100010000;
    rom[14130] = 25'b1111111111111111100010011;
    rom[14131] = 25'b1111111111111111100010110;
    rom[14132] = 25'b1111111111111111100011010;
    rom[14133] = 25'b1111111111111111100011100;
    rom[14134] = 25'b1111111111111111100100000;
    rom[14135] = 25'b1111111111111111100100011;
    rom[14136] = 25'b1111111111111111100100111;
    rom[14137] = 25'b1111111111111111100101010;
    rom[14138] = 25'b1111111111111111100101101;
    rom[14139] = 25'b1111111111111111100110000;
    rom[14140] = 25'b1111111111111111100110011;
    rom[14141] = 25'b1111111111111111100110111;
    rom[14142] = 25'b1111111111111111100111010;
    rom[14143] = 25'b1111111111111111100111101;
    rom[14144] = 25'b1111111111111111101000000;
    rom[14145] = 25'b1111111111111111101000100;
    rom[14146] = 25'b1111111111111111101000110;
    rom[14147] = 25'b1111111111111111101001001;
    rom[14148] = 25'b1111111111111111101001101;
    rom[14149] = 25'b1111111111111111101010000;
    rom[14150] = 25'b1111111111111111101010011;
    rom[14151] = 25'b1111111111111111101010110;
    rom[14152] = 25'b1111111111111111101011001;
    rom[14153] = 25'b1111111111111111101011100;
    rom[14154] = 25'b1111111111111111101100000;
    rom[14155] = 25'b1111111111111111101100010;
    rom[14156] = 25'b1111111111111111101100110;
    rom[14157] = 25'b1111111111111111101101001;
    rom[14158] = 25'b1111111111111111101101100;
    rom[14159] = 25'b1111111111111111101101111;
    rom[14160] = 25'b1111111111111111101110001;
    rom[14161] = 25'b1111111111111111101110101;
    rom[14162] = 25'b1111111111111111101110111;
    rom[14163] = 25'b1111111111111111101111011;
    rom[14164] = 25'b1111111111111111101111101;
    rom[14165] = 25'b1111111111111111110000001;
    rom[14166] = 25'b1111111111111111110000011;
    rom[14167] = 25'b1111111111111111110000111;
    rom[14168] = 25'b1111111111111111110001001;
    rom[14169] = 25'b1111111111111111110001101;
    rom[14170] = 25'b1111111111111111110001111;
    rom[14171] = 25'b1111111111111111110010011;
    rom[14172] = 25'b1111111111111111110010101;
    rom[14173] = 25'b1111111111111111110011000;
    rom[14174] = 25'b1111111111111111110011011;
    rom[14175] = 25'b1111111111111111110011110;
    rom[14176] = 25'b1111111111111111110100000;
    rom[14177] = 25'b1111111111111111110100100;
    rom[14178] = 25'b1111111111111111110100110;
    rom[14179] = 25'b1111111111111111110101001;
    rom[14180] = 25'b1111111111111111110101100;
    rom[14181] = 25'b1111111111111111110101111;
    rom[14182] = 25'b1111111111111111110110001;
    rom[14183] = 25'b1111111111111111110110101;
    rom[14184] = 25'b1111111111111111110110111;
    rom[14185] = 25'b1111111111111111110111010;
    rom[14186] = 25'b1111111111111111110111100;
    rom[14187] = 25'b1111111111111111111000000;
    rom[14188] = 25'b1111111111111111111000010;
    rom[14189] = 25'b1111111111111111111000101;
    rom[14190] = 25'b1111111111111111111000111;
    rom[14191] = 25'b1111111111111111111001010;
    rom[14192] = 25'b1111111111111111111001100;
    rom[14193] = 25'b1111111111111111111010000;
    rom[14194] = 25'b1111111111111111111010010;
    rom[14195] = 25'b1111111111111111111010101;
    rom[14196] = 25'b1111111111111111111011000;
    rom[14197] = 25'b1111111111111111111011010;
    rom[14198] = 25'b1111111111111111111011101;
    rom[14199] = 25'b1111111111111111111011111;
    rom[14200] = 25'b1111111111111111111100010;
    rom[14201] = 25'b1111111111111111111100100;
    rom[14202] = 25'b1111111111111111111100111;
    rom[14203] = 25'b1111111111111111111101001;
    rom[14204] = 25'b1111111111111111111101100;
    rom[14205] = 25'b1111111111111111111101110;
    rom[14206] = 25'b1111111111111111111110001;
    rom[14207] = 25'b1111111111111111111110100;
    rom[14208] = 25'b1111111111111111111110110;
    rom[14209] = 25'b1111111111111111111111001;
    rom[14210] = 25'b1111111111111111111111011;
    rom[14211] = 25'b1111111111111111111111110;
    rom[14212] = 25'b0000000000000000000000000;
    rom[14213] = 25'b0000000000000000000000001;
    rom[14214] = 25'b0000000000000000000000100;
    rom[14215] = 25'b0000000000000000000000110;
    rom[14216] = 25'b0000000000000000000001001;
    rom[14217] = 25'b0000000000000000000001011;
    rom[14218] = 25'b0000000000000000000001110;
    rom[14219] = 25'b0000000000000000000010000;
    rom[14220] = 25'b0000000000000000000010010;
    rom[14221] = 25'b0000000000000000000010101;
    rom[14222] = 25'b0000000000000000000010111;
    rom[14223] = 25'b0000000000000000000011001;
    rom[14224] = 25'b0000000000000000000011100;
    rom[14225] = 25'b0000000000000000000011110;
    rom[14226] = 25'b0000000000000000000100000;
    rom[14227] = 25'b0000000000000000000100010;
    rom[14228] = 25'b0000000000000000000100101;
    rom[14229] = 25'b0000000000000000000100111;
    rom[14230] = 25'b0000000000000000000101001;
    rom[14231] = 25'b0000000000000000000101100;
    rom[14232] = 25'b0000000000000000000101101;
    rom[14233] = 25'b0000000000000000000110000;
    rom[14234] = 25'b0000000000000000000110010;
    rom[14235] = 25'b0000000000000000000110100;
    rom[14236] = 25'b0000000000000000000110110;
    rom[14237] = 25'b0000000000000000000111000;
    rom[14238] = 25'b0000000000000000000111010;
    rom[14239] = 25'b0000000000000000000111101;
    rom[14240] = 25'b0000000000000000000111110;
    rom[14241] = 25'b0000000000000000001000001;
    rom[14242] = 25'b0000000000000000001000011;
    rom[14243] = 25'b0000000000000000001000101;
    rom[14244] = 25'b0000000000000000001000111;
    rom[14245] = 25'b0000000000000000001001001;
    rom[14246] = 25'b0000000000000000001001011;
    rom[14247] = 25'b0000000000000000001001101;
    rom[14248] = 25'b0000000000000000001001111;
    rom[14249] = 25'b0000000000000000001010001;
    rom[14250] = 25'b0000000000000000001010011;
    rom[14251] = 25'b0000000000000000001010101;
    rom[14252] = 25'b0000000000000000001010111;
    rom[14253] = 25'b0000000000000000001011001;
    rom[14254] = 25'b0000000000000000001011011;
    rom[14255] = 25'b0000000000000000001011101;
    rom[14256] = 25'b0000000000000000001011111;
    rom[14257] = 25'b0000000000000000001100000;
    rom[14258] = 25'b0000000000000000001100010;
    rom[14259] = 25'b0000000000000000001100101;
    rom[14260] = 25'b0000000000000000001100110;
    rom[14261] = 25'b0000000000000000001101000;
    rom[14262] = 25'b0000000000000000001101010;
    rom[14263] = 25'b0000000000000000001101100;
    rom[14264] = 25'b0000000000000000001101101;
    rom[14265] = 25'b0000000000000000001101111;
    rom[14266] = 25'b0000000000000000001110001;
    rom[14267] = 25'b0000000000000000001110011;
    rom[14268] = 25'b0000000000000000001110101;
    rom[14269] = 25'b0000000000000000001110111;
    rom[14270] = 25'b0000000000000000001111000;
    rom[14271] = 25'b0000000000000000001111010;
    rom[14272] = 25'b0000000000000000001111100;
    rom[14273] = 25'b0000000000000000001111101;
    rom[14274] = 25'b0000000000000000001111111;
    rom[14275] = 25'b0000000000000000010000001;
    rom[14276] = 25'b0000000000000000010000010;
    rom[14277] = 25'b0000000000000000010000100;
    rom[14278] = 25'b0000000000000000010000101;
    rom[14279] = 25'b0000000000000000010000111;
    rom[14280] = 25'b0000000000000000010001000;
    rom[14281] = 25'b0000000000000000010001010;
    rom[14282] = 25'b0000000000000000010001100;
    rom[14283] = 25'b0000000000000000010001110;
    rom[14284] = 25'b0000000000000000010001111;
    rom[14285] = 25'b0000000000000000010010000;
    rom[14286] = 25'b0000000000000000010010010;
    rom[14287] = 25'b0000000000000000010010011;
    rom[14288] = 25'b0000000000000000010010101;
    rom[14289] = 25'b0000000000000000010010111;
    rom[14290] = 25'b0000000000000000010011000;
    rom[14291] = 25'b0000000000000000010011001;
    rom[14292] = 25'b0000000000000000010011011;
    rom[14293] = 25'b0000000000000000010011100;
    rom[14294] = 25'b0000000000000000010011110;
    rom[14295] = 25'b0000000000000000010011111;
    rom[14296] = 25'b0000000000000000010100000;
    rom[14297] = 25'b0000000000000000010100010;
    rom[14298] = 25'b0000000000000000010100100;
    rom[14299] = 25'b0000000000000000010100100;
    rom[14300] = 25'b0000000000000000010100110;
    rom[14301] = 25'b0000000000000000010100111;
    rom[14302] = 25'b0000000000000000010101001;
    rom[14303] = 25'b0000000000000000010101010;
    rom[14304] = 25'b0000000000000000010101011;
    rom[14305] = 25'b0000000000000000010101101;
    rom[14306] = 25'b0000000000000000010101110;
    rom[14307] = 25'b0000000000000000010110000;
    rom[14308] = 25'b0000000000000000010110000;
    rom[14309] = 25'b0000000000000000010110001;
    rom[14310] = 25'b0000000000000000010110011;
    rom[14311] = 25'b0000000000000000010110100;
    rom[14312] = 25'b0000000000000000010110110;
    rom[14313] = 25'b0000000000000000010110110;
    rom[14314] = 25'b0000000000000000010111000;
    rom[14315] = 25'b0000000000000000010111001;
    rom[14316] = 25'b0000000000000000010111010;
    rom[14317] = 25'b0000000000000000010111011;
    rom[14318] = 25'b0000000000000000010111100;
    rom[14319] = 25'b0000000000000000010111101;
    rom[14320] = 25'b0000000000000000010111111;
    rom[14321] = 25'b0000000000000000011000000;
    rom[14322] = 25'b0000000000000000011000001;
    rom[14323] = 25'b0000000000000000011000001;
    rom[14324] = 25'b0000000000000000011000011;
    rom[14325] = 25'b0000000000000000011000100;
    rom[14326] = 25'b0000000000000000011000101;
    rom[14327] = 25'b0000000000000000011000110;
    rom[14328] = 25'b0000000000000000011000111;
    rom[14329] = 25'b0000000000000000011001000;
    rom[14330] = 25'b0000000000000000011001001;
    rom[14331] = 25'b0000000000000000011001010;
    rom[14332] = 25'b0000000000000000011001011;
    rom[14333] = 25'b0000000000000000011001100;
    rom[14334] = 25'b0000000000000000011001100;
    rom[14335] = 25'b0000000000000000011001101;
    rom[14336] = 25'b0000000000000000011001111;
    rom[14337] = 25'b0000000000000000011010000;
    rom[14338] = 25'b0000000000000000011010001;
    rom[14339] = 25'b0000000000000000011010010;
    rom[14340] = 25'b0000000000000000011010010;
    rom[14341] = 25'b0000000000000000011010011;
    rom[14342] = 25'b0000000000000000011010100;
    rom[14343] = 25'b0000000000000000011010101;
    rom[14344] = 25'b0000000000000000011010110;
    rom[14345] = 25'b0000000000000000011010111;
    rom[14346] = 25'b0000000000000000011011000;
    rom[14347] = 25'b0000000000000000011011000;
    rom[14348] = 25'b0000000000000000011011001;
    rom[14349] = 25'b0000000000000000011011001;
    rom[14350] = 25'b0000000000000000011011010;
    rom[14351] = 25'b0000000000000000011011011;
    rom[14352] = 25'b0000000000000000011011100;
    rom[14353] = 25'b0000000000000000011011101;
    rom[14354] = 25'b0000000000000000011011101;
    rom[14355] = 25'b0000000000000000011011110;
    rom[14356] = 25'b0000000000000000011011110;
    rom[14357] = 25'b0000000000000000011011111;
    rom[14358] = 25'b0000000000000000011100000;
    rom[14359] = 25'b0000000000000000011100001;
    rom[14360] = 25'b0000000000000000011100010;
    rom[14361] = 25'b0000000000000000011100010;
    rom[14362] = 25'b0000000000000000011100011;
    rom[14363] = 25'b0000000000000000011100011;
    rom[14364] = 25'b0000000000000000011100011;
    rom[14365] = 25'b0000000000000000011100100;
    rom[14366] = 25'b0000000000000000011100101;
    rom[14367] = 25'b0000000000000000011100110;
    rom[14368] = 25'b0000000000000000011100110;
    rom[14369] = 25'b0000000000000000011100111;
    rom[14370] = 25'b0000000000000000011101000;
    rom[14371] = 25'b0000000000000000011101000;
    rom[14372] = 25'b0000000000000000011101001;
    rom[14373] = 25'b0000000000000000011101001;
    rom[14374] = 25'b0000000000000000011101001;
    rom[14375] = 25'b0000000000000000011101010;
    rom[14376] = 25'b0000000000000000011101010;
    rom[14377] = 25'b0000000000000000011101011;
    rom[14378] = 25'b0000000000000000011101011;
    rom[14379] = 25'b0000000000000000011101100;
    rom[14380] = 25'b0000000000000000011101100;
    rom[14381] = 25'b0000000000000000011101101;
    rom[14382] = 25'b0000000000000000011101101;
    rom[14383] = 25'b0000000000000000011101110;
    rom[14384] = 25'b0000000000000000011101110;
    rom[14385] = 25'b0000000000000000011101110;
    rom[14386] = 25'b0000000000000000011101110;
    rom[14387] = 25'b0000000000000000011101110;
    rom[14388] = 25'b0000000000000000011101111;
    rom[14389] = 25'b0000000000000000011101111;
    rom[14390] = 25'b0000000000000000011110000;
    rom[14391] = 25'b0000000000000000011110000;
    rom[14392] = 25'b0000000000000000011110000;
    rom[14393] = 25'b0000000000000000011110001;
    rom[14394] = 25'b0000000000000000011110001;
    rom[14395] = 25'b0000000000000000011110010;
    rom[14396] = 25'b0000000000000000011110010;
    rom[14397] = 25'b0000000000000000011110010;
    rom[14398] = 25'b0000000000000000011110010;
    rom[14399] = 25'b0000000000000000011110011;
    rom[14400] = 25'b0000000000000000011110011;
    rom[14401] = 25'b0000000000000000011110011;
    rom[14402] = 25'b0000000000000000011110100;
    rom[14403] = 25'b0000000000000000011110100;
    rom[14404] = 25'b0000000000000000011110100;
    rom[14405] = 25'b0000000000000000011110100;
    rom[14406] = 25'b0000000000000000011110100;
    rom[14407] = 25'b0000000000000000011110100;
    rom[14408] = 25'b0000000000000000011110100;
    rom[14409] = 25'b0000000000000000011110100;
    rom[14410] = 25'b0000000000000000011110100;
    rom[14411] = 25'b0000000000000000011110100;
    rom[14412] = 25'b0000000000000000011110101;
    rom[14413] = 25'b0000000000000000011110101;
    rom[14414] = 25'b0000000000000000011110101;
    rom[14415] = 25'b0000000000000000011110101;
    rom[14416] = 25'b0000000000000000011110101;
    rom[14417] = 25'b0000000000000000011110101;
    rom[14418] = 25'b0000000000000000011110101;
    rom[14419] = 25'b0000000000000000011110101;
    rom[14420] = 25'b0000000000000000011110101;
    rom[14421] = 25'b0000000000000000011110110;
    rom[14422] = 25'b0000000000000000011110110;
    rom[14423] = 25'b0000000000000000011110110;
    rom[14424] = 25'b0000000000000000011110110;
    rom[14425] = 25'b0000000000000000011110110;
    rom[14426] = 25'b0000000000000000011110110;
    rom[14427] = 25'b0000000000000000011110110;
    rom[14428] = 25'b0000000000000000011110110;
    rom[14429] = 25'b0000000000000000011110110;
    rom[14430] = 25'b0000000000000000011110110;
    rom[14431] = 25'b0000000000000000011110110;
    rom[14432] = 25'b0000000000000000011110110;
    rom[14433] = 25'b0000000000000000011110101;
    rom[14434] = 25'b0000000000000000011110101;
    rom[14435] = 25'b0000000000000000011110101;
    rom[14436] = 25'b0000000000000000011110101;
    rom[14437] = 25'b0000000000000000011110101;
    rom[14438] = 25'b0000000000000000011110101;
    rom[14439] = 25'b0000000000000000011110101;
    rom[14440] = 25'b0000000000000000011110101;
    rom[14441] = 25'b0000000000000000011110101;
    rom[14442] = 25'b0000000000000000011110101;
    rom[14443] = 25'b0000000000000000011110100;
    rom[14444] = 25'b0000000000000000011110100;
    rom[14445] = 25'b0000000000000000011110100;
    rom[14446] = 25'b0000000000000000011110100;
    rom[14447] = 25'b0000000000000000011110100;
    rom[14448] = 25'b0000000000000000011110100;
    rom[14449] = 25'b0000000000000000011110100;
    rom[14450] = 25'b0000000000000000011110100;
    rom[14451] = 25'b0000000000000000011110100;
    rom[14452] = 25'b0000000000000000011110100;
    rom[14453] = 25'b0000000000000000011110011;
    rom[14454] = 25'b0000000000000000011110011;
    rom[14455] = 25'b0000000000000000011110011;
    rom[14456] = 25'b0000000000000000011110011;
    rom[14457] = 25'b0000000000000000011110010;
    rom[14458] = 25'b0000000000000000011110010;
    rom[14459] = 25'b0000000000000000011110010;
    rom[14460] = 25'b0000000000000000011110001;
    rom[14461] = 25'b0000000000000000011110001;
    rom[14462] = 25'b0000000000000000011110001;
    rom[14463] = 25'b0000000000000000011110001;
    rom[14464] = 25'b0000000000000000011110000;
    rom[14465] = 25'b0000000000000000011110000;
    rom[14466] = 25'b0000000000000000011110000;
    rom[14467] = 25'b0000000000000000011101111;
    rom[14468] = 25'b0000000000000000011101111;
    rom[14469] = 25'b0000000000000000011101110;
    rom[14470] = 25'b0000000000000000011101110;
    rom[14471] = 25'b0000000000000000011101110;
    rom[14472] = 25'b0000000000000000011101110;
    rom[14473] = 25'b0000000000000000011101110;
    rom[14474] = 25'b0000000000000000011101101;
    rom[14475] = 25'b0000000000000000011101101;
    rom[14476] = 25'b0000000000000000011101101;
    rom[14477] = 25'b0000000000000000011101100;
    rom[14478] = 25'b0000000000000000011101100;
    rom[14479] = 25'b0000000000000000011101011;
    rom[14480] = 25'b0000000000000000011101011;
    rom[14481] = 25'b0000000000000000011101010;
    rom[14482] = 25'b0000000000000000011101010;
    rom[14483] = 25'b0000000000000000011101001;
    rom[14484] = 25'b0000000000000000011101001;
    rom[14485] = 25'b0000000000000000011101001;
    rom[14486] = 25'b0000000000000000011101001;
    rom[14487] = 25'b0000000000000000011101001;
    rom[14488] = 25'b0000000000000000011101000;
    rom[14489] = 25'b0000000000000000011101000;
    rom[14490] = 25'b0000000000000000011100111;
    rom[14491] = 25'b0000000000000000011100110;
    rom[14492] = 25'b0000000000000000011100110;
    rom[14493] = 25'b0000000000000000011100101;
    rom[14494] = 25'b0000000000000000011100101;
    rom[14495] = 25'b0000000000000000011100100;
    rom[14496] = 25'b0000000000000000011100100;
    rom[14497] = 25'b0000000000000000011100011;
    rom[14498] = 25'b0000000000000000011100011;
    rom[14499] = 25'b0000000000000000011100011;
    rom[14500] = 25'b0000000000000000011100010;
    rom[14501] = 25'b0000000000000000011100010;
    rom[14502] = 25'b0000000000000000011100001;
    rom[14503] = 25'b0000000000000000011100001;
    rom[14504] = 25'b0000000000000000011100000;
    rom[14505] = 25'b0000000000000000011011111;
    rom[14506] = 25'b0000000000000000011011111;
    rom[14507] = 25'b0000000000000000011011110;
    rom[14508] = 25'b0000000000000000011011110;
    rom[14509] = 25'b0000000000000000011011101;
    rom[14510] = 25'b0000000000000000011011101;
    rom[14511] = 25'b0000000000000000011011101;
    rom[14512] = 25'b0000000000000000011011100;
    rom[14513] = 25'b0000000000000000011011011;
    rom[14514] = 25'b0000000000000000011011011;
    rom[14515] = 25'b0000000000000000011011010;
    rom[14516] = 25'b0000000000000000011011001;
    rom[14517] = 25'b0000000000000000011011001;
    rom[14518] = 25'b0000000000000000011011000;
    rom[14519] = 25'b0000000000000000011011000;
    rom[14520] = 25'b0000000000000000011011000;
    rom[14521] = 25'b0000000000000000011010111;
    rom[14522] = 25'b0000000000000000011010110;
    rom[14523] = 25'b0000000000000000011010101;
    rom[14524] = 25'b0000000000000000011010101;
    rom[14525] = 25'b0000000000000000011010100;
    rom[14526] = 25'b0000000000000000011010011;
    rom[14527] = 25'b0000000000000000011010011;
    rom[14528] = 25'b0000000000000000011010010;
    rom[14529] = 25'b0000000000000000011010010;
    rom[14530] = 25'b0000000000000000011010001;
    rom[14531] = 25'b0000000000000000011010001;
    rom[14532] = 25'b0000000000000000011010000;
    rom[14533] = 25'b0000000000000000011001111;
    rom[14534] = 25'b0000000000000000011001110;
    rom[14535] = 25'b0000000000000000011001101;
    rom[14536] = 25'b0000000000000000011001101;
    rom[14537] = 25'b0000000000000000011001100;
    rom[14538] = 25'b0000000000000000011001100;
    rom[14539] = 25'b0000000000000000011001011;
    rom[14540] = 25'b0000000000000000011001011;
    rom[14541] = 25'b0000000000000000011001010;
    rom[14542] = 25'b0000000000000000011001001;
    rom[14543] = 25'b0000000000000000011001000;
    rom[14544] = 25'b0000000000000000011000111;
    rom[14545] = 25'b0000000000000000011000111;
    rom[14546] = 25'b0000000000000000011000111;
    rom[14547] = 25'b0000000000000000011000110;
    rom[14548] = 25'b0000000000000000011000101;
    rom[14549] = 25'b0000000000000000011000100;
    rom[14550] = 25'b0000000000000000011000011;
    rom[14551] = 25'b0000000000000000011000011;
    rom[14552] = 25'b0000000000000000011000010;
    rom[14553] = 25'b0000000000000000011000001;
    rom[14554] = 25'b0000000000000000011000001;
    rom[14555] = 25'b0000000000000000011000000;
    rom[14556] = 25'b0000000000000000010111111;
    rom[14557] = 25'b0000000000000000010111111;
    rom[14558] = 25'b0000000000000000010111110;
    rom[14559] = 25'b0000000000000000010111101;
    rom[14560] = 25'b0000000000000000010111100;
    rom[14561] = 25'b0000000000000000010111011;
    rom[14562] = 25'b0000000000000000010111011;
    rom[14563] = 25'b0000000000000000010111010;
    rom[14564] = 25'b0000000000000000010111010;
    rom[14565] = 25'b0000000000000000010111001;
    rom[14566] = 25'b0000000000000000010111000;
    rom[14567] = 25'b0000000000000000010110111;
    rom[14568] = 25'b0000000000000000010110110;
    rom[14569] = 25'b0000000000000000010110110;
    rom[14570] = 25'b0000000000000000010110101;
    rom[14571] = 25'b0000000000000000010110100;
    rom[14572] = 25'b0000000000000000010110011;
    rom[14573] = 25'b0000000000000000010110011;
    rom[14574] = 25'b0000000000000000010110010;
    rom[14575] = 25'b0000000000000000010110001;
    rom[14576] = 25'b0000000000000000010110000;
    rom[14577] = 25'b0000000000000000010110000;
    rom[14578] = 25'b0000000000000000010101111;
    rom[14579] = 25'b0000000000000000010101110;
    rom[14580] = 25'b0000000000000000010101101;
    rom[14581] = 25'b0000000000000000010101100;
    rom[14582] = 25'b0000000000000000010101011;
    rom[14583] = 25'b0000000000000000010101010;
    rom[14584] = 25'b0000000000000000010101010;
    rom[14585] = 25'b0000000000000000010101010;
    rom[14586] = 25'b0000000000000000010101001;
    rom[14587] = 25'b0000000000000000010101000;
    rom[14588] = 25'b0000000000000000010100111;
    rom[14589] = 25'b0000000000000000010100110;
    rom[14590] = 25'b0000000000000000010100101;
    rom[14591] = 25'b0000000000000000010100100;
    rom[14592] = 25'b0000000000000000010100100;
    rom[14593] = 25'b0000000000000000010100011;
    rom[14594] = 25'b0000000000000000010100010;
    rom[14595] = 25'b0000000000000000010100001;
    rom[14596] = 25'b0000000000000000010100000;
    rom[14597] = 25'b0000000000000000010011111;
    rom[14598] = 25'b0000000000000000010011111;
    rom[14599] = 25'b0000000000000000010011110;
    rom[14600] = 25'b0000000000000000010011101;
    rom[14601] = 25'b0000000000000000010011100;
    rom[14602] = 25'b0000000000000000010011011;
    rom[14603] = 25'b0000000000000000010011010;
    rom[14604] = 25'b0000000000000000010011010;
    rom[14605] = 25'b0000000000000000010011001;
    rom[14606] = 25'b0000000000000000010011001;
    rom[14607] = 25'b0000000000000000010011000;
    rom[14608] = 25'b0000000000000000010010111;
    rom[14609] = 25'b0000000000000000010010110;
    rom[14610] = 25'b0000000000000000010010101;
    rom[14611] = 25'b0000000000000000010010100;
    rom[14612] = 25'b0000000000000000010010011;
    rom[14613] = 25'b0000000000000000010010011;
    rom[14614] = 25'b0000000000000000010010010;
    rom[14615] = 25'b0000000000000000010010001;
    rom[14616] = 25'b0000000000000000010010000;
    rom[14617] = 25'b0000000000000000010001111;
    rom[14618] = 25'b0000000000000000010001110;
    rom[14619] = 25'b0000000000000000010001110;
    rom[14620] = 25'b0000000000000000010001101;
    rom[14621] = 25'b0000000000000000010001100;
    rom[14622] = 25'b0000000000000000010001011;
    rom[14623] = 25'b0000000000000000010001010;
    rom[14624] = 25'b0000000000000000010001001;
    rom[14625] = 25'b0000000000000000010001000;
    rom[14626] = 25'b0000000000000000010001000;
    rom[14627] = 25'b0000000000000000010000111;
    rom[14628] = 25'b0000000000000000010000110;
    rom[14629] = 25'b0000000000000000010000101;
    rom[14630] = 25'b0000000000000000010000100;
    rom[14631] = 25'b0000000000000000010000011;
    rom[14632] = 25'b0000000000000000010000010;
    rom[14633] = 25'b0000000000000000010000010;
    rom[14634] = 25'b0000000000000000010000001;
    rom[14635] = 25'b0000000000000000010000000;
    rom[14636] = 25'b0000000000000000001111111;
    rom[14637] = 25'b0000000000000000001111110;
    rom[14638] = 25'b0000000000000000001111101;
    rom[14639] = 25'b0000000000000000001111101;
    rom[14640] = 25'b0000000000000000001111100;
    rom[14641] = 25'b0000000000000000001111011;
    rom[14642] = 25'b0000000000000000001111010;
    rom[14643] = 25'b0000000000000000001111001;
    rom[14644] = 25'b0000000000000000001111000;
    rom[14645] = 25'b0000000000000000001111000;
    rom[14646] = 25'b0000000000000000001110111;
    rom[14647] = 25'b0000000000000000001110111;
    rom[14648] = 25'b0000000000000000001110110;
    rom[14649] = 25'b0000000000000000001110101;
    rom[14650] = 25'b0000000000000000001110100;
    rom[14651] = 25'b0000000000000000001110011;
    rom[14652] = 25'b0000000000000000001110010;
    rom[14653] = 25'b0000000000000000001110001;
    rom[14654] = 25'b0000000000000000001110001;
    rom[14655] = 25'b0000000000000000001110000;
    rom[14656] = 25'b0000000000000000001101111;
    rom[14657] = 25'b0000000000000000001101110;
    rom[14658] = 25'b0000000000000000001101101;
    rom[14659] = 25'b0000000000000000001101100;
    rom[14660] = 25'b0000000000000000001101100;
    rom[14661] = 25'b0000000000000000001101011;
    rom[14662] = 25'b0000000000000000001101010;
    rom[14663] = 25'b0000000000000000001101001;
    rom[14664] = 25'b0000000000000000001101000;
    rom[14665] = 25'b0000000000000000001100111;
    rom[14666] = 25'b0000000000000000001100110;
    rom[14667] = 25'b0000000000000000001100110;
    rom[14668] = 25'b0000000000000000001100101;
    rom[14669] = 25'b0000000000000000001100100;
    rom[14670] = 25'b0000000000000000001100011;
    rom[14671] = 25'b0000000000000000001100010;
    rom[14672] = 25'b0000000000000000001100001;
    rom[14673] = 25'b0000000000000000001100000;
    rom[14674] = 25'b0000000000000000001100000;
    rom[14675] = 25'b0000000000000000001011111;
    rom[14676] = 25'b0000000000000000001011110;
    rom[14677] = 25'b0000000000000000001011101;
    rom[14678] = 25'b0000000000000000001011100;
    rom[14679] = 25'b0000000000000000001011011;
    rom[14680] = 25'b0000000000000000001011011;
    rom[14681] = 25'b0000000000000000001011011;
    rom[14682] = 25'b0000000000000000001011010;
    rom[14683] = 25'b0000000000000000001011001;
    rom[14684] = 25'b0000000000000000001011000;
    rom[14685] = 25'b0000000000000000001010111;
    rom[14686] = 25'b0000000000000000001010110;
    rom[14687] = 25'b0000000000000000001010101;
    rom[14688] = 25'b0000000000000000001010101;
    rom[14689] = 25'b0000000000000000001010100;
    rom[14690] = 25'b0000000000000000001010011;
    rom[14691] = 25'b0000000000000000001010010;
    rom[14692] = 25'b0000000000000000001010001;
    rom[14693] = 25'b0000000000000000001010000;
    rom[14694] = 25'b0000000000000000001001111;
    rom[14695] = 25'b0000000000000000001001111;
    rom[14696] = 25'b0000000000000000001001110;
    rom[14697] = 25'b0000000000000000001001110;
    rom[14698] = 25'b0000000000000000001001101;
    rom[14699] = 25'b0000000000000000001001100;
    rom[14700] = 25'b0000000000000000001001011;
    rom[14701] = 25'b0000000000000000001001010;
    rom[14702] = 25'b0000000000000000001001001;
    rom[14703] = 25'b0000000000000000001001001;
    rom[14704] = 25'b0000000000000000001001000;
    rom[14705] = 25'b0000000000000000001000111;
    rom[14706] = 25'b0000000000000000001000110;
    rom[14707] = 25'b0000000000000000001000101;
    rom[14708] = 25'b0000000000000000001000100;
    rom[14709] = 25'b0000000000000000001000100;
    rom[14710] = 25'b0000000000000000001000100;
    rom[14711] = 25'b0000000000000000001000011;
    rom[14712] = 25'b0000000000000000001000010;
    rom[14713] = 25'b0000000000000000001000001;
    rom[14714] = 25'b0000000000000000001000000;
    rom[14715] = 25'b0000000000000000000111111;
    rom[14716] = 25'b0000000000000000000111110;
    rom[14717] = 25'b0000000000000000000111110;
    rom[14718] = 25'b0000000000000000000111101;
    rom[14719] = 25'b0000000000000000000111101;
    rom[14720] = 25'b0000000000000000000111100;
    rom[14721] = 25'b0000000000000000000111011;
    rom[14722] = 25'b0000000000000000000111010;
    rom[14723] = 25'b0000000000000000000111001;
    rom[14724] = 25'b0000000000000000000111000;
    rom[14725] = 25'b0000000000000000000111000;
    rom[14726] = 25'b0000000000000000000110111;
    rom[14727] = 25'b0000000000000000000110111;
    rom[14728] = 25'b0000000000000000000110110;
    rom[14729] = 25'b0000000000000000000110101;
    rom[14730] = 25'b0000000000000000000110100;
    rom[14731] = 25'b0000000000000000000110011;
    rom[14732] = 25'b0000000000000000000110011;
    rom[14733] = 25'b0000000000000000000110010;
    rom[14734] = 25'b0000000000000000000110001;
    rom[14735] = 25'b0000000000000000000110001;
    rom[14736] = 25'b0000000000000000000110000;
    rom[14737] = 25'b0000000000000000000101111;
    rom[14738] = 25'b0000000000000000000101110;
    rom[14739] = 25'b0000000000000000000101101;
    rom[14740] = 25'b0000000000000000000101101;
    rom[14741] = 25'b0000000000000000000101101;
    rom[14742] = 25'b0000000000000000000101100;
    rom[14743] = 25'b0000000000000000000101011;
    rom[14744] = 25'b0000000000000000000101010;
    rom[14745] = 25'b0000000000000000000101001;
    rom[14746] = 25'b0000000000000000000101000;
    rom[14747] = 25'b0000000000000000000101000;
    rom[14748] = 25'b0000000000000000000100111;
    rom[14749] = 25'b0000000000000000000100111;
    rom[14750] = 25'b0000000000000000000100110;
    rom[14751] = 25'b0000000000000000000100101;
    rom[14752] = 25'b0000000000000000000100101;
    rom[14753] = 25'b0000000000000000000100100;
    rom[14754] = 25'b0000000000000000000100011;
    rom[14755] = 25'b0000000000000000000100010;
    rom[14756] = 25'b0000000000000000000100010;
    rom[14757] = 25'b0000000000000000000100010;
    rom[14758] = 25'b0000000000000000000100001;
    rom[14759] = 25'b0000000000000000000100000;
    rom[14760] = 25'b0000000000000000000011111;
    rom[14761] = 25'b0000000000000000000011110;
    rom[14762] = 25'b0000000000000000000011110;
    rom[14763] = 25'b0000000000000000000011101;
    rom[14764] = 25'b0000000000000000000011100;
    rom[14765] = 25'b0000000000000000000011100;
    rom[14766] = 25'b0000000000000000000011100;
    rom[14767] = 25'b0000000000000000000011011;
    rom[14768] = 25'b0000000000000000000011010;
    rom[14769] = 25'b0000000000000000000011001;
    rom[14770] = 25'b0000000000000000000011001;
    rom[14771] = 25'b0000000000000000000011000;
    rom[14772] = 25'b0000000000000000000010111;
    rom[14773] = 25'b0000000000000000000010110;
    rom[14774] = 25'b0000000000000000000010110;
    rom[14775] = 25'b0000000000000000000010110;
    rom[14776] = 25'b0000000000000000000010101;
    rom[14777] = 25'b0000000000000000000010100;
    rom[14778] = 25'b0000000000000000000010100;
    rom[14779] = 25'b0000000000000000000010011;
    rom[14780] = 25'b0000000000000000000010010;
    rom[14781] = 25'b0000000000000000000010001;
    rom[14782] = 25'b0000000000000000000010001;
    rom[14783] = 25'b0000000000000000000010001;
    rom[14784] = 25'b0000000000000000000010000;
    rom[14785] = 25'b0000000000000000000010000;
    rom[14786] = 25'b0000000000000000000001111;
    rom[14787] = 25'b0000000000000000000001110;
    rom[14788] = 25'b0000000000000000000001101;
    rom[14789] = 25'b0000000000000000000001101;
    rom[14790] = 25'b0000000000000000000001100;
    rom[14791] = 25'b0000000000000000000001011;
    rom[14792] = 25'b0000000000000000000001011;
    rom[14793] = 25'b0000000000000000000001011;
    rom[14794] = 25'b0000000000000000000001010;
    rom[14795] = 25'b0000000000000000000001010;
    rom[14796] = 25'b0000000000000000000001001;
    rom[14797] = 25'b0000000000000000000001000;
    rom[14798] = 25'b0000000000000000000001000;
    rom[14799] = 25'b0000000000000000000000111;
    rom[14800] = 25'b0000000000000000000000110;
    rom[14801] = 25'b0000000000000000000000110;
    rom[14802] = 25'b0000000000000000000000101;
    rom[14803] = 25'b0000000000000000000000101;
    rom[14804] = 25'b0000000000000000000000101;
    rom[14805] = 25'b0000000000000000000000100;
    rom[14806] = 25'b0000000000000000000000011;
    rom[14807] = 25'b0000000000000000000000011;
    rom[14808] = 25'b0000000000000000000000010;
    rom[14809] = 25'b0000000000000000000000001;
    rom[14810] = 25'b0000000000000000000000001;
    rom[14811] = 25'b0000000000000000000000000;
    rom[14812] = 25'b0000000000000000000000000;
    rom[14813] = 25'b0000000000000000000000000;
    rom[14814] = 25'b0000000000000000000000000;
    rom[14815] = 25'b0000000000000000000000000;
    rom[14816] = 25'b1111111111111111111111111;
    rom[14817] = 25'b1111111111111111111111111;
    rom[14818] = 25'b1111111111111111111111110;
    rom[14819] = 25'b1111111111111111111111101;
    rom[14820] = 25'b1111111111111111111111101;
    rom[14821] = 25'b1111111111111111111111100;
    rom[14822] = 25'b1111111111111111111111100;
    rom[14823] = 25'b1111111111111111111111011;
    rom[14824] = 25'b1111111111111111111111010;
    rom[14825] = 25'b1111111111111111111111010;
    rom[14826] = 25'b1111111111111111111111010;
    rom[14827] = 25'b1111111111111111111111010;
    rom[14828] = 25'b1111111111111111111111001;
    rom[14829] = 25'b1111111111111111111111001;
    rom[14830] = 25'b1111111111111111111111000;
    rom[14831] = 25'b1111111111111111111110111;
    rom[14832] = 25'b1111111111111111111110111;
    rom[14833] = 25'b1111111111111111111110110;
    rom[14834] = 25'b1111111111111111111110110;
    rom[14835] = 25'b1111111111111111111110101;
    rom[14836] = 25'b1111111111111111111110101;
    rom[14837] = 25'b1111111111111111111110100;
    rom[14838] = 25'b1111111111111111111110100;
    rom[14839] = 25'b1111111111111111111110100;
    rom[14840] = 25'b1111111111111111111110100;
    rom[14841] = 25'b1111111111111111111110011;
    rom[14842] = 25'b1111111111111111111110010;
    rom[14843] = 25'b1111111111111111111110010;
    rom[14844] = 25'b1111111111111111111110001;
    rom[14845] = 25'b1111111111111111111110001;
    rom[14846] = 25'b1111111111111111111110000;
    rom[14847] = 25'b1111111111111111111110000;
    rom[14848] = 25'b1111111111111111111101111;
    rom[14849] = 25'b1111111111111111111101111;
    rom[14850] = 25'b1111111111111111111101110;
    rom[14851] = 25'b1111111111111111111101110;
    rom[14852] = 25'b1111111111111111111101110;
    rom[14853] = 25'b1111111111111111111101110;
    rom[14854] = 25'b1111111111111111111101101;
    rom[14855] = 25'b1111111111111111111101101;
    rom[14856] = 25'b1111111111111111111101100;
    rom[14857] = 25'b1111111111111111111101100;
    rom[14858] = 25'b1111111111111111111101100;
    rom[14859] = 25'b1111111111111111111101011;
    rom[14860] = 25'b1111111111111111111101011;
    rom[14861] = 25'b1111111111111111111101010;
    rom[14862] = 25'b1111111111111111111101010;
    rom[14863] = 25'b1111111111111111111101001;
    rom[14864] = 25'b1111111111111111111101001;
    rom[14865] = 25'b1111111111111111111101001;
    rom[14866] = 25'b1111111111111111111101001;
    rom[14867] = 25'b1111111111111111111101000;
    rom[14868] = 25'b1111111111111111111101000;
    rom[14869] = 25'b1111111111111111111101000;
    rom[14870] = 25'b1111111111111111111100111;
    rom[14871] = 25'b1111111111111111111100111;
    rom[14872] = 25'b1111111111111111111100110;
    rom[14873] = 25'b1111111111111111111100110;
    rom[14874] = 25'b1111111111111111111100101;
    rom[14875] = 25'b1111111111111111111100101;
    rom[14876] = 25'b1111111111111111111100101;
    rom[14877] = 25'b1111111111111111111100100;
    rom[14878] = 25'b1111111111111111111100100;
    rom[14879] = 25'b1111111111111111111100011;
    rom[14880] = 25'b1111111111111111111100011;
    rom[14881] = 25'b1111111111111111111100011;
    rom[14882] = 25'b1111111111111111111100011;
    rom[14883] = 25'b1111111111111111111100011;
    rom[14884] = 25'b1111111111111111111100010;
    rom[14885] = 25'b1111111111111111111100010;
    rom[14886] = 25'b1111111111111111111100010;
    rom[14887] = 25'b1111111111111111111100001;
    rom[14888] = 25'b1111111111111111111100001;
    rom[14889] = 25'b1111111111111111111100001;
    rom[14890] = 25'b1111111111111111111100000;
    rom[14891] = 25'b1111111111111111111100000;
    rom[14892] = 25'b1111111111111111111100000;
    rom[14893] = 25'b1111111111111111111011111;
    rom[14894] = 25'b1111111111111111111011111;
    rom[14895] = 25'b1111111111111111111011110;
    rom[14896] = 25'b1111111111111111111011110;
    rom[14897] = 25'b1111111111111111111011110;
    rom[14898] = 25'b1111111111111111111011101;
    rom[14899] = 25'b1111111111111111111011101;
    rom[14900] = 25'b1111111111111111111011101;
    rom[14901] = 25'b1111111111111111111011101;
    rom[14902] = 25'b1111111111111111111011101;
    rom[14903] = 25'b1111111111111111111011101;
    rom[14904] = 25'b1111111111111111111011100;
    rom[14905] = 25'b1111111111111111111011100;
    rom[14906] = 25'b1111111111111111111011100;
    rom[14907] = 25'b1111111111111111111011100;
    rom[14908] = 25'b1111111111111111111011011;
    rom[14909] = 25'b1111111111111111111011011;
    rom[14910] = 25'b1111111111111111111011011;
    rom[14911] = 25'b1111111111111111111011010;
    rom[14912] = 25'b1111111111111111111011010;
    rom[14913] = 25'b1111111111111111111011010;
    rom[14914] = 25'b1111111111111111111011001;
    rom[14915] = 25'b1111111111111111111011001;
    rom[14916] = 25'b1111111111111111111011001;
    rom[14917] = 25'b1111111111111111111011001;
    rom[14918] = 25'b1111111111111111111011000;
    rom[14919] = 25'b1111111111111111111011000;
    rom[14920] = 25'b1111111111111111111011000;
    rom[14921] = 25'b1111111111111111111011000;
    rom[14922] = 25'b1111111111111111111011000;
    rom[14923] = 25'b1111111111111111111011000;
    rom[14924] = 25'b1111111111111111111011000;
    rom[14925] = 25'b1111111111111111111011000;
    rom[14926] = 25'b1111111111111111111010111;
    rom[14927] = 25'b1111111111111111111010111;
    rom[14928] = 25'b1111111111111111111010111;
    rom[14929] = 25'b1111111111111111111010111;
    rom[14930] = 25'b1111111111111111111010110;
    rom[14931] = 25'b1111111111111111111010110;
    rom[14932] = 25'b1111111111111111111010110;
    rom[14933] = 25'b1111111111111111111010110;
    rom[14934] = 25'b1111111111111111111010101;
    rom[14935] = 25'b1111111111111111111010101;
    rom[14936] = 25'b1111111111111111111010101;
    rom[14937] = 25'b1111111111111111111010101;
    rom[14938] = 25'b1111111111111111111010100;
    rom[14939] = 25'b1111111111111111111010100;
    rom[14940] = 25'b1111111111111111111010100;
    rom[14941] = 25'b1111111111111111111010100;
    rom[14942] = 25'b1111111111111111111010100;
    rom[14943] = 25'b1111111111111111111010011;
    rom[14944] = 25'b1111111111111111111010011;
    rom[14945] = 25'b1111111111111111111010011;
    rom[14946] = 25'b1111111111111111111010011;
    rom[14947] = 25'b1111111111111111111010011;
    rom[14948] = 25'b1111111111111111111010011;
    rom[14949] = 25'b1111111111111111111010010;
    rom[14950] = 25'b1111111111111111111010010;
    rom[14951] = 25'b1111111111111111111010010;
    rom[14952] = 25'b1111111111111111111010010;
    rom[14953] = 25'b1111111111111111111010010;
    rom[14954] = 25'b1111111111111111111010010;
    rom[14955] = 25'b1111111111111111111010010;
    rom[14956] = 25'b1111111111111111111010010;
    rom[14957] = 25'b1111111111111111111010010;
    rom[14958] = 25'b1111111111111111111010010;
    rom[14959] = 25'b1111111111111111111010010;
    rom[14960] = 25'b1111111111111111111010010;
    rom[14961] = 25'b1111111111111111111010001;
    rom[14962] = 25'b1111111111111111111010001;
    rom[14963] = 25'b1111111111111111111010001;
    rom[14964] = 25'b1111111111111111111010001;
    rom[14965] = 25'b1111111111111111111010001;
    rom[14966] = 25'b1111111111111111111010001;
    rom[14967] = 25'b1111111111111111111010001;
    rom[14968] = 25'b1111111111111111111010000;
    rom[14969] = 25'b1111111111111111111010000;
    rom[14970] = 25'b1111111111111111111010000;
    rom[14971] = 25'b1111111111111111111010000;
    rom[14972] = 25'b1111111111111111111010000;
    rom[14973] = 25'b1111111111111111111010000;
    rom[14974] = 25'b1111111111111111111010000;
    rom[14975] = 25'b1111111111111111111010000;
    rom[14976] = 25'b1111111111111111111001111;
    rom[14977] = 25'b1111111111111111111001111;
    rom[14978] = 25'b1111111111111111111001111;
    rom[14979] = 25'b1111111111111111111001111;
    rom[14980] = 25'b1111111111111111111001111;
    rom[14981] = 25'b1111111111111111111001111;
    rom[14982] = 25'b1111111111111111111001111;
    rom[14983] = 25'b1111111111111111111001111;
    rom[14984] = 25'b1111111111111111111001111;
    rom[14985] = 25'b1111111111111111111001111;
    rom[14986] = 25'b1111111111111111111001110;
    rom[14987] = 25'b1111111111111111111001110;
    rom[14988] = 25'b1111111111111111111001110;
    rom[14989] = 25'b1111111111111111111001110;
    rom[14990] = 25'b1111111111111111111001110;
    rom[14991] = 25'b1111111111111111111001110;
    rom[14992] = 25'b1111111111111111111001110;
    rom[14993] = 25'b1111111111111111111001110;
    rom[14994] = 25'b1111111111111111111001110;
    rom[14995] = 25'b1111111111111111111001110;
    rom[14996] = 25'b1111111111111111111001110;
    rom[14997] = 25'b1111111111111111111001110;
    rom[14998] = 25'b1111111111111111111001110;
    rom[14999] = 25'b1111111111111111111001110;
    rom[15000] = 25'b1111111111111111111001110;
    rom[15001] = 25'b1111111111111111111001110;
    rom[15002] = 25'b1111111111111111111001101;
    rom[15003] = 25'b1111111111111111111001101;
    rom[15004] = 25'b1111111111111111111001101;
    rom[15005] = 25'b1111111111111111111001101;
    rom[15006] = 25'b1111111111111111111001101;
    rom[15007] = 25'b1111111111111111111001101;
    rom[15008] = 25'b1111111111111111111001101;
    rom[15009] = 25'b1111111111111111111001101;
    rom[15010] = 25'b1111111111111111111001101;
    rom[15011] = 25'b1111111111111111111001101;
    rom[15012] = 25'b1111111111111111111001101;
    rom[15013] = 25'b1111111111111111111001101;
    rom[15014] = 25'b1111111111111111111001101;
    rom[15015] = 25'b1111111111111111111001101;
    rom[15016] = 25'b1111111111111111111001101;
    rom[15017] = 25'b1111111111111111111001101;
    rom[15018] = 25'b1111111111111111111001101;
    rom[15019] = 25'b1111111111111111111001101;
    rom[15020] = 25'b1111111111111111111001101;
    rom[15021] = 25'b1111111111111111111001101;
    rom[15022] = 25'b1111111111111111111001101;
    rom[15023] = 25'b1111111111111111111001101;
    rom[15024] = 25'b1111111111111111111001101;
    rom[15025] = 25'b1111111111111111111001101;
    rom[15026] = 25'b1111111111111111111001101;
    rom[15027] = 25'b1111111111111111111001101;
    rom[15028] = 25'b1111111111111111111001101;
    rom[15029] = 25'b1111111111111111111001101;
    rom[15030] = 25'b1111111111111111111001101;
    rom[15031] = 25'b1111111111111111111001101;
    rom[15032] = 25'b1111111111111111111001101;
    rom[15033] = 25'b1111111111111111111001101;
    rom[15034] = 25'b1111111111111111111001101;
    rom[15035] = 25'b1111111111111111111001101;
    rom[15036] = 25'b1111111111111111111001101;
    rom[15037] = 25'b1111111111111111111001101;
    rom[15038] = 25'b1111111111111111111001101;
    rom[15039] = 25'b1111111111111111111001101;
    rom[15040] = 25'b1111111111111111111001101;
    rom[15041] = 25'b1111111111111111111001101;
    rom[15042] = 25'b1111111111111111111001101;
    rom[15043] = 25'b1111111111111111111001110;
    rom[15044] = 25'b1111111111111111111001110;
    rom[15045] = 25'b1111111111111111111001110;
    rom[15046] = 25'b1111111111111111111001110;
    rom[15047] = 25'b1111111111111111111001110;
    rom[15048] = 25'b1111111111111111111001110;
    rom[15049] = 25'b1111111111111111111001110;
    rom[15050] = 25'b1111111111111111111001110;
    rom[15051] = 25'b1111111111111111111001110;
    rom[15052] = 25'b1111111111111111111001110;
    rom[15053] = 25'b1111111111111111111001110;
    rom[15054] = 25'b1111111111111111111001110;
    rom[15055] = 25'b1111111111111111111001110;
    rom[15056] = 25'b1111111111111111111001110;
    rom[15057] = 25'b1111111111111111111001110;
    rom[15058] = 25'b1111111111111111111001110;
    rom[15059] = 25'b1111111111111111111001110;
    rom[15060] = 25'b1111111111111111111001110;
    rom[15061] = 25'b1111111111111111111001111;
    rom[15062] = 25'b1111111111111111111001111;
    rom[15063] = 25'b1111111111111111111001111;
    rom[15064] = 25'b1111111111111111111001111;
    rom[15065] = 25'b1111111111111111111001111;
    rom[15066] = 25'b1111111111111111111001111;
    rom[15067] = 25'b1111111111111111111001111;
    rom[15068] = 25'b1111111111111111111001111;
    rom[15069] = 25'b1111111111111111111001111;
    rom[15070] = 25'b1111111111111111111001111;
    rom[15071] = 25'b1111111111111111111001111;
    rom[15072] = 25'b1111111111111111111001111;
    rom[15073] = 25'b1111111111111111111010000;
    rom[15074] = 25'b1111111111111111111010000;
    rom[15075] = 25'b1111111111111111111010000;
    rom[15076] = 25'b1111111111111111111010000;
    rom[15077] = 25'b1111111111111111111010000;
    rom[15078] = 25'b1111111111111111111010000;
    rom[15079] = 25'b1111111111111111111010000;
    rom[15080] = 25'b1111111111111111111010000;
    rom[15081] = 25'b1111111111111111111010000;
    rom[15082] = 25'b1111111111111111111010000;
    rom[15083] = 25'b1111111111111111111010001;
    rom[15084] = 25'b1111111111111111111010001;
    rom[15085] = 25'b1111111111111111111010001;
    rom[15086] = 25'b1111111111111111111010001;
    rom[15087] = 25'b1111111111111111111010001;
    rom[15088] = 25'b1111111111111111111010001;
    rom[15089] = 25'b1111111111111111111010001;
    rom[15090] = 25'b1111111111111111111010001;
    rom[15091] = 25'b1111111111111111111010001;
    rom[15092] = 25'b1111111111111111111010010;
    rom[15093] = 25'b1111111111111111111010010;
    rom[15094] = 25'b1111111111111111111010010;
    rom[15095] = 25'b1111111111111111111010010;
    rom[15096] = 25'b1111111111111111111010010;
    rom[15097] = 25'b1111111111111111111010010;
    rom[15098] = 25'b1111111111111111111010010;
    rom[15099] = 25'b1111111111111111111010010;
    rom[15100] = 25'b1111111111111111111010010;
    rom[15101] = 25'b1111111111111111111010010;
    rom[15102] = 25'b1111111111111111111010010;
    rom[15103] = 25'b1111111111111111111010010;
    rom[15104] = 25'b1111111111111111111010010;
    rom[15105] = 25'b1111111111111111111010010;
    rom[15106] = 25'b1111111111111111111010010;
    rom[15107] = 25'b1111111111111111111010010;
    rom[15108] = 25'b1111111111111111111010011;
    rom[15109] = 25'b1111111111111111111010011;
    rom[15110] = 25'b1111111111111111111010011;
    rom[15111] = 25'b1111111111111111111010011;
    rom[15112] = 25'b1111111111111111111010011;
    rom[15113] = 25'b1111111111111111111010011;
    rom[15114] = 25'b1111111111111111111010011;
    rom[15115] = 25'b1111111111111111111010100;
    rom[15116] = 25'b1111111111111111111010100;
    rom[15117] = 25'b1111111111111111111010100;
    rom[15118] = 25'b1111111111111111111010100;
    rom[15119] = 25'b1111111111111111111010100;
    rom[15120] = 25'b1111111111111111111010100;
    rom[15121] = 25'b1111111111111111111010100;
    rom[15122] = 25'b1111111111111111111010101;
    rom[15123] = 25'b1111111111111111111010101;
    rom[15124] = 25'b1111111111111111111010101;
    rom[15125] = 25'b1111111111111111111010101;
    rom[15126] = 25'b1111111111111111111010101;
    rom[15127] = 25'b1111111111111111111010101;
    rom[15128] = 25'b1111111111111111111010110;
    rom[15129] = 25'b1111111111111111111010110;
    rom[15130] = 25'b1111111111111111111010110;
    rom[15131] = 25'b1111111111111111111010110;
    rom[15132] = 25'b1111111111111111111010110;
    rom[15133] = 25'b1111111111111111111010110;
    rom[15134] = 25'b1111111111111111111010111;
    rom[15135] = 25'b1111111111111111111010111;
    rom[15136] = 25'b1111111111111111111010111;
    rom[15137] = 25'b1111111111111111111010111;
    rom[15138] = 25'b1111111111111111111010111;
    rom[15139] = 25'b1111111111111111111010111;
    rom[15140] = 25'b1111111111111111111011000;
    rom[15141] = 25'b1111111111111111111011000;
    rom[15142] = 25'b1111111111111111111011000;
    rom[15143] = 25'b1111111111111111111011000;
    rom[15144] = 25'b1111111111111111111011000;
    rom[15145] = 25'b1111111111111111111011000;
    rom[15146] = 25'b1111111111111111111011000;
    rom[15147] = 25'b1111111111111111111011000;
    rom[15148] = 25'b1111111111111111111011000;
    rom[15149] = 25'b1111111111111111111011000;
    rom[15150] = 25'b1111111111111111111011000;
    rom[15151] = 25'b1111111111111111111011000;
    rom[15152] = 25'b1111111111111111111011001;
    rom[15153] = 25'b1111111111111111111011001;
    rom[15154] = 25'b1111111111111111111011001;
    rom[15155] = 25'b1111111111111111111011001;
    rom[15156] = 25'b1111111111111111111011001;
    rom[15157] = 25'b1111111111111111111011001;
    rom[15158] = 25'b1111111111111111111011010;
    rom[15159] = 25'b1111111111111111111011010;
    rom[15160] = 25'b1111111111111111111011010;
    rom[15161] = 25'b1111111111111111111011010;
    rom[15162] = 25'b1111111111111111111011010;
    rom[15163] = 25'b1111111111111111111011011;
    rom[15164] = 25'b1111111111111111111011011;
    rom[15165] = 25'b1111111111111111111011011;
    rom[15166] = 25'b1111111111111111111011011;
    rom[15167] = 25'b1111111111111111111011011;
    rom[15168] = 25'b1111111111111111111011011;
    rom[15169] = 25'b1111111111111111111011100;
    rom[15170] = 25'b1111111111111111111011100;
    rom[15171] = 25'b1111111111111111111011100;
    rom[15172] = 25'b1111111111111111111011100;
    rom[15173] = 25'b1111111111111111111011100;
    rom[15174] = 25'b1111111111111111111011101;
    rom[15175] = 25'b1111111111111111111011101;
    rom[15176] = 25'b1111111111111111111011101;
    rom[15177] = 25'b1111111111111111111011101;
    rom[15178] = 25'b1111111111111111111011101;
    rom[15179] = 25'b1111111111111111111011101;
    rom[15180] = 25'b1111111111111111111011101;
    rom[15181] = 25'b1111111111111111111011101;
    rom[15182] = 25'b1111111111111111111011101;
    rom[15183] = 25'b1111111111111111111011101;
    rom[15184] = 25'b1111111111111111111011101;
    rom[15185] = 25'b1111111111111111111011110;
    rom[15186] = 25'b1111111111111111111011110;
    rom[15187] = 25'b1111111111111111111011110;
    rom[15188] = 25'b1111111111111111111011110;
    rom[15189] = 25'b1111111111111111111011110;
    rom[15190] = 25'b1111111111111111111011111;
    rom[15191] = 25'b1111111111111111111011111;
    rom[15192] = 25'b1111111111111111111011111;
    rom[15193] = 25'b1111111111111111111011111;
    rom[15194] = 25'b1111111111111111111011111;
    rom[15195] = 25'b1111111111111111111100000;
    rom[15196] = 25'b1111111111111111111100000;
    rom[15197] = 25'b1111111111111111111100000;
    rom[15198] = 25'b1111111111111111111100000;
    rom[15199] = 25'b1111111111111111111100000;
    rom[15200] = 25'b1111111111111111111100001;
    rom[15201] = 25'b1111111111111111111100001;
    rom[15202] = 25'b1111111111111111111100001;
    rom[15203] = 25'b1111111111111111111100001;
    rom[15204] = 25'b1111111111111111111100001;
    rom[15205] = 25'b1111111111111111111100010;
    rom[15206] = 25'b1111111111111111111100010;
    rom[15207] = 25'b1111111111111111111100010;
    rom[15208] = 25'b1111111111111111111100010;
    rom[15209] = 25'b1111111111111111111100010;
    rom[15210] = 25'b1111111111111111111100011;
    rom[15211] = 25'b1111111111111111111100011;
    rom[15212] = 25'b1111111111111111111100011;
    rom[15213] = 25'b1111111111111111111100011;
    rom[15214] = 25'b1111111111111111111100011;
    rom[15215] = 25'b1111111111111111111100011;
    rom[15216] = 25'b1111111111111111111100011;
    rom[15217] = 25'b1111111111111111111100011;
    rom[15218] = 25'b1111111111111111111100011;
    rom[15219] = 25'b1111111111111111111100011;
    rom[15220] = 25'b1111111111111111111100100;
    rom[15221] = 25'b1111111111111111111100100;
    rom[15222] = 25'b1111111111111111111100100;
    rom[15223] = 25'b1111111111111111111100100;
    rom[15224] = 25'b1111111111111111111100100;
    rom[15225] = 25'b1111111111111111111100101;
    rom[15226] = 25'b1111111111111111111100101;
    rom[15227] = 25'b1111111111111111111100101;
    rom[15228] = 25'b1111111111111111111100101;
    rom[15229] = 25'b1111111111111111111100101;
    rom[15230] = 25'b1111111111111111111100110;
    rom[15231] = 25'b1111111111111111111100110;
    rom[15232] = 25'b1111111111111111111100110;
    rom[15233] = 25'b1111111111111111111100110;
    rom[15234] = 25'b1111111111111111111100110;
    rom[15235] = 25'b1111111111111111111100111;
    rom[15236] = 25'b1111111111111111111100111;
    rom[15237] = 25'b1111111111111111111100111;
    rom[15238] = 25'b1111111111111111111100111;
    rom[15239] = 25'b1111111111111111111100111;
    rom[15240] = 25'b1111111111111111111101000;
    rom[15241] = 25'b1111111111111111111101000;
    rom[15242] = 25'b1111111111111111111101000;
    rom[15243] = 25'b1111111111111111111101000;
    rom[15244] = 25'b1111111111111111111101000;
    rom[15245] = 25'b1111111111111111111101001;
    rom[15246] = 25'b1111111111111111111101001;
    rom[15247] = 25'b1111111111111111111101001;
    rom[15248] = 25'b1111111111111111111101001;
    rom[15249] = 25'b1111111111111111111101001;
    rom[15250] = 25'b1111111111111111111101001;
    rom[15251] = 25'b1111111111111111111101001;
    rom[15252] = 25'b1111111111111111111101001;
    rom[15253] = 25'b1111111111111111111101001;
    rom[15254] = 25'b1111111111111111111101001;
    rom[15255] = 25'b1111111111111111111101010;
    rom[15256] = 25'b1111111111111111111101010;
    rom[15257] = 25'b1111111111111111111101010;
    rom[15258] = 25'b1111111111111111111101010;
    rom[15259] = 25'b1111111111111111111101010;
    rom[15260] = 25'b1111111111111111111101010;
    rom[15261] = 25'b1111111111111111111101011;
    rom[15262] = 25'b1111111111111111111101011;
    rom[15263] = 25'b1111111111111111111101011;
    rom[15264] = 25'b1111111111111111111101011;
    rom[15265] = 25'b1111111111111111111101011;
    rom[15266] = 25'b1111111111111111111101100;
    rom[15267] = 25'b1111111111111111111101100;
    rom[15268] = 25'b1111111111111111111101100;
    rom[15269] = 25'b1111111111111111111101100;
    rom[15270] = 25'b1111111111111111111101100;
    rom[15271] = 25'b1111111111111111111101101;
    rom[15272] = 25'b1111111111111111111101101;
    rom[15273] = 25'b1111111111111111111101101;
    rom[15274] = 25'b1111111111111111111101101;
    rom[15275] = 25'b1111111111111111111101101;
    rom[15276] = 25'b1111111111111111111101110;
    rom[15277] = 25'b1111111111111111111101110;
    rom[15278] = 25'b1111111111111111111101110;
    rom[15279] = 25'b1111111111111111111101110;
    rom[15280] = 25'b1111111111111111111101110;
    rom[15281] = 25'b1111111111111111111101110;
    rom[15282] = 25'b1111111111111111111101110;
    rom[15283] = 25'b1111111111111111111101110;
    rom[15284] = 25'b1111111111111111111101110;
    rom[15285] = 25'b1111111111111111111101110;
    rom[15286] = 25'b1111111111111111111101110;
    rom[15287] = 25'b1111111111111111111101111;
    rom[15288] = 25'b1111111111111111111101111;
    rom[15289] = 25'b1111111111111111111101111;
    rom[15290] = 25'b1111111111111111111101111;
    rom[15291] = 25'b1111111111111111111101111;
    rom[15292] = 25'b1111111111111111111110000;
    rom[15293] = 25'b1111111111111111111110000;
    rom[15294] = 25'b1111111111111111111110000;
    rom[15295] = 25'b1111111111111111111110000;
    rom[15296] = 25'b1111111111111111111110000;
    rom[15297] = 25'b1111111111111111111110001;
    rom[15298] = 25'b1111111111111111111110001;
    rom[15299] = 25'b1111111111111111111110001;
    rom[15300] = 25'b1111111111111111111110001;
    rom[15301] = 25'b1111111111111111111110001;
    rom[15302] = 25'b1111111111111111111110001;
    rom[15303] = 25'b1111111111111111111110010;
    rom[15304] = 25'b1111111111111111111110010;
    rom[15305] = 25'b1111111111111111111110010;
    rom[15306] = 25'b1111111111111111111110010;
    rom[15307] = 25'b1111111111111111111110010;
    rom[15308] = 25'b1111111111111111111110011;
    rom[15309] = 25'b1111111111111111111110011;
    rom[15310] = 25'b1111111111111111111110011;
    rom[15311] = 25'b1111111111111111111110011;
    rom[15312] = 25'b1111111111111111111110011;
    rom[15313] = 25'b1111111111111111111110011;
    rom[15314] = 25'b1111111111111111111110100;
    rom[15315] = 25'b1111111111111111111110100;
    rom[15316] = 25'b1111111111111111111110100;
    rom[15317] = 25'b1111111111111111111110100;
    rom[15318] = 25'b1111111111111111111110100;
    rom[15319] = 25'b1111111111111111111110100;
    rom[15320] = 25'b1111111111111111111110100;
    rom[15321] = 25'b1111111111111111111110100;
    rom[15322] = 25'b1111111111111111111110100;
    rom[15323] = 25'b1111111111111111111110100;
    rom[15324] = 25'b1111111111111111111110100;
    rom[15325] = 25'b1111111111111111111110100;
    rom[15326] = 25'b1111111111111111111110101;
    rom[15327] = 25'b1111111111111111111110101;
    rom[15328] = 25'b1111111111111111111110101;
    rom[15329] = 25'b1111111111111111111110101;
    rom[15330] = 25'b1111111111111111111110101;
    rom[15331] = 25'b1111111111111111111110110;
    rom[15332] = 25'b1111111111111111111110110;
    rom[15333] = 25'b1111111111111111111110110;
    rom[15334] = 25'b1111111111111111111110110;
    rom[15335] = 25'b1111111111111111111110110;
    rom[15336] = 25'b1111111111111111111110110;
    rom[15337] = 25'b1111111111111111111110111;
    rom[15338] = 25'b1111111111111111111110111;
    rom[15339] = 25'b1111111111111111111110111;
    rom[15340] = 25'b1111111111111111111110111;
    rom[15341] = 25'b1111111111111111111110111;
    rom[15342] = 25'b1111111111111111111110111;
    rom[15343] = 25'b1111111111111111111110111;
    rom[15344] = 25'b1111111111111111111111000;
    rom[15345] = 25'b1111111111111111111111000;
    rom[15346] = 25'b1111111111111111111111000;
    rom[15347] = 25'b1111111111111111111111000;
    rom[15348] = 25'b1111111111111111111111000;
    rom[15349] = 25'b1111111111111111111111000;
    rom[15350] = 25'b1111111111111111111111001;
    rom[15351] = 25'b1111111111111111111111001;
    rom[15352] = 25'b1111111111111111111111001;
    rom[15353] = 25'b1111111111111111111111001;
    rom[15354] = 25'b1111111111111111111111001;
    rom[15355] = 25'b1111111111111111111111001;
    rom[15356] = 25'b1111111111111111111111010;
    rom[15357] = 25'b1111111111111111111111010;
    rom[15358] = 25'b1111111111111111111111010;
    rom[15359] = 25'b1111111111111111111111010;
    rom[15360] = 25'b1111111111111111111111010;
    rom[15361] = 25'b1111111111111111111111010;
    rom[15362] = 25'b1111111111111111111111010;
    rom[15363] = 25'b1111111111111111111111010;
    rom[15364] = 25'b1111111111111111111111010;
    rom[15365] = 25'b1111111111111111111111010;
    rom[15366] = 25'b1111111111111111111111010;
    rom[15367] = 25'b1111111111111111111111010;
    rom[15368] = 25'b1111111111111111111111010;
    rom[15369] = 25'b1111111111111111111111010;
    rom[15370] = 25'b1111111111111111111111011;
    rom[15371] = 25'b1111111111111111111111011;
    rom[15372] = 25'b1111111111111111111111011;
    rom[15373] = 25'b1111111111111111111111011;
    rom[15374] = 25'b1111111111111111111111011;
    rom[15375] = 25'b1111111111111111111111011;
    rom[15376] = 25'b1111111111111111111111011;
    rom[15377] = 25'b1111111111111111111111100;
    rom[15378] = 25'b1111111111111111111111100;
    rom[15379] = 25'b1111111111111111111111100;
    rom[15380] = 25'b1111111111111111111111100;
    rom[15381] = 25'b1111111111111111111111100;
    rom[15382] = 25'b1111111111111111111111100;
    rom[15383] = 25'b1111111111111111111111100;
    rom[15384] = 25'b1111111111111111111111101;
    rom[15385] = 25'b1111111111111111111111101;
    rom[15386] = 25'b1111111111111111111111101;
    rom[15387] = 25'b1111111111111111111111101;
    rom[15388] = 25'b1111111111111111111111101;
    rom[15389] = 25'b1111111111111111111111101;
    rom[15390] = 25'b1111111111111111111111101;
    rom[15391] = 25'b1111111111111111111111110;
    rom[15392] = 25'b1111111111111111111111110;
    rom[15393] = 25'b1111111111111111111111110;
    rom[15394] = 25'b1111111111111111111111110;
    rom[15395] = 25'b1111111111111111111111110;
    rom[15396] = 25'b1111111111111111111111110;
    rom[15397] = 25'b1111111111111111111111110;
    rom[15398] = 25'b1111111111111111111111110;
    rom[15399] = 25'b1111111111111111111111111;
    rom[15400] = 25'b1111111111111111111111111;
    rom[15401] = 25'b1111111111111111111111111;
    rom[15402] = 25'b1111111111111111111111111;
    rom[15403] = 25'b1111111111111111111111111;
    rom[15404] = 25'b1111111111111111111111111;
    rom[15405] = 25'b1111111111111111111111111;
    rom[15406] = 25'b1111111111111111111111111;
    rom[15407] = 25'b0000000000000000000000000;
    rom[15408] = 25'b0000000000000000000000000;
    rom[15409] = 25'b0000000000000000000000000;
    rom[15410] = 25'b0000000000000000000000000;
    rom[15411] = 25'b0000000000000000000000000;
    rom[15412] = 25'b0000000000000000000000000;
    rom[15413] = 25'b0000000000000000000000000;
    rom[15414] = 25'b0000000000000000000000000;
    rom[15415] = 25'b0000000000000000000000000;
    rom[15416] = 25'b0000000000000000000000000;
    rom[15417] = 25'b0000000000000000000000000;
    rom[15418] = 25'b0000000000000000000000000;
    rom[15419] = 25'b0000000000000000000000000;
    rom[15420] = 25'b0000000000000000000000000;
    rom[15421] = 25'b0000000000000000000000000;
    rom[15422] = 25'b0000000000000000000000000;
    rom[15423] = 25'b0000000000000000000000000;
    rom[15424] = 25'b0000000000000000000000000;
    rom[15425] = 25'b0000000000000000000000000;
    rom[15426] = 25'b0000000000000000000000000;
    rom[15427] = 25'b0000000000000000000000000;
    rom[15428] = 25'b0000000000000000000000000;
    rom[15429] = 25'b0000000000000000000000000;
    rom[15430] = 25'b0000000000000000000000000;
    rom[15431] = 25'b0000000000000000000000000;
    rom[15432] = 25'b0000000000000000000000000;
    rom[15433] = 25'b0000000000000000000000000;
    rom[15434] = 25'b0000000000000000000000001;
    rom[15435] = 25'b0000000000000000000000001;
    rom[15436] = 25'b0000000000000000000000001;
    rom[15437] = 25'b0000000000000000000000001;
    rom[15438] = 25'b0000000000000000000000001;
    rom[15439] = 25'b0000000000000000000000001;
    rom[15440] = 25'b0000000000000000000000001;
    rom[15441] = 25'b0000000000000000000000001;
    rom[15442] = 25'b0000000000000000000000001;
    rom[15443] = 25'b0000000000000000000000001;
    rom[15444] = 25'b0000000000000000000000010;
    rom[15445] = 25'b0000000000000000000000010;
    rom[15446] = 25'b0000000000000000000000010;
    rom[15447] = 25'b0000000000000000000000010;
    rom[15448] = 25'b0000000000000000000000010;
    rom[15449] = 25'b0000000000000000000000010;
    rom[15450] = 25'b0000000000000000000000010;
    rom[15451] = 25'b0000000000000000000000010;
    rom[15452] = 25'b0000000000000000000000010;
    rom[15453] = 25'b0000000000000000000000010;
    rom[15454] = 25'b0000000000000000000000010;
    rom[15455] = 25'b0000000000000000000000011;
    rom[15456] = 25'b0000000000000000000000011;
    rom[15457] = 25'b0000000000000000000000011;
    rom[15458] = 25'b0000000000000000000000011;
    rom[15459] = 25'b0000000000000000000000011;
    rom[15460] = 25'b0000000000000000000000011;
    rom[15461] = 25'b0000000000000000000000011;
    rom[15462] = 25'b0000000000000000000000011;
    rom[15463] = 25'b0000000000000000000000011;
    rom[15464] = 25'b0000000000000000000000011;
    rom[15465] = 25'b0000000000000000000000011;
    rom[15466] = 25'b0000000000000000000000100;
    rom[15467] = 25'b0000000000000000000000100;
    rom[15468] = 25'b0000000000000000000000100;
    rom[15469] = 25'b0000000000000000000000100;
    rom[15470] = 25'b0000000000000000000000100;
    rom[15471] = 25'b0000000000000000000000100;
    rom[15472] = 25'b0000000000000000000000100;
    rom[15473] = 25'b0000000000000000000000100;
    rom[15474] = 25'b0000000000000000000000100;
    rom[15475] = 25'b0000000000000000000000100;
    rom[15476] = 25'b0000000000000000000000100;
    rom[15477] = 25'b0000000000000000000000100;
    rom[15478] = 25'b0000000000000000000000100;
    rom[15479] = 25'b0000000000000000000000101;
    rom[15480] = 25'b0000000000000000000000101;
    rom[15481] = 25'b0000000000000000000000101;
    rom[15482] = 25'b0000000000000000000000101;
    rom[15483] = 25'b0000000000000000000000101;
    rom[15484] = 25'b0000000000000000000000101;
    rom[15485] = 25'b0000000000000000000000101;
    rom[15486] = 25'b0000000000000000000000101;
    rom[15487] = 25'b0000000000000000000000101;
    rom[15488] = 25'b0000000000000000000000101;
    rom[15489] = 25'b0000000000000000000000101;
    rom[15490] = 25'b0000000000000000000000101;
    rom[15491] = 25'b0000000000000000000000101;
    rom[15492] = 25'b0000000000000000000000101;
    rom[15493] = 25'b0000000000000000000000101;
    rom[15494] = 25'b0000000000000000000000101;
    rom[15495] = 25'b0000000000000000000000101;
    rom[15496] = 25'b0000000000000000000000101;
    rom[15497] = 25'b0000000000000000000000101;
    rom[15498] = 25'b0000000000000000000000101;
    rom[15499] = 25'b0000000000000000000000101;
    rom[15500] = 25'b0000000000000000000000101;
    rom[15501] = 25'b0000000000000000000000101;
    rom[15502] = 25'b0000000000000000000000101;
    rom[15503] = 25'b0000000000000000000000101;
    rom[15504] = 25'b0000000000000000000000101;
    rom[15505] = 25'b0000000000000000000000101;
    rom[15506] = 25'b0000000000000000000000101;
    rom[15507] = 25'b0000000000000000000000101;
    rom[15508] = 25'b0000000000000000000000101;
    rom[15509] = 25'b0000000000000000000000101;
    rom[15510] = 25'b0000000000000000000000101;
    rom[15511] = 25'b0000000000000000000000110;
    rom[15512] = 25'b0000000000000000000000110;
    rom[15513] = 25'b0000000000000000000000110;
    rom[15514] = 25'b0000000000000000000000110;
    rom[15515] = 25'b0000000000000000000000110;
    rom[15516] = 25'b0000000000000000000000110;
    rom[15517] = 25'b0000000000000000000000110;
    rom[15518] = 25'b0000000000000000000000110;
    rom[15519] = 25'b0000000000000000000000110;
    rom[15520] = 25'b0000000000000000000000110;
    rom[15521] = 25'b0000000000000000000000110;
    rom[15522] = 25'b0000000000000000000000110;
    rom[15523] = 25'b0000000000000000000000110;
    rom[15524] = 25'b0000000000000000000000110;
    rom[15525] = 25'b0000000000000000000000110;
    rom[15526] = 25'b0000000000000000000000110;
    rom[15527] = 25'b0000000000000000000000110;
    rom[15528] = 25'b0000000000000000000000110;
    rom[15529] = 25'b0000000000000000000000110;
    rom[15530] = 25'b0000000000000000000000110;
    rom[15531] = 25'b0000000000000000000000110;
    rom[15532] = 25'b0000000000000000000000111;
    rom[15533] = 25'b0000000000000000000000111;
    rom[15534] = 25'b0000000000000000000000111;
    rom[15535] = 25'b0000000000000000000000111;
    rom[15536] = 25'b0000000000000000000000111;
    rom[15537] = 25'b0000000000000000000000111;
    rom[15538] = 25'b0000000000000000000000111;
    rom[15539] = 25'b0000000000000000000000111;
    rom[15540] = 25'b0000000000000000000000111;
    rom[15541] = 25'b0000000000000000000000111;
    rom[15542] = 25'b0000000000000000000000111;
    rom[15543] = 25'b0000000000000000000000111;
    rom[15544] = 25'b0000000000000000000000111;
    rom[15545] = 25'b0000000000000000000000111;
    rom[15546] = 25'b0000000000000000000000111;
    rom[15547] = 25'b0000000000000000000000111;
    rom[15548] = 25'b0000000000000000000000111;
    rom[15549] = 25'b0000000000000000000000111;
    rom[15550] = 25'b0000000000000000000000111;
    rom[15551] = 25'b0000000000000000000000111;
    rom[15552] = 25'b0000000000000000000000111;
    rom[15553] = 25'b0000000000000000000000111;
    rom[15554] = 25'b0000000000000000000000111;
    rom[15555] = 25'b0000000000000000000000111;
    rom[15556] = 25'b0000000000000000000000111;
    rom[15557] = 25'b0000000000000000000000111;
    rom[15558] = 25'b0000000000000000000000111;
    rom[15559] = 25'b0000000000000000000000111;
    rom[15560] = 25'b0000000000000000000000111;
    rom[15561] = 25'b0000000000000000000000111;
    rom[15562] = 25'b0000000000000000000000111;
    rom[15563] = 25'b0000000000000000000000111;
    rom[15564] = 25'b0000000000000000000001000;
    rom[15565] = 25'b0000000000000000000001000;
    rom[15566] = 25'b0000000000000000000001000;
    rom[15567] = 25'b0000000000000000000001000;
    rom[15568] = 25'b0000000000000000000001000;
    rom[15569] = 25'b0000000000000000000001000;
    rom[15570] = 25'b0000000000000000000001000;
    rom[15571] = 25'b0000000000000000000001000;
    rom[15572] = 25'b0000000000000000000001000;
    rom[15573] = 25'b0000000000000000000001000;
    rom[15574] = 25'b0000000000000000000001000;
    rom[15575] = 25'b0000000000000000000001000;
    rom[15576] = 25'b0000000000000000000001000;
    rom[15577] = 25'b0000000000000000000001000;
    rom[15578] = 25'b0000000000000000000001000;
    rom[15579] = 25'b0000000000000000000001000;
    rom[15580] = 25'b0000000000000000000001000;
    rom[15581] = 25'b0000000000000000000001000;
    rom[15582] = 25'b0000000000000000000001000;
    rom[15583] = 25'b0000000000000000000001000;
    rom[15584] = 25'b0000000000000000000001000;
    rom[15585] = 25'b0000000000000000000001000;
    rom[15586] = 25'b0000000000000000000001000;
    rom[15587] = 25'b0000000000000000000001000;
    rom[15588] = 25'b0000000000000000000001000;
    rom[15589] = 25'b0000000000000000000001000;
    rom[15590] = 25'b0000000000000000000001000;
    rom[15591] = 25'b0000000000000000000001000;
    rom[15592] = 25'b0000000000000000000001000;
    rom[15593] = 25'b0000000000000000000001000;
    rom[15594] = 25'b0000000000000000000001000;
    rom[15595] = 25'b0000000000000000000001000;
    rom[15596] = 25'b0000000000000000000001000;
    rom[15597] = 25'b0000000000000000000001000;
    rom[15598] = 25'b0000000000000000000001000;
    rom[15599] = 25'b0000000000000000000001000;
    rom[15600] = 25'b0000000000000000000001000;
    rom[15601] = 25'b0000000000000000000001000;
    rom[15602] = 25'b0000000000000000000001000;
    rom[15603] = 25'b0000000000000000000001000;
    rom[15604] = 25'b0000000000000000000001000;
    rom[15605] = 25'b0000000000000000000001000;
    rom[15606] = 25'b0000000000000000000001000;
    rom[15607] = 25'b0000000000000000000001000;
    rom[15608] = 25'b0000000000000000000001000;
    rom[15609] = 25'b0000000000000000000001000;
    rom[15610] = 25'b0000000000000000000001000;
    rom[15611] = 25'b0000000000000000000001000;
    rom[15612] = 25'b0000000000000000000001000;
    rom[15613] = 25'b0000000000000000000001000;
    rom[15614] = 25'b0000000000000000000001000;
    rom[15615] = 25'b0000000000000000000001000;
    rom[15616] = 25'b0000000000000000000001000;
    rom[15617] = 25'b0000000000000000000001000;
    rom[15618] = 25'b0000000000000000000001000;
    rom[15619] = 25'b0000000000000000000001000;
    rom[15620] = 25'b0000000000000000000001000;
    rom[15621] = 25'b0000000000000000000001000;
    rom[15622] = 25'b0000000000000000000001000;
    rom[15623] = 25'b0000000000000000000001000;
    rom[15624] = 25'b0000000000000000000001000;
    rom[15625] = 25'b0000000000000000000001000;
    rom[15626] = 25'b0000000000000000000001000;
    rom[15627] = 25'b0000000000000000000001000;
    rom[15628] = 25'b0000000000000000000001000;
    rom[15629] = 25'b0000000000000000000001000;
    rom[15630] = 25'b0000000000000000000001000;
    rom[15631] = 25'b0000000000000000000001000;
    rom[15632] = 25'b0000000000000000000001000;
    rom[15633] = 25'b0000000000000000000001000;
    rom[15634] = 25'b0000000000000000000001000;
    rom[15635] = 25'b0000000000000000000001000;
    rom[15636] = 25'b0000000000000000000001000;
    rom[15637] = 25'b0000000000000000000001000;
    rom[15638] = 25'b0000000000000000000001000;
    rom[15639] = 25'b0000000000000000000001000;
    rom[15640] = 25'b0000000000000000000001000;
    rom[15641] = 25'b0000000000000000000001000;
    rom[15642] = 25'b0000000000000000000001000;
    rom[15643] = 25'b0000000000000000000001000;
    rom[15644] = 25'b0000000000000000000001000;
    rom[15645] = 25'b0000000000000000000001000;
    rom[15646] = 25'b0000000000000000000001000;
    rom[15647] = 25'b0000000000000000000001000;
    rom[15648] = 25'b0000000000000000000001000;
    rom[15649] = 25'b0000000000000000000001000;
    rom[15650] = 25'b0000000000000000000001000;
    rom[15651] = 25'b0000000000000000000001000;
    rom[15652] = 25'b0000000000000000000001000;
    rom[15653] = 25'b0000000000000000000001000;
    rom[15654] = 25'b0000000000000000000001000;
    rom[15655] = 25'b0000000000000000000001000;
    rom[15656] = 25'b0000000000000000000001000;
    rom[15657] = 25'b0000000000000000000001000;
    rom[15658] = 25'b0000000000000000000001000;
    rom[15659] = 25'b0000000000000000000001000;
    rom[15660] = 25'b0000000000000000000001000;
    rom[15661] = 25'b0000000000000000000001000;
    rom[15662] = 25'b0000000000000000000001000;
    rom[15663] = 25'b0000000000000000000001000;
    rom[15664] = 25'b0000000000000000000001000;
    rom[15665] = 25'b0000000000000000000001000;
    rom[15666] = 25'b0000000000000000000001000;
    rom[15667] = 25'b0000000000000000000001000;
    rom[15668] = 25'b0000000000000000000001000;
    rom[15669] = 25'b0000000000000000000001000;
    rom[15670] = 25'b0000000000000000000001000;
    rom[15671] = 25'b0000000000000000000001000;
    rom[15672] = 25'b0000000000000000000001000;
    rom[15673] = 25'b0000000000000000000001000;
    rom[15674] = 25'b0000000000000000000001000;
    rom[15675] = 25'b0000000000000000000000111;
    rom[15676] = 25'b0000000000000000000000111;
    rom[15677] = 25'b0000000000000000000000111;
    rom[15678] = 25'b0000000000000000000000111;
    rom[15679] = 25'b0000000000000000000000111;
    rom[15680] = 25'b0000000000000000000000111;
    rom[15681] = 25'b0000000000000000000000111;
    rom[15682] = 25'b0000000000000000000000111;
    rom[15683] = 25'b0000000000000000000000111;
    rom[15684] = 25'b0000000000000000000000111;
    rom[15685] = 25'b0000000000000000000000111;
    rom[15686] = 25'b0000000000000000000000111;
    rom[15687] = 25'b0000000000000000000000111;
    rom[15688] = 25'b0000000000000000000000111;
    rom[15689] = 25'b0000000000000000000000111;
    rom[15690] = 25'b0000000000000000000000111;
    rom[15691] = 25'b0000000000000000000000111;
    rom[15692] = 25'b0000000000000000000000111;
    rom[15693] = 25'b0000000000000000000000111;
    rom[15694] = 25'b0000000000000000000000111;
    rom[15695] = 25'b0000000000000000000000111;
    rom[15696] = 25'b0000000000000000000000111;
    rom[15697] = 25'b0000000000000000000000111;
    rom[15698] = 25'b0000000000000000000000111;
    rom[15699] = 25'b0000000000000000000000111;
    rom[15700] = 25'b0000000000000000000000111;
    rom[15701] = 25'b0000000000000000000000111;
    rom[15702] = 25'b0000000000000000000000111;
    rom[15703] = 25'b0000000000000000000000111;
    rom[15704] = 25'b0000000000000000000000111;
    rom[15705] = 25'b0000000000000000000000111;
    rom[15706] = 25'b0000000000000000000000111;
    rom[15707] = 25'b0000000000000000000000111;
    rom[15708] = 25'b0000000000000000000000111;
    rom[15709] = 25'b0000000000000000000000111;
    rom[15710] = 25'b0000000000000000000000111;
    rom[15711] = 25'b0000000000000000000000111;
    rom[15712] = 25'b0000000000000000000000111;
    rom[15713] = 25'b0000000000000000000000111;
    rom[15714] = 25'b0000000000000000000000111;
    rom[15715] = 25'b0000000000000000000000111;
    rom[15716] = 25'b0000000000000000000000111;
    rom[15717] = 25'b0000000000000000000000110;
    rom[15718] = 25'b0000000000000000000000110;
    rom[15719] = 25'b0000000000000000000000110;
    rom[15720] = 25'b0000000000000000000000110;
    rom[15721] = 25'b0000000000000000000000110;
    rom[15722] = 25'b0000000000000000000000110;
    rom[15723] = 25'b0000000000000000000000110;
    rom[15724] = 25'b0000000000000000000000110;
    rom[15725] = 25'b0000000000000000000000110;
    rom[15726] = 25'b0000000000000000000000110;
    rom[15727] = 25'b0000000000000000000000110;
    rom[15728] = 25'b0000000000000000000000110;
    rom[15729] = 25'b0000000000000000000000110;
    rom[15730] = 25'b0000000000000000000000110;
    rom[15731] = 25'b0000000000000000000000110;
    rom[15732] = 25'b0000000000000000000000110;
    rom[15733] = 25'b0000000000000000000000110;
    rom[15734] = 25'b0000000000000000000000110;
    rom[15735] = 25'b0000000000000000000000110;
    rom[15736] = 25'b0000000000000000000000110;
    rom[15737] = 25'b0000000000000000000000110;
    rom[15738] = 25'b0000000000000000000000110;
    rom[15739] = 25'b0000000000000000000000110;
    rom[15740] = 25'b0000000000000000000000110;
    rom[15741] = 25'b0000000000000000000000110;
    rom[15742] = 25'b0000000000000000000000110;
    rom[15743] = 25'b0000000000000000000000110;
    rom[15744] = 25'b0000000000000000000000110;
    rom[15745] = 25'b0000000000000000000000110;
    rom[15746] = 25'b0000000000000000000000110;
    rom[15747] = 25'b0000000000000000000000110;
    rom[15748] = 25'b0000000000000000000000110;
    rom[15749] = 25'b0000000000000000000000110;
    rom[15750] = 25'b0000000000000000000000110;
    rom[15751] = 25'b0000000000000000000000101;
    rom[15752] = 25'b0000000000000000000000101;
    rom[15753] = 25'b0000000000000000000000101;
    rom[15754] = 25'b0000000000000000000000101;
    rom[15755] = 25'b0000000000000000000000101;
    rom[15756] = 25'b0000000000000000000000101;
    rom[15757] = 25'b0000000000000000000000101;
    rom[15758] = 25'b0000000000000000000000101;
    rom[15759] = 25'b0000000000000000000000101;
    rom[15760] = 25'b0000000000000000000000101;
    rom[15761] = 25'b0000000000000000000000101;
    rom[15762] = 25'b0000000000000000000000101;
    rom[15763] = 25'b0000000000000000000000101;
    rom[15764] = 25'b0000000000000000000000101;
    rom[15765] = 25'b0000000000000000000000101;
    rom[15766] = 25'b0000000000000000000000101;
    rom[15767] = 25'b0000000000000000000000101;
    rom[15768] = 25'b0000000000000000000000101;
    rom[15769] = 25'b0000000000000000000000101;
    rom[15770] = 25'b0000000000000000000000101;
    rom[15771] = 25'b0000000000000000000000101;
    rom[15772] = 25'b0000000000000000000000101;
    rom[15773] = 25'b0000000000000000000000101;
    rom[15774] = 25'b0000000000000000000000101;
    rom[15775] = 25'b0000000000000000000000101;
    rom[15776] = 25'b0000000000000000000000101;
    rom[15777] = 25'b0000000000000000000000101;
    rom[15778] = 25'b0000000000000000000000101;
    rom[15779] = 25'b0000000000000000000000101;
    rom[15780] = 25'b0000000000000000000000101;
    rom[15781] = 25'b0000000000000000000000101;
    rom[15782] = 25'b0000000000000000000000101;
    rom[15783] = 25'b0000000000000000000000101;
    rom[15784] = 25'b0000000000000000000000101;
    rom[15785] = 25'b0000000000000000000000101;
    rom[15786] = 25'b0000000000000000000000101;
    rom[15787] = 25'b0000000000000000000000101;
    rom[15788] = 25'b0000000000000000000000101;
    rom[15789] = 25'b0000000000000000000000101;
    rom[15790] = 25'b0000000000000000000000101;
    rom[15791] = 25'b0000000000000000000000101;
    rom[15792] = 25'b0000000000000000000000101;
    rom[15793] = 25'b0000000000000000000000101;
    rom[15794] = 25'b0000000000000000000000101;
    rom[15795] = 25'b0000000000000000000000101;
    rom[15796] = 25'b0000000000000000000000101;
    rom[15797] = 25'b0000000000000000000000101;
    rom[15798] = 25'b0000000000000000000000101;
    rom[15799] = 25'b0000000000000000000000101;
    rom[15800] = 25'b0000000000000000000000101;
    rom[15801] = 25'b0000000000000000000000101;
    rom[15802] = 25'b0000000000000000000000101;
    rom[15803] = 25'b0000000000000000000000101;
    rom[15804] = 25'b0000000000000000000000101;
    rom[15805] = 25'b0000000000000000000000101;
    rom[15806] = 25'b0000000000000000000000101;
    rom[15807] = 25'b0000000000000000000000101;
    rom[15808] = 25'b0000000000000000000000101;
    rom[15809] = 25'b0000000000000000000000101;
    rom[15810] = 25'b0000000000000000000000100;
    rom[15811] = 25'b0000000000000000000000100;
    rom[15812] = 25'b0000000000000000000000100;
    rom[15813] = 25'b0000000000000000000000100;
    rom[15814] = 25'b0000000000000000000000100;
    rom[15815] = 25'b0000000000000000000000100;
    rom[15816] = 25'b0000000000000000000000100;
    rom[15817] = 25'b0000000000000000000000100;
    rom[15818] = 25'b0000000000000000000000100;
    rom[15819] = 25'b0000000000000000000000100;
    rom[15820] = 25'b0000000000000000000000100;
    rom[15821] = 25'b0000000000000000000000100;
    rom[15822] = 25'b0000000000000000000000100;
    rom[15823] = 25'b0000000000000000000000100;
    rom[15824] = 25'b0000000000000000000000100;
    rom[15825] = 25'b0000000000000000000000100;
    rom[15826] = 25'b0000000000000000000000100;
    rom[15827] = 25'b0000000000000000000000100;
    rom[15828] = 25'b0000000000000000000000100;
    rom[15829] = 25'b0000000000000000000000100;
    rom[15830] = 25'b0000000000000000000000100;
    rom[15831] = 25'b0000000000000000000000100;
    rom[15832] = 25'b0000000000000000000000100;
    rom[15833] = 25'b0000000000000000000000100;
    rom[15834] = 25'b0000000000000000000000100;
    rom[15835] = 25'b0000000000000000000000100;
    rom[15836] = 25'b0000000000000000000000100;
    rom[15837] = 25'b0000000000000000000000100;
    rom[15838] = 25'b0000000000000000000000100;
    rom[15839] = 25'b0000000000000000000000011;
    rom[15840] = 25'b0000000000000000000000011;
    rom[15841] = 25'b0000000000000000000000011;
    rom[15842] = 25'b0000000000000000000000011;
    rom[15843] = 25'b0000000000000000000000011;
    rom[15844] = 25'b0000000000000000000000011;
    rom[15845] = 25'b0000000000000000000000011;
    rom[15846] = 25'b0000000000000000000000011;
    rom[15847] = 25'b0000000000000000000000011;
    rom[15848] = 25'b0000000000000000000000011;
    rom[15849] = 25'b0000000000000000000000011;
    rom[15850] = 25'b0000000000000000000000011;
    rom[15851] = 25'b0000000000000000000000011;
    rom[15852] = 25'b0000000000000000000000011;
    rom[15853] = 25'b0000000000000000000000011;
    rom[15854] = 25'b0000000000000000000000011;
    rom[15855] = 25'b0000000000000000000000011;
    rom[15856] = 25'b0000000000000000000000011;
    rom[15857] = 25'b0000000000000000000000011;
    rom[15858] = 25'b0000000000000000000000011;
    rom[15859] = 25'b0000000000000000000000011;
    rom[15860] = 25'b0000000000000000000000011;
    rom[15861] = 25'b0000000000000000000000011;
    rom[15862] = 25'b0000000000000000000000011;
    rom[15863] = 25'b0000000000000000000000011;
    rom[15864] = 25'b0000000000000000000000011;
    rom[15865] = 25'b0000000000000000000000011;
    rom[15866] = 25'b0000000000000000000000011;
    rom[15867] = 25'b0000000000000000000000011;
    rom[15868] = 25'b0000000000000000000000010;
    rom[15869] = 25'b0000000000000000000000010;
    rom[15870] = 25'b0000000000000000000000010;
    rom[15871] = 25'b0000000000000000000000010;
    rom[15872] = 25'b0000000000000000000000010;
    rom[15873] = 25'b0000000000000000000000010;
    rom[15874] = 25'b0000000000000000000000010;
    rom[15875] = 25'b0000000000000000000000010;
    rom[15876] = 25'b0000000000000000000000010;
    rom[15877] = 25'b0000000000000000000000010;
    rom[15878] = 25'b0000000000000000000000010;
    rom[15879] = 25'b0000000000000000000000010;
    rom[15880] = 25'b0000000000000000000000010;
    rom[15881] = 25'b0000000000000000000000010;
    rom[15882] = 25'b0000000000000000000000010;
    rom[15883] = 25'b0000000000000000000000010;
    rom[15884] = 25'b0000000000000000000000010;
    rom[15885] = 25'b0000000000000000000000010;
    rom[15886] = 25'b0000000000000000000000010;
    rom[15887] = 25'b0000000000000000000000010;
    rom[15888] = 25'b0000000000000000000000010;
    rom[15889] = 25'b0000000000000000000000010;
    rom[15890] = 25'b0000000000000000000000010;
    rom[15891] = 25'b0000000000000000000000010;
    rom[15892] = 25'b0000000000000000000000010;
    rom[15893] = 25'b0000000000000000000000010;
    rom[15894] = 25'b0000000000000000000000010;
    rom[15895] = 25'b0000000000000000000000010;
    rom[15896] = 25'b0000000000000000000000010;
    rom[15897] = 25'b0000000000000000000000010;
    rom[15898] = 25'b0000000000000000000000010;
    rom[15899] = 25'b0000000000000000000000010;
    rom[15900] = 25'b0000000000000000000000001;
    rom[15901] = 25'b0000000000000000000000001;
    rom[15902] = 25'b0000000000000000000000001;
    rom[15903] = 25'b0000000000000000000000001;
    rom[15904] = 25'b0000000000000000000000001;
    rom[15905] = 25'b0000000000000000000000001;
    rom[15906] = 25'b0000000000000000000000001;
    rom[15907] = 25'b0000000000000000000000001;
    rom[15908] = 25'b0000000000000000000000001;
    rom[15909] = 25'b0000000000000000000000001;
    rom[15910] = 25'b0000000000000000000000001;
    rom[15911] = 25'b0000000000000000000000001;
    rom[15912] = 25'b0000000000000000000000001;
    rom[15913] = 25'b0000000000000000000000001;
    rom[15914] = 25'b0000000000000000000000001;
    rom[15915] = 25'b0000000000000000000000001;
    rom[15916] = 25'b0000000000000000000000001;
    rom[15917] = 25'b0000000000000000000000001;
    rom[15918] = 25'b0000000000000000000000001;
    rom[15919] = 25'b0000000000000000000000001;
    rom[15920] = 25'b0000000000000000000000001;
    rom[15921] = 25'b0000000000000000000000001;
    rom[15922] = 25'b0000000000000000000000001;
    rom[15923] = 25'b0000000000000000000000001;
    rom[15924] = 25'b0000000000000000000000001;
    rom[15925] = 25'b0000000000000000000000001;
    rom[15926] = 25'b0000000000000000000000001;
    rom[15927] = 25'b0000000000000000000000001;
    rom[15928] = 25'b0000000000000000000000001;
    rom[15929] = 25'b0000000000000000000000001;
    rom[15930] = 25'b0000000000000000000000001;
    rom[15931] = 25'b0000000000000000000000001;
    rom[15932] = 25'b0000000000000000000000001;
    rom[15933] = 25'b0000000000000000000000001;
    rom[15934] = 25'b0000000000000000000000000;
    rom[15935] = 25'b0000000000000000000000000;
    rom[15936] = 25'b0000000000000000000000000;
    rom[15937] = 25'b0000000000000000000000000;
    rom[15938] = 25'b0000000000000000000000000;
    rom[15939] = 25'b0000000000000000000000000;
    rom[15940] = 25'b0000000000000000000000000;
    rom[15941] = 25'b0000000000000000000000000;
    rom[15942] = 25'b0000000000000000000000000;
    rom[15943] = 25'b0000000000000000000000000;
    rom[15944] = 25'b0000000000000000000000000;
    rom[15945] = 25'b0000000000000000000000000;
    rom[15946] = 25'b0000000000000000000000000;
    rom[15947] = 25'b0000000000000000000000000;
    rom[15948] = 25'b0000000000000000000000000;
    rom[15949] = 25'b0000000000000000000000000;
    rom[15950] = 25'b0000000000000000000000000;
    rom[15951] = 25'b0000000000000000000000000;
    rom[15952] = 25'b0000000000000000000000000;
    rom[15953] = 25'b0000000000000000000000000;
    rom[15954] = 25'b0000000000000000000000000;
    rom[15955] = 25'b0000000000000000000000000;
    rom[15956] = 25'b0000000000000000000000000;
    rom[15957] = 25'b0000000000000000000000000;
    rom[15958] = 25'b0000000000000000000000000;
    rom[15959] = 25'b0000000000000000000000000;
    rom[15960] = 25'b0000000000000000000000000;
    rom[15961] = 25'b0000000000000000000000000;
    rom[15962] = 25'b0000000000000000000000000;
    rom[15963] = 25'b0000000000000000000000000;
    rom[15964] = 25'b0000000000000000000000000;
    rom[15965] = 25'b0000000000000000000000000;
    rom[15966] = 25'b0000000000000000000000000;
    rom[15967] = 25'b0000000000000000000000000;
    rom[15968] = 25'b0000000000000000000000000;
    rom[15969] = 25'b0000000000000000000000000;
    rom[15970] = 25'b0000000000000000000000000;
    rom[15971] = 25'b0000000000000000000000000;
    rom[15972] = 25'b0000000000000000000000000;
    rom[15973] = 25'b0000000000000000000000000;
    rom[15974] = 25'b0000000000000000000000000;
    rom[15975] = 25'b0000000000000000000000000;
    rom[15976] = 25'b0000000000000000000000000;
    rom[15977] = 25'b0000000000000000000000000;
    rom[15978] = 25'b0000000000000000000000000;
    rom[15979] = 25'b0000000000000000000000000;
    rom[15980] = 25'b0000000000000000000000000;
    rom[15981] = 25'b0000000000000000000000000;
    rom[15982] = 25'b0000000000000000000000000;
    rom[15983] = 25'b0000000000000000000000000;
    rom[15984] = 25'b0000000000000000000000000;
    rom[15985] = 25'b0000000000000000000000000;
    rom[15986] = 25'b0000000000000000000000000;
    rom[15987] = 25'b0000000000000000000000000;
    rom[15988] = 25'b0000000000000000000000000;
    rom[15989] = 25'b0000000000000000000000000;
    rom[15990] = 25'b0000000000000000000000000;
    rom[15991] = 25'b0000000000000000000000000;
    rom[15992] = 25'b0000000000000000000000000;
    rom[15993] = 25'b0000000000000000000000000;
    rom[15994] = 25'b0000000000000000000000000;
    rom[15995] = 25'b0000000000000000000000000;
    rom[15996] = 25'b0000000000000000000000000;
    rom[15997] = 25'b0000000000000000000000000;
    rom[15998] = 25'b0000000000000000000000000;
    rom[15999] = 25'b0000000000000000000000000;
    rom[16000] = 25'b0000000000000000000000000;
    rom[16001] = 25'b0000000000000000000000000;
    rom[16002] = 25'b0000000000000000000000000;
    rom[16003] = 25'b0000000000000000000000000;
    rom[16004] = 25'b0000000000000000000000000;
    rom[16005] = 25'b0000000000000000000000000;
    rom[16006] = 25'b0000000000000000000000000;
    rom[16007] = 25'b0000000000000000000000000;
    rom[16008] = 25'b0000000000000000000000000;
    rom[16009] = 25'b0000000000000000000000000;
    rom[16010] = 25'b0000000000000000000000000;
    rom[16011] = 25'b0000000000000000000000000;
    rom[16012] = 25'b0000000000000000000000000;
    rom[16013] = 25'b0000000000000000000000000;
    rom[16014] = 25'b0000000000000000000000000;
    rom[16015] = 25'b0000000000000000000000000;
    rom[16016] = 25'b0000000000000000000000000;
    rom[16017] = 25'b0000000000000000000000000;
    rom[16018] = 25'b0000000000000000000000000;
    rom[16019] = 25'b0000000000000000000000000;
    rom[16020] = 25'b0000000000000000000000000;
    rom[16021] = 25'b0000000000000000000000000;
    rom[16022] = 25'b0000000000000000000000000;
    rom[16023] = 25'b0000000000000000000000000;
    rom[16024] = 25'b0000000000000000000000000;
    rom[16025] = 25'b0000000000000000000000000;
    rom[16026] = 25'b0000000000000000000000000;
    rom[16027] = 25'b0000000000000000000000000;
    rom[16028] = 25'b0000000000000000000000000;
    rom[16029] = 25'b0000000000000000000000000;
    rom[16030] = 25'b0000000000000000000000000;
    rom[16031] = 25'b0000000000000000000000000;
    rom[16032] = 25'b0000000000000000000000000;
    rom[16033] = 25'b0000000000000000000000000;
    rom[16034] = 25'b0000000000000000000000000;
    rom[16035] = 25'b0000000000000000000000000;
    rom[16036] = 25'b0000000000000000000000000;
    rom[16037] = 25'b0000000000000000000000000;
    rom[16038] = 25'b0000000000000000000000000;
    rom[16039] = 25'b0000000000000000000000000;
    rom[16040] = 25'b0000000000000000000000000;
    rom[16041] = 25'b0000000000000000000000000;
    rom[16042] = 25'b0000000000000000000000000;
    rom[16043] = 25'b0000000000000000000000000;
    rom[16044] = 25'b0000000000000000000000000;
    rom[16045] = 25'b0000000000000000000000000;
    rom[16046] = 25'b0000000000000000000000000;
    rom[16047] = 25'b0000000000000000000000000;
    rom[16048] = 25'b0000000000000000000000000;
    rom[16049] = 25'b0000000000000000000000000;
    rom[16050] = 25'b0000000000000000000000000;
    rom[16051] = 25'b0000000000000000000000000;
    rom[16052] = 25'b0000000000000000000000000;
    rom[16053] = 25'b0000000000000000000000000;
    rom[16054] = 25'b0000000000000000000000000;
    rom[16055] = 25'b0000000000000000000000000;
    rom[16056] = 25'b0000000000000000000000000;
    rom[16057] = 25'b0000000000000000000000000;
    rom[16058] = 25'b0000000000000000000000000;
    rom[16059] = 25'b0000000000000000000000000;
    rom[16060] = 25'b0000000000000000000000000;
    rom[16061] = 25'b0000000000000000000000000;
    rom[16062] = 25'b0000000000000000000000000;
    rom[16063] = 25'b0000000000000000000000000;
    rom[16064] = 25'b0000000000000000000000000;
    rom[16065] = 25'b0000000000000000000000000;
    rom[16066] = 25'b0000000000000000000000000;
    rom[16067] = 25'b0000000000000000000000000;
    rom[16068] = 25'b0000000000000000000000000;
    rom[16069] = 25'b0000000000000000000000000;
    rom[16070] = 25'b0000000000000000000000000;
    rom[16071] = 25'b0000000000000000000000000;
    rom[16072] = 25'b0000000000000000000000000;
    rom[16073] = 25'b0000000000000000000000000;
    rom[16074] = 25'b0000000000000000000000000;
    rom[16075] = 25'b0000000000000000000000000;
    rom[16076] = 25'b0000000000000000000000000;
    rom[16077] = 25'b0000000000000000000000000;
    rom[16078] = 25'b0000000000000000000000000;
    rom[16079] = 25'b0000000000000000000000000;
    rom[16080] = 25'b0000000000000000000000000;
    rom[16081] = 25'b0000000000000000000000000;
    rom[16082] = 25'b0000000000000000000000000;
    rom[16083] = 25'b0000000000000000000000000;
    rom[16084] = 25'b0000000000000000000000000;
    rom[16085] = 25'b0000000000000000000000000;
    rom[16086] = 25'b0000000000000000000000000;
    rom[16087] = 25'b0000000000000000000000000;
    rom[16088] = 25'b0000000000000000000000000;
    rom[16089] = 25'b0000000000000000000000000;
    rom[16090] = 25'b0000000000000000000000000;
    rom[16091] = 25'b0000000000000000000000000;
    rom[16092] = 25'b0000000000000000000000000;
    rom[16093] = 25'b0000000000000000000000000;
    rom[16094] = 25'b0000000000000000000000000;
    rom[16095] = 25'b1111111111111111111111111;
    rom[16096] = 25'b1111111111111111111111111;
    rom[16097] = 25'b1111111111111111111111111;
    rom[16098] = 25'b1111111111111111111111111;
    rom[16099] = 25'b1111111111111111111111111;
    rom[16100] = 25'b1111111111111111111111111;
    rom[16101] = 25'b1111111111111111111111111;
    rom[16102] = 25'b1111111111111111111111111;
    rom[16103] = 25'b1111111111111111111111111;
    rom[16104] = 25'b1111111111111111111111111;
    rom[16105] = 25'b1111111111111111111111111;
    rom[16106] = 25'b1111111111111111111111111;
    rom[16107] = 25'b1111111111111111111111111;
    rom[16108] = 25'b1111111111111111111111111;
    rom[16109] = 25'b1111111111111111111111111;
    rom[16110] = 25'b1111111111111111111111111;
    rom[16111] = 25'b1111111111111111111111111;
    rom[16112] = 25'b1111111111111111111111111;
    rom[16113] = 25'b1111111111111111111111111;
    rom[16114] = 25'b1111111111111111111111111;
    rom[16115] = 25'b1111111111111111111111111;
    rom[16116] = 25'b1111111111111111111111111;
    rom[16117] = 25'b1111111111111111111111111;
    rom[16118] = 25'b1111111111111111111111111;
    rom[16119] = 25'b1111111111111111111111111;
    rom[16120] = 25'b1111111111111111111111111;
    rom[16121] = 25'b1111111111111111111111111;
    rom[16122] = 25'b1111111111111111111111111;
    rom[16123] = 25'b1111111111111111111111111;
    rom[16124] = 25'b1111111111111111111111111;
    rom[16125] = 25'b1111111111111111111111111;
    rom[16126] = 25'b1111111111111111111111111;
    rom[16127] = 25'b1111111111111111111111111;
    rom[16128] = 25'b1111111111111111111111111;
    rom[16129] = 25'b1111111111111111111111111;
    rom[16130] = 25'b1111111111111111111111111;
    rom[16131] = 25'b1111111111111111111111111;
    rom[16132] = 25'b1111111111111111111111111;
    rom[16133] = 25'b1111111111111111111111111;
    rom[16134] = 25'b1111111111111111111111111;
    rom[16135] = 25'b1111111111111111111111111;
    rom[16136] = 25'b1111111111111111111111111;
    rom[16137] = 25'b1111111111111111111111111;
    rom[16138] = 25'b1111111111111111111111111;
    rom[16139] = 25'b1111111111111111111111111;
    rom[16140] = 25'b1111111111111111111111111;
    rom[16141] = 25'b1111111111111111111111111;
    rom[16142] = 25'b1111111111111111111111111;
    rom[16143] = 25'b1111111111111111111111111;
    rom[16144] = 25'b1111111111111111111111111;
    rom[16145] = 25'b1111111111111111111111111;
    rom[16146] = 25'b1111111111111111111111111;
    rom[16147] = 25'b1111111111111111111111111;
    rom[16148] = 25'b1111111111111111111111111;
    rom[16149] = 25'b1111111111111111111111111;
    rom[16150] = 25'b1111111111111111111111111;
    rom[16151] = 25'b1111111111111111111111111;
    rom[16152] = 25'b1111111111111111111111111;
    rom[16153] = 25'b1111111111111111111111111;
    rom[16154] = 25'b1111111111111111111111111;
    rom[16155] = 25'b1111111111111111111111111;
    rom[16156] = 25'b1111111111111111111111111;
    rom[16157] = 25'b1111111111111111111111111;
    rom[16158] = 25'b1111111111111111111111111;
    rom[16159] = 25'b1111111111111111111111111;
    rom[16160] = 25'b1111111111111111111111111;
    rom[16161] = 25'b1111111111111111111111111;
    rom[16162] = 25'b1111111111111111111111111;
    rom[16163] = 25'b1111111111111111111111111;
    rom[16164] = 25'b1111111111111111111111111;
    rom[16165] = 25'b1111111111111111111111111;
    rom[16166] = 25'b1111111111111111111111111;
    rom[16167] = 25'b1111111111111111111111111;
    rom[16168] = 25'b1111111111111111111111111;
    rom[16169] = 25'b1111111111111111111111111;
    rom[16170] = 25'b1111111111111111111111111;
    rom[16171] = 25'b1111111111111111111111111;
    rom[16172] = 25'b1111111111111111111111111;
    rom[16173] = 25'b1111111111111111111111111;
    rom[16174] = 25'b1111111111111111111111111;
    rom[16175] = 25'b1111111111111111111111111;
    rom[16176] = 25'b1111111111111111111111111;
    rom[16177] = 25'b1111111111111111111111111;
    rom[16178] = 25'b1111111111111111111111111;
    rom[16179] = 25'b1111111111111111111111111;
    rom[16180] = 25'b1111111111111111111111111;
    rom[16181] = 25'b1111111111111111111111111;
    rom[16182] = 25'b1111111111111111111111111;
    rom[16183] = 25'b1111111111111111111111111;
    rom[16184] = 25'b1111111111111111111111111;
    rom[16185] = 25'b1111111111111111111111111;
    rom[16186] = 25'b1111111111111111111111111;
    rom[16187] = 25'b1111111111111111111111111;
    rom[16188] = 25'b1111111111111111111111111;
    rom[16189] = 25'b1111111111111111111111111;
    rom[16190] = 25'b1111111111111111111111111;
    rom[16191] = 25'b1111111111111111111111111;
    rom[16192] = 25'b1111111111111111111111111;
    rom[16193] = 25'b1111111111111111111111111;
    rom[16194] = 25'b1111111111111111111111111;
    rom[16195] = 25'b1111111111111111111111111;
    rom[16196] = 25'b1111111111111111111111111;
    rom[16197] = 25'b1111111111111111111111111;
    rom[16198] = 25'b1111111111111111111111111;
    rom[16199] = 25'b1111111111111111111111111;
    rom[16200] = 25'b1111111111111111111111111;
    rom[16201] = 25'b1111111111111111111111111;
    rom[16202] = 25'b1111111111111111111111111;
    rom[16203] = 25'b1111111111111111111111111;
    rom[16204] = 25'b1111111111111111111111111;
    rom[16205] = 25'b1111111111111111111111111;
    rom[16206] = 25'b1111111111111111111111111;
    rom[16207] = 25'b1111111111111111111111111;
    rom[16208] = 25'b1111111111111111111111111;
    rom[16209] = 25'b1111111111111111111111111;
    rom[16210] = 25'b1111111111111111111111111;
    rom[16211] = 25'b1111111111111111111111111;
    rom[16212] = 25'b1111111111111111111111111;
    rom[16213] = 25'b1111111111111111111111111;
    rom[16214] = 25'b1111111111111111111111111;
    rom[16215] = 25'b1111111111111111111111111;
    rom[16216] = 25'b1111111111111111111111111;
    rom[16217] = 25'b1111111111111111111111111;
    rom[16218] = 25'b1111111111111111111111111;
    rom[16219] = 25'b1111111111111111111111111;
    rom[16220] = 25'b1111111111111111111111111;
    rom[16221] = 25'b1111111111111111111111111;
    rom[16222] = 25'b1111111111111111111111111;
    rom[16223] = 25'b1111111111111111111111111;
    rom[16224] = 25'b1111111111111111111111111;
    rom[16225] = 25'b1111111111111111111111111;
    rom[16226] = 25'b1111111111111111111111111;
    rom[16227] = 25'b1111111111111111111111111;
    rom[16228] = 25'b1111111111111111111111111;
    rom[16229] = 25'b1111111111111111111111111;
    rom[16230] = 25'b1111111111111111111111111;
    rom[16231] = 25'b1111111111111111111111111;
    rom[16232] = 25'b1111111111111111111111111;
    rom[16233] = 25'b1111111111111111111111111;
    rom[16234] = 25'b1111111111111111111111111;
    rom[16235] = 25'b1111111111111111111111111;
    rom[16236] = 25'b1111111111111111111111111;
    rom[16237] = 25'b1111111111111111111111111;
    rom[16238] = 25'b1111111111111111111111111;
    rom[16239] = 25'b1111111111111111111111111;
    rom[16240] = 25'b1111111111111111111111111;
    rom[16241] = 25'b1111111111111111111111111;
    rom[16242] = 25'b1111111111111111111111111;
    rom[16243] = 25'b1111111111111111111111111;
    rom[16244] = 25'b1111111111111111111111111;
    rom[16245] = 25'b1111111111111111111111111;
    rom[16246] = 25'b1111111111111111111111111;
    rom[16247] = 25'b1111111111111111111111111;
    rom[16248] = 25'b1111111111111111111111111;
    rom[16249] = 25'b1111111111111111111111111;
    rom[16250] = 25'b1111111111111111111111111;
    rom[16251] = 25'b1111111111111111111111111;
    rom[16252] = 25'b1111111111111111111111111;
    rom[16253] = 25'b1111111111111111111111111;
    rom[16254] = 25'b1111111111111111111111111;
    rom[16255] = 25'b1111111111111111111111111;
    rom[16256] = 25'b1111111111111111111111111;
    rom[16257] = 25'b1111111111111111111111111;
    rom[16258] = 25'b1111111111111111111111111;
    rom[16259] = 25'b1111111111111111111111111;
    rom[16260] = 25'b1111111111111111111111111;
    rom[16261] = 25'b1111111111111111111111111;
    rom[16262] = 25'b1111111111111111111111111;
    rom[16263] = 25'b1111111111111111111111111;
    rom[16264] = 25'b1111111111111111111111111;
    rom[16265] = 25'b1111111111111111111111111;
    rom[16266] = 25'b1111111111111111111111111;
    rom[16267] = 25'b1111111111111111111111111;
    rom[16268] = 25'b1111111111111111111111111;
    rom[16269] = 25'b1111111111111111111111111;
    rom[16270] = 25'b1111111111111111111111111;
    rom[16271] = 25'b1111111111111111111111111;
    rom[16272] = 25'b1111111111111111111111111;
    rom[16273] = 25'b1111111111111111111111111;
    rom[16274] = 25'b1111111111111111111111111;
    rom[16275] = 25'b1111111111111111111111111;
    rom[16276] = 25'b1111111111111111111111111;
    rom[16277] = 25'b1111111111111111111111111;
    rom[16278] = 25'b1111111111111111111111111;
    rom[16279] = 25'b1111111111111111111111111;
    rom[16280] = 25'b1111111111111111111111111;
    rom[16281] = 25'b1111111111111111111111111;
    rom[16282] = 25'b1111111111111111111111111;
    rom[16283] = 25'b1111111111111111111111111;
    rom[16284] = 25'b1111111111111111111111111;
    rom[16285] = 25'b1111111111111111111111111;
    rom[16286] = 25'b1111111111111111111111111;
    rom[16287] = 25'b1111111111111111111111111;
    rom[16288] = 25'b1111111111111111111111111;
    rom[16289] = 25'b1111111111111111111111111;
    rom[16290] = 25'b1111111111111111111111111;
    rom[16291] = 25'b1111111111111111111111111;
    rom[16292] = 25'b1111111111111111111111111;
    rom[16293] = 25'b1111111111111111111111111;
    rom[16294] = 25'b1111111111111111111111111;
    rom[16295] = 25'b1111111111111111111111111;
    rom[16296] = 25'b1111111111111111111111111;
    rom[16297] = 25'b1111111111111111111111111;
    rom[16298] = 25'b1111111111111111111111111;
    rom[16299] = 25'b1111111111111111111111111;
    rom[16300] = 25'b1111111111111111111111111;
    rom[16301] = 25'b1111111111111111111111111;
    rom[16302] = 25'b1111111111111111111111111;
    rom[16303] = 25'b1111111111111111111111111;
    rom[16304] = 25'b1111111111111111111111111;
    rom[16305] = 25'b1111111111111111111111111;
    rom[16306] = 25'b1111111111111111111111111;
    rom[16307] = 25'b1111111111111111111111111;
    rom[16308] = 25'b1111111111111111111111111;
    rom[16309] = 25'b1111111111111111111111111;
    rom[16310] = 25'b1111111111111111111111111;
    rom[16311] = 25'b1111111111111111111111111;
    rom[16312] = 25'b1111111111111111111111111;
    rom[16313] = 25'b1111111111111111111111111;
    rom[16314] = 25'b1111111111111111111111111;
    rom[16315] = 25'b1111111111111111111111111;
    rom[16316] = 25'b1111111111111111111111111;
    rom[16317] = 25'b1111111111111111111111111;
    rom[16318] = 25'b1111111111111111111111111;
    rom[16319] = 25'b1111111111111111111111111;
    rom[16320] = 25'b1111111111111111111111111;
    rom[16321] = 25'b1111111111111111111111111;
    rom[16322] = 25'b1111111111111111111111111;
    rom[16323] = 25'b1111111111111111111111111;
    rom[16324] = 25'b1111111111111111111111111;
    rom[16325] = 25'b1111111111111111111111111;
    rom[16326] = 25'b1111111111111111111111111;
    rom[16327] = 25'b1111111111111111111111111;
    rom[16328] = 25'b1111111111111111111111111;
    rom[16329] = 25'b1111111111111111111111111;
    rom[16330] = 25'b1111111111111111111111111;
    rom[16331] = 25'b1111111111111111111111111;
    rom[16332] = 25'b1111111111111111111111111;
    rom[16333] = 25'b1111111111111111111111111;
    rom[16334] = 25'b1111111111111111111111111;
    rom[16335] = 25'b1111111111111111111111111;
    rom[16336] = 25'b1111111111111111111111111;
    rom[16337] = 25'b1111111111111111111111111;
    rom[16338] = 25'b1111111111111111111111111;
    rom[16339] = 25'b1111111111111111111111111;
    rom[16340] = 25'b1111111111111111111111111;
    rom[16341] = 25'b1111111111111111111111111;
    rom[16342] = 25'b1111111111111111111111111;
    rom[16343] = 25'b1111111111111111111111111;
    rom[16344] = 25'b1111111111111111111111111;
    rom[16345] = 25'b1111111111111111111111111;
    rom[16346] = 25'b1111111111111111111111111;
    rom[16347] = 25'b1111111111111111111111111;
    rom[16348] = 25'b1111111111111111111111111;
    rom[16349] = 25'b1111111111111111111111111;
    rom[16350] = 25'b1111111111111111111111111;
    rom[16351] = 25'b1111111111111111111111111;
    rom[16352] = 25'b1111111111111111111111111;
    rom[16353] = 25'b1111111111111111111111111;
    rom[16354] = 25'b1111111111111111111111111;
    rom[16355] = 25'b1111111111111111111111111;
    rom[16356] = 25'b1111111111111111111111111;
    rom[16357] = 25'b1111111111111111111111111;
    rom[16358] = 25'b1111111111111111111111111;
    rom[16359] = 25'b1111111111111111111111111;
    rom[16360] = 25'b1111111111111111111111111;
    rom[16361] = 25'b1111111111111111111111111;
    rom[16362] = 25'b1111111111111111111111111;
    rom[16363] = 25'b1111111111111111111111111;
    rom[16364] = 25'b1111111111111111111111111;
    rom[16365] = 25'b1111111111111111111111111;
    rom[16366] = 25'b1111111111111111111111111;
    rom[16367] = 25'b1111111111111111111111111;
    rom[16368] = 25'b1111111111111111111111111;
    rom[16369] = 25'b1111111111111111111111111;
    rom[16370] = 25'b1111111111111111111111111;
    rom[16371] = 25'b1111111111111111111111111;
    rom[16372] = 25'b1111111111111111111111111;
    rom[16373] = 25'b1111111111111111111111111;
    rom[16374] = 25'b1111111111111111111111111;
    rom[16375] = 25'b1111111111111111111111111;
    rom[16376] = 25'b1111111111111111111111111;
    rom[16377] = 25'b1111111111111111111111111;
    rom[16378] = 25'b1111111111111111111111111;
    rom[16379] = 25'b1111111111111111111111111;
    rom[16380] = 25'b1111111111111111111111111;
    rom[16381] = 25'b1111111111111111111111111;
    rom[16382] = 25'b1111111111111111111111111;
    rom[16383] = 25'b1111111111111111111111111;
end

// port a
always @(posedge clk)
begin
    if (wea_d == 1'b1) begin
      rom[addra_d] <= dia_d;
    end
    wea_d <= wea;
    dia_d <= dia;
    addra_d <= addra;
end

// port b
always @(posedge clk)
begin
    addrb_d <= addrb;
    rom_pipea <= rom[addrb_d];
    dob_d <= rom_pipea;
end

endmodule
