
/*****************************************************************************/
//
// Author      : Phil Vallance
// File        : exp_shift_sp_rom.v
// Description : Implements a single port RAM with block ram. The ram is a fully
//               pipelined implementation -- 3 clock cycles from new read address
//               to new data                                                     
//
//
/*****************************************************************************/


module exp_shift_sp_rom
(
  input clk, 

  input [7:0] addra,
  output [15:0] doa
);

(* rom_style = "distributed" *) reg [15:0] rom [255:0];
reg [7:0] addra_d;
reg [15:0] doa_d;
reg [15:0] rom_pipea;

assign doa = doa_d;

initial
begin
    rom[0] = 16'b1000000000000000;
    rom[1] = 16'b0111111110100111;
    rom[2] = 16'b0111111101001111;
    rom[3] = 16'b0111111011110111;
    rom[4] = 16'b0111111010011111;
    rom[5] = 16'b0111111001000111;
    rom[6] = 16'b0111110111110000;
    rom[7] = 16'b0111110110011001;
    rom[8] = 16'b0111110101000010;
    rom[9] = 16'b0111110011101011;
    rom[10] = 16'b0111110010010101;
    rom[11] = 16'b0111110000111110;
    rom[12] = 16'b0111101111101000;
    rom[13] = 16'b0111101110010011;
    rom[14] = 16'b0111101100111101;
    rom[15] = 16'b0111101011101000;
    rom[16] = 16'b0111101010010011;
    rom[17] = 16'b0111101000111110;
    rom[18] = 16'b0111100111101001;
    rom[19] = 16'b0111100110010101;
    rom[20] = 16'b0111100101000001;
    rom[21] = 16'b0111100011101101;
    rom[22] = 16'b0111100010011001;
    rom[23] = 16'b0111100001000110;
    rom[24] = 16'b0111011111110010;
    rom[25] = 16'b0111011110011111;
    rom[26] = 16'b0111011101001101;
    rom[27] = 16'b0111011011111010;
    rom[28] = 16'b0111011010101000;
    rom[29] = 16'b0111011001010101;
    rom[30] = 16'b0111011000000100;
    rom[31] = 16'b0111010110110010;
    rom[32] = 16'b0111010101100000;
    rom[33] = 16'b0111010100001111;
    rom[34] = 16'b0111010010111110;
    rom[35] = 16'b0111010001101101;
    rom[36] = 16'b0111010000011101;
    rom[37] = 16'b0111001111001100;
    rom[38] = 16'b0111001101111100;
    rom[39] = 16'b0111001100101100;
    rom[40] = 16'b0111001011011101;
    rom[41] = 16'b0111001010001101;
    rom[42] = 16'b0111001000111110;
    rom[43] = 16'b0111000111101111;
    rom[44] = 16'b0111000110100000;
    rom[45] = 16'b0111000101010001;
    rom[46] = 16'b0111000100000011;
    rom[47] = 16'b0111000010110100;
    rom[48] = 16'b0111000001100110;
    rom[49] = 16'b0111000000011001;
    rom[50] = 16'b0110111111001011;
    rom[51] = 16'b0110111101111110;
    rom[52] = 16'b0110111100110000;
    rom[53] = 16'b0110111011100100;
    rom[54] = 16'b0110111010010111;
    rom[55] = 16'b0110111001001010;
    rom[56] = 16'b0110110111111110;
    rom[57] = 16'b0110110110110010;
    rom[58] = 16'b0110110101100110;
    rom[59] = 16'b0110110100011010;
    rom[60] = 16'b0110110011001111;
    rom[61] = 16'b0110110010000011;
    rom[62] = 16'b0110110000111000;
    rom[63] = 16'b0110101111101101;
    rom[64] = 16'b0110101110100010;
    rom[65] = 16'b0110101101011000;
    rom[66] = 16'b0110101100001110;
    rom[67] = 16'b0110101011000100;
    rom[68] = 16'b0110101001111010;
    rom[69] = 16'b0110101000110000;
    rom[70] = 16'b0110100111100110;
    rom[71] = 16'b0110100110011101;
    rom[72] = 16'b0110100101010100;
    rom[73] = 16'b0110100100001011;
    rom[74] = 16'b0110100011000010;
    rom[75] = 16'b0110100001111010;
    rom[76] = 16'b0110100000110010;
    rom[77] = 16'b0110011111101001;
    rom[78] = 16'b0110011110100010;
    rom[79] = 16'b0110011101011010;
    rom[80] = 16'b0110011100010010;
    rom[81] = 16'b0110011011001011;
    rom[82] = 16'b0110011010000100;
    rom[83] = 16'b0110011000111101;
    rom[84] = 16'b0110010111110110;
    rom[85] = 16'b0110010110101111;
    rom[86] = 16'b0110010101101001;
    rom[87] = 16'b0110010100100011;
    rom[88] = 16'b0110010011011101;
    rom[89] = 16'b0110010010010111;
    rom[90] = 16'b0110010001010001;
    rom[91] = 16'b0110010000001100;
    rom[92] = 16'b0110001111000111;
    rom[93] = 16'b0110001110000010;
    rom[94] = 16'b0110001100111101;
    rom[95] = 16'b0110001011111000;
    rom[96] = 16'b0110001010110100;
    rom[97] = 16'b0110001001101111;
    rom[98] = 16'b0110001000101011;
    rom[99] = 16'b0110000111100111;
    rom[100] = 16'b0110000110100011;
    rom[101] = 16'b0110000101100000;
    rom[102] = 16'b0110000100011100;
    rom[103] = 16'b0110000011011001;
    rom[104] = 16'b0110000010010110;
    rom[105] = 16'b0110000001010011;
    rom[106] = 16'b0110000000010001;
    rom[107] = 16'b0101111111001110;
    rom[108] = 16'b0101111110001100;
    rom[109] = 16'b0101111101001010;
    rom[110] = 16'b0101111100001000;
    rom[111] = 16'b0101111011000110;
    rom[112] = 16'b0101111010000100;
    rom[113] = 16'b0101111001000011;
    rom[114] = 16'b0101111000000010;
    rom[115] = 16'b0101110111000001;
    rom[116] = 16'b0101110110000000;
    rom[117] = 16'b0101110100111111;
    rom[118] = 16'b0101110011111110;
    rom[119] = 16'b0101110010111110;
    rom[120] = 16'b0101110001111110;
    rom[121] = 16'b0101110000111110;
    rom[122] = 16'b0101101111111110;
    rom[123] = 16'b0101101110111110;
    rom[124] = 16'b0101101101111111;
    rom[125] = 16'b0101101100111111;
    rom[126] = 16'b0101101100000000;
    rom[127] = 16'b0101101011000001;
    rom[128] = 16'b0101101010000010;
    rom[129] = 16'b0101101001000100;
    rom[130] = 16'b0101101000000101;
    rom[131] = 16'b0101100111000111;
    rom[132] = 16'b0101100110001001;
    rom[133] = 16'b0101100101001011;
    rom[134] = 16'b0101100100001101;
    rom[135] = 16'b0101100011001111;
    rom[136] = 16'b0101100010010010;
    rom[137] = 16'b0101100001010101;
    rom[138] = 16'b0101100000011000;
    rom[139] = 16'b0101011111011011;
    rom[140] = 16'b0101011110011110;
    rom[141] = 16'b0101011101100001;
    rom[142] = 16'b0101011100100101;
    rom[143] = 16'b0101011011101000;
    rom[144] = 16'b0101011010101100;
    rom[145] = 16'b0101011001110000;
    rom[146] = 16'b0101011000110100;
    rom[147] = 16'b0101010111111001;
    rom[148] = 16'b0101010110111101;
    rom[149] = 16'b0101010110000010;
    rom[150] = 16'b0101010101000111;
    rom[151] = 16'b0101010100001100;
    rom[152] = 16'b0101010011010001;
    rom[153] = 16'b0101010010010110;
    rom[154] = 16'b0101010001011011;
    rom[155] = 16'b0101010000100001;
    rom[156] = 16'b0101001111100111;
    rom[157] = 16'b0101001110101101;
    rom[158] = 16'b0101001101110011;
    rom[159] = 16'b0101001100111001;
    rom[160] = 16'b0101001011111111;
    rom[161] = 16'b0101001011000110;
    rom[162] = 16'b0101001010001101;
    rom[163] = 16'b0101001001010100;
    rom[164] = 16'b0101001000011011;
    rom[165] = 16'b0101000111100010;
    rom[166] = 16'b0101000110101001;
    rom[167] = 16'b0101000101110001;
    rom[168] = 16'b0101000100111000;
    rom[169] = 16'b0101000100000000;
    rom[170] = 16'b0101000011001000;
    rom[171] = 16'b0101000010010000;
    rom[172] = 16'b0101000001011000;
    rom[173] = 16'b0101000000100001;
    rom[174] = 16'b0100111111101001;
    rom[175] = 16'b0100111110110010;
    rom[176] = 16'b0100111101111011;
    rom[177] = 16'b0100111101000100;
    rom[178] = 16'b0100111100001101;
    rom[179] = 16'b0100111011010110;
    rom[180] = 16'b0100111010011111;
    rom[181] = 16'b0100111001101001;
    rom[182] = 16'b0100111000110011;
    rom[183] = 16'b0100110111111101;
    rom[184] = 16'b0100110111000111;
    rom[185] = 16'b0100110110010001;
    rom[186] = 16'b0100110101011011;
    rom[187] = 16'b0100110100100110;
    rom[188] = 16'b0100110011110000;
    rom[189] = 16'b0100110010111011;
    rom[190] = 16'b0100110010000110;
    rom[191] = 16'b0100110001010001;
    rom[192] = 16'b0100110000011100;
    rom[193] = 16'b0100101111100111;
    rom[194] = 16'b0100101110110011;
    rom[195] = 16'b0100101101111110;
    rom[196] = 16'b0100101101001010;
    rom[197] = 16'b0100101100010110;
    rom[198] = 16'b0100101011100010;
    rom[199] = 16'b0100101010101110;
    rom[200] = 16'b0100101001111010;
    rom[201] = 16'b0100101001000111;
    rom[202] = 16'b0100101000010011;
    rom[203] = 16'b0100100111100000;
    rom[204] = 16'b0100100110101101;
    rom[205] = 16'b0100100101111010;
    rom[206] = 16'b0100100101000111;
    rom[207] = 16'b0100100100010100;
    rom[208] = 16'b0100100011100010;
    rom[209] = 16'b0100100010101111;
    rom[210] = 16'b0100100001111101;
    rom[211] = 16'b0100100001001011;
    rom[212] = 16'b0100100000011001;
    rom[213] = 16'b0100011111100111;
    rom[214] = 16'b0100011110110101;
    rom[215] = 16'b0100011110000100;
    rom[216] = 16'b0100011101010010;
    rom[217] = 16'b0100011100100001;
    rom[218] = 16'b0100011011110000;
    rom[219] = 16'b0100011010111110;
    rom[220] = 16'b0100011010001101;
    rom[221] = 16'b0100011001011101;
    rom[222] = 16'b0100011000101100;
    rom[223] = 16'b0100010111111011;
    rom[224] = 16'b0100010111001011;
    rom[225] = 16'b0100010110011011;
    rom[226] = 16'b0100010101101010;
    rom[227] = 16'b0100010100111010;
    rom[228] = 16'b0100010100001010;
    rom[229] = 16'b0100010011011011;
    rom[230] = 16'b0100010010101011;
    rom[231] = 16'b0100010001111011;
    rom[232] = 16'b0100010001001100;
    rom[233] = 16'b0100010000011101;
    rom[234] = 16'b0100001111101110;
    rom[235] = 16'b0100001110111111;
    rom[236] = 16'b0100001110010000;
    rom[237] = 16'b0100001101100001;
    rom[238] = 16'b0100001100110010;
    rom[239] = 16'b0100001100000100;
    rom[240] = 16'b0100001011010101;
    rom[241] = 16'b0100001010100111;
    rom[242] = 16'b0100001001111001;
    rom[243] = 16'b0100001001001011;
    rom[244] = 16'b0100001000011101;
    rom[245] = 16'b0100000111101111;
    rom[246] = 16'b0100000111000010;
    rom[247] = 16'b0100000110010100;
    rom[248] = 16'b0100000101100111;
    rom[249] = 16'b0100000100111001;
    rom[250] = 16'b0100000100001100;
    rom[251] = 16'b0100000011011111;
    rom[252] = 16'b0100000010110010;
    rom[253] = 16'b0100000010000110;
    rom[254] = 16'b0100000001011001;
    rom[255] = 16'b0100000000101100;
end


always @(posedge clk)
begin
    addra_d <= addra;
    rom_pipea <= rom[addra_d];
    doa_d <= rom_pipea;
end
endmodule
