//
// Macros used only in simulation.
//
//
`ifndef SIM_BIN_WRITE
`define SIM_BIN_WRITE 1 // Default: 100 ms
`endif
